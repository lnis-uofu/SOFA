VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_1__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 134.32 BY 97.92 ;
  SYMMETRY X Y ;
  PIN pReset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.12 97.435 58.26 97.92 ;
    END
  END pReset[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.75 97.12 99.05 97.92 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.6 97.435 75.74 97.92 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.68 97.435 51.82 97.92 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.35 97.12 80.65 97.92 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.23 97.12 70.53 97.92 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.03 97.12 61.33 97.92 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.03 97.12 84.33 97.92 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.56 97.435 87.7 97.92 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.31 97.12 92.61 97.92 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.8 97.435 84.94 97.92 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.72 97.435 85.86 97.92 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.04 97.435 82.18 97.92 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.55 97.12 66.85 97.92 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 82.19 97.12 82.49 97.92 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.47 97.12 90.77 97.92 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.04 97.435 59.18 97.92 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.52 97.435 99.66 97.92 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.94 97.435 66.08 97.92 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.92 97.435 95.06 97.92 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.51 97.12 78.81 97.92 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.39 97.12 68.69 97.92 ;
    END
  END chany_top_in[20]
  PIN chany_top_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.87 97.12 63.17 97.92 ;
    END
  END chany_top_in[21]
  PIN chany_top_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.44 97.435 100.58 97.92 ;
    END
  END chany_top_in[22]
  PIN chany_top_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.44 97.435 77.58 97.92 ;
    END
  END chany_top_in[23]
  PIN chany_top_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 76.67 97.12 76.97 97.92 ;
    END
  END chany_top_in[24]
  PIN chany_top_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 64.71 97.12 65.01 97.92 ;
    END
  END chany_top_in[25]
  PIN chany_top_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.15 97.12 94.45 97.92 ;
    END
  END chany_top_in[26]
  PIN chany_top_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94 97.435 94.14 97.92 ;
    END
  END chany_top_in[27]
  PIN chany_top_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.87 97.12 86.17 97.92 ;
    END
  END chany_top_in[28]
  PIN chany_top_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.86 97.435 90 97.92 ;
    END
  END chany_top_in[29]
  PIN top_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 30.36 91.56 30.955 91.7 ;
    END
  END top_left_grid_pin_44_[0]
  PIN top_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.96 86.555 14.1 87.04 ;
    END
  END top_left_grid_pin_45_[0]
  PIN top_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 30.36 90.88 30.955 91.02 ;
    END
  END top_left_grid_pin_46_[0]
  PIN top_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.82 86.555 9.96 87.04 ;
    END
  END top_left_grid_pin_47_[0]
  PIN top_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 30.36 91.99 31.16 92.29 ;
    END
  END top_left_grid_pin_48_[0]
  PIN top_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.56 86.555 18.7 87.04 ;
    END
  END top_left_grid_pin_49_[0]
  PIN top_left_grid_pin_50_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 30.36 88.84 30.955 88.98 ;
    END
  END top_left_grid_pin_50_[0]
  PIN top_left_grid_pin_51_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.64 86.555 17.78 87.04 ;
    END
  END top_left_grid_pin_51_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 68.78 134.32 68.92 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 69.46 134.32 69.6 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 43.03 134.32 43.33 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 41.67 134.32 41.97 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 26.71 134.32 27.01 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 52.55 134.32 52.85 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 51.19 134.32 51.49 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 49.74 134.32 49.88 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 45.75 134.32 46.05 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 40.31 134.32 40.61 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 52.46 134.32 52.6 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 44.3 134.32 44.44 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 29.43 134.32 29.73 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 47.11 134.32 47.41 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 53.14 134.32 53.28 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 79.66 134.32 79.8 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 44.39 134.32 44.69 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 41.58 134.32 41.72 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 60.71 134.32 61.01 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 36.14 134.32 36.28 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 47.7 134.32 47.84 ;
    END
  END chanx_right_in[20]
  PIN chanx_right_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 74.9 134.32 75.04 ;
    END
  END chanx_right_in[21]
  PIN chanx_right_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 50.42 134.32 50.56 ;
    END
  END chanx_right_in[22]
  PIN chanx_right_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 34.44 134.32 34.58 ;
    END
  END chanx_right_in[23]
  PIN chanx_right_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 49.83 134.32 50.13 ;
    END
  END chanx_right_in[24]
  PIN chanx_right_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 42.26 134.32 42.4 ;
    END
  END chanx_right_in[25]
  PIN chanx_right_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 62.07 134.32 62.37 ;
    END
  END chanx_right_in[26]
  PIN chanx_right_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 53.91 134.32 54.21 ;
    END
  END chanx_right_in[27]
  PIN chanx_right_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 29 134.32 29.14 ;
    END
  END chanx_right_in[28]
  PIN chanx_right_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 48.47 134.32 48.77 ;
    END
  END chanx_right_in[29]
  PIN right_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 6.22 103.96 6.36 ;
    END
  END right_bottom_grid_pin_36_[0]
  PIN right_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 12.68 134.32 12.82 ;
    END
  END right_bottom_grid_pin_37_[0]
  PIN right_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.14 10.88 121.28 11.365 ;
    END
  END right_bottom_grid_pin_38_[0]
  PIN right_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 14.38 134.32 14.52 ;
    END
  END right_bottom_grid_pin_39_[0]
  PIN right_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.9 10.88 124.04 11.365 ;
    END
  END right_bottom_grid_pin_40_[0]
  PIN right_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 1.8 103.96 1.94 ;
    END
  END right_bottom_grid_pin_41_[0]
  PIN right_bottom_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 6.9 103.96 7.04 ;
    END
  END right_bottom_grid_pin_42_[0]
  PIN right_bottom_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.82 10.88 124.96 11.365 ;
    END
  END right_bottom_grid_pin_43_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.27 0 58.57 0.8 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.36 0 55.5 0.485 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.39 0 68.69 0.8 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94 0 94.14 0.485 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.35 0 80.65 0.8 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.75 0 99.05 0.8 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.82 0 78.96 0.485 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.55 0 66.85 0.8 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 76.67 0 76.97 0.8 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.95 0 85.25 0.8 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.31 0 92.61 0.8 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.12 0 58.26 0.485 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.08 0 93.22 0.485 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 71.15 0 71.45 0.8 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.88 0 84.02 0.485 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.52 0 99.66 0.485 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.44 0 100.58 0.485 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 64.71 0 65.01 0.8 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.24 0 68.38 0.485 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.72 0 85.86 0.485 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.78 0 44.92 0.485 ;
    END
  END chany_bottom_in[20]
  PIN chany_bottom_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.87 0 63.17 0.8 ;
    END
  END chany_bottom_in[21]
  PIN chany_bottom_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.04 0 59.18 0.485 ;
    END
  END chany_bottom_in[22]
  PIN chany_bottom_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.48 0 65.62 0.485 ;
    END
  END chany_bottom_in[23]
  PIN chany_bottom_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.47 0 90.77 0.8 ;
    END
  END chany_bottom_in[24]
  PIN chany_bottom_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.56 0 87.7 0.485 ;
    END
  END chany_bottom_in[25]
  PIN chany_bottom_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.15 0 94.45 0.8 ;
    END
  END chany_bottom_in[26]
  PIN chany_bottom_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.24 0 91.38 0.485 ;
    END
  END chany_bottom_in[27]
  PIN chany_bottom_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.51 0 78.81 0.8 ;
    END
  END chany_bottom_in[28]
  PIN chany_bottom_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.16 0 69.3 0.485 ;
    END
  END chany_bottom_in[29]
  PIN bottom_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.44 10.88 8.58 11.365 ;
    END
  END bottom_left_grid_pin_44_[0]
  PIN bottom_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.2 10.88 11.34 11.365 ;
    END
  END bottom_left_grid_pin_45_[0]
  PIN bottom_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 30.36 5.63 31.16 5.93 ;
    END
  END bottom_left_grid_pin_46_[0]
  PIN bottom_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.94 10.88 20.08 11.365 ;
    END
  END bottom_left_grid_pin_47_[0]
  PIN bottom_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 30.36 6.22 30.955 6.36 ;
    END
  END bottom_left_grid_pin_48_[0]
  PIN bottom_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.1 10.88 18.24 11.365 ;
    END
  END bottom_left_grid_pin_49_[0]
  PIN bottom_left_grid_pin_50_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.72 10.88 16.86 11.365 ;
    END
  END bottom_left_grid_pin_50_[0]
  PIN bottom_left_grid_pin_51_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.8 10.88 15.94 11.365 ;
    END
  END bottom_left_grid_pin_51_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 49.83 0.8 50.13 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 50.42 0.595 50.56 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 69.46 0.595 69.6 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 79.66 0.595 79.8 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 30.79 0.8 31.09 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 47.7 0.595 47.84 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.55 0.8 52.85 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 45.75 0.8 46.05 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 51.19 0.8 51.49 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 53.14 0.595 53.28 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 40.31 0.8 40.61 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.39 0.8 44.69 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.03 0.8 43.33 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 44.98 0.595 45.12 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 74.9 0.595 75.04 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 29 0.595 29.14 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 77.62 0.595 77.76 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 82.38 0.595 82.52 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 52.46 0.595 52.6 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 72.18 0.595 72.32 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 47.11 0.8 47.41 ;
    END
  END chanx_left_in[20]
  PIN chanx_left_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 71.5 0.595 71.64 ;
    END
  END chanx_left_in[21]
  PIN chanx_left_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.47 0.8 48.77 ;
    END
  END chanx_left_in[22]
  PIN chanx_left_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 55.52 0.595 55.66 ;
    END
  END chanx_left_in[23]
  PIN chanx_left_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 53.91 0.8 54.21 ;
    END
  END chanx_left_in[24]
  PIN chanx_left_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 47.02 0.595 47.16 ;
    END
  END chanx_left_in[25]
  PIN chanx_left_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 49.74 0.595 49.88 ;
    END
  END chanx_left_in[26]
  PIN chanx_left_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 41.67 0.8 41.97 ;
    END
  END chanx_left_in[27]
  PIN chanx_left_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 80.34 0.595 80.48 ;
    END
  END chanx_left_in[28]
  PIN chanx_left_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.23 0.8 36.53 ;
    END
  END chanx_left_in[29]
  PIN left_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.12 10.88 12.26 11.365 ;
    END
  END left_bottom_grid_pin_36_[0]
  PIN left_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.6 10.88 6.74 11.365 ;
    END
  END left_bottom_grid_pin_37_[0]
  PIN left_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.28 10.88 10.42 11.365 ;
    END
  END left_bottom_grid_pin_38_[0]
  PIN left_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.36 10.88 9.5 11.365 ;
    END
  END left_bottom_grid_pin_39_[0]
  PIN left_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.04 10.88 13.18 11.365 ;
    END
  END left_bottom_grid_pin_40_[0]
  PIN left_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.96 10.88 14.1 11.365 ;
    END
  END left_bottom_grid_pin_41_[0]
  PIN left_bottom_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.52 10.88 7.66 11.365 ;
    END
  END left_bottom_grid_pin_42_[0]
  PIN left_bottom_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.88 10.88 15.02 11.365 ;
    END
  END left_bottom_grid_pin_43_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 71.5 134.32 71.64 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.12 97.435 81.26 97.92 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.2 97.435 80.34 97.92 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.48 97.435 42.62 97.92 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.64 97.435 86.78 97.92 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.92 97.435 72.06 97.92 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 97.435 41.24 97.92 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.88 97.435 84.02 97.92 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.3 97.435 73.44 97.92 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.7 97.435 68.84 97.92 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.18 97.435 63.32 97.92 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.8 97.435 61.94 97.92 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.92 97.435 49.06 97.92 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.27 97.12 58.57 97.92 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.36 97.435 78.5 97.92 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.32 97.435 44.46 97.92 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.36 97.435 101.5 97.92 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.28 97.435 79.42 97.92 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.62 97.435 46.76 97.92 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.86 97.435 67 97.92 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.07 97.12 72.37 97.92 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48 97.435 48.14 97.92 ;
    END
  END chany_top_out[20]
  PIN chany_top_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.08 97.435 93.22 97.92 ;
    END
  END chany_top_out[21]
  PIN chany_top_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.88 97.435 61.02 97.92 ;
    END
  END chany_top_out[22]
  PIN chany_top_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.88 97.435 38.02 97.92 ;
    END
  END chany_top_out[23]
  PIN chany_top_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.52 97.435 76.66 97.92 ;
    END
  END chany_top_out[24]
  PIN chany_top_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.78 97.435 67.92 97.92 ;
    END
  END chany_top_out[25]
  PIN chany_top_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.96 97.435 37.1 97.92 ;
    END
  END chany_top_out[26]
  PIN chany_top_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 97.435 65.16 97.92 ;
    END
  END chany_top_out[27]
  PIN chany_top_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.62 97.435 69.76 97.92 ;
    END
  END chany_top_out[28]
  PIN chany_top_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 97.435 64.24 97.92 ;
    END
  END chany_top_out[29]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 56.2 134.32 56.34 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 36.82 134.32 36.96 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 27.98 134.32 28.12 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 38.86 134.32 39 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 76.94 134.32 77.08 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 31.04 134.32 31.18 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 55.52 134.32 55.66 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 55.27 134.32 55.57 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 57.99 134.32 58.29 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 56.63 134.32 56.93 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 37.59 134.32 37.89 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 59.35 134.32 59.65 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 31.72 134.32 31.86 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 77.62 134.32 77.76 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 32.15 134.32 32.45 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 33.51 134.32 33.81 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 74.22 134.32 74.36 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 72.18 134.32 72.32 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 39.54 134.32 39.68 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 25.35 134.32 25.65 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 28.07 134.32 28.37 ;
    END
  END chanx_right_out[20]
  PIN chanx_right_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 34.87 134.32 35.17 ;
    END
  END chanx_right_out[21]
  PIN chanx_right_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 25.94 134.32 26.08 ;
    END
  END chanx_right_out[22]
  PIN chanx_right_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 22.54 134.32 22.68 ;
    END
  END chanx_right_out[23]
  PIN chanx_right_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 30.79 134.32 31.09 ;
    END
  END chanx_right_out[24]
  PIN chanx_right_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 23.22 134.32 23.36 ;
    END
  END chanx_right_out[25]
  PIN chanx_right_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 38.95 134.32 39.25 ;
    END
  END chanx_right_out[26]
  PIN chanx_right_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 36.23 134.32 36.53 ;
    END
  END chanx_right_out[27]
  PIN chanx_right_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 25.26 134.32 25.4 ;
    END
  END chanx_right_out[28]
  PIN chanx_right_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 33.76 134.32 33.9 ;
    END
  END chanx_right_out[29]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.14 0 75.28 0.485 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.7 0 45.84 0.485 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.48 0 42.62 0.485 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.38 0 72.52 0.485 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.79 0 87.09 0.8 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.56 0 41.7 0.485 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.14 0 52.28 0.485 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.36 0 101.5 0.485 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.64 0 40.78 0.485 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.22 0 74.36 0.485 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.98 0 77.12 0.485 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.64 0 86.78 0.485 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.72 0 62.86 0.485 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.99 0 73.29 0.8 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.56 0 64.7 0.485 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.2 0 57.34 0.485 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.16 0 92.3 0.485 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.03 0 61.33 0.8 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.64 0 63.78 0.485 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.4 0 66.54 0.485 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.06 0 76.2 0.485 ;
    END
  END chany_bottom_out[20]
  PIN chany_bottom_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.3 0 73.44 0.485 ;
    END
  END chany_bottom_out[21]
  PIN chany_bottom_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.8 0 84.94 0.485 ;
    END
  END chany_bottom_out[22]
  PIN chany_bottom_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.8 0 61.94 0.485 ;
    END
  END chany_bottom_out[23]
  PIN chany_bottom_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 0 56.42 0.485 ;
    END
  END chany_bottom_out[24]
  PIN chany_bottom_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.32 0 67.46 0.485 ;
    END
  END chany_bottom_out[25]
  PIN chany_bottom_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.48 0 88.62 0.485 ;
    END
  END chany_bottom_out[26]
  PIN chany_bottom_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.2 0 80.34 0.485 ;
    END
  END chany_bottom_out[27]
  PIN chany_bottom_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.9 0 78.04 0.485 ;
    END
  END chany_bottom_out[28]
  PIN chany_bottom_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.32 0 90.46 0.485 ;
    END
  END chany_bottom_out[29]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 31.04 0.595 31.18 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 28.07 0.8 28.37 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 39.54 0.595 39.68 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 36.82 0.595 36.96 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 25.94 0.595 26.08 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 32.15 0.8 32.45 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 38.86 0.595 39 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 26.71 0.8 27.01 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 34.44 0.595 34.58 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 44.3 0.595 44.44 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.51 0.8 33.81 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.43 0.8 29.73 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 31.72 0.595 31.86 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 76.94 0.595 77.08 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.35 0.8 25.65 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 41.58 0.595 41.72 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.63 0.8 56.93 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 42.26 0.595 42.4 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 28.32 0.595 28.46 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 83.06 0.595 83.2 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 36.14 0.595 36.28 ;
    END
  END chanx_left_out[20]
  PIN chanx_left_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.59 0.8 37.89 ;
    END
  END chanx_left_out[21]
  PIN chanx_left_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 25.26 0.595 25.4 ;
    END
  END chanx_left_out[22]
  PIN chanx_left_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 74.22 0.595 74.36 ;
    END
  END chanx_left_out[23]
  PIN chanx_left_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 68.78 0.595 68.92 ;
    END
  END chanx_left_out[24]
  PIN chanx_left_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 55.27 0.8 55.57 ;
    END
  END chanx_left_out[25]
  PIN chanx_left_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 38.95 0.8 39.25 ;
    END
  END chanx_left_out[26]
  PIN chanx_left_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 34.87 0.8 35.17 ;
    END
  END chanx_left_out[27]
  PIN chanx_left_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 33.76 0.595 33.9 ;
    END
  END chanx_left_out[28]
  PIN chanx_left_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 22.54 0.595 22.68 ;
    END
  END chanx_left_out[29]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 56.2 0.595 56.34 ;
    END
  END ccff_tail[0]
  PIN Test_en_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.12 0 81.26 0.485 ;
    END
  END Test_en_S_in
  PIN Test_en_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.96 97.435 83.1 97.92 ;
    END
  END Test_en_N_out
  PIN pReset_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.88 0 61.02 0.485 ;
    END
  END pReset_S_in
  PIN pReset_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 15.4 134.32 15.54 ;
    END
  END pReset_E_in
  PIN pReset_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.63 0.8 22.93 ;
    END
  END pReset_W_in
  PIN pReset_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.66 97.435 34.8 97.92 ;
    END
  END pReset_N_out
  PIN pReset_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 20.16 0.595 20.3 ;
    END
  END pReset_W_out
  PIN pReset_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 47.02 134.32 47.16 ;
    END
  END pReset_E_out
  PIN Reset_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.04 0 82.18 0.485 ;
    END
  END Reset_S_in
  PIN Reset_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.68 97.435 74.82 97.92 ;
    END
  END Reset_N_out
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 33.74 97.435 33.88 97.92 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_1_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71 97.435 71.14 97.92 ;
    END
  END prog_clk_1_N_in
  PIN prog_clk_1_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.46 0 71.6 0.485 ;
    END
  END prog_clk_1_S_in
  PIN prog_clk_1_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 22.63 134.32 22.93 ;
    END
  END prog_clk_1_E_out
  PIN prog_clk_1_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 23.99 0.8 24.29 ;
    END
  END prog_clk_1_W_out
  PIN prog_clk_2_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.76 97.435 96.9 97.92 ;
    END
  END prog_clk_2_N_in
  PIN prog_clk_2_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 60.96 134.32 61.1 ;
    END
  END prog_clk_2_E_in
  PIN prog_clk_2_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.91 0 97.21 0.8 ;
    END
  END prog_clk_2_S_in
  PIN prog_clk_2_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 58.24 0.595 58.38 ;
    END
  END prog_clk_2_W_in
  PIN prog_clk_2_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 60.96 0.595 61.1 ;
    END
  END prog_clk_2_W_out
  PIN prog_clk_2_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.92 0 95.06 0.485 ;
    END
  END prog_clk_2_S_out
  PIN prog_clk_2_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.84 97.435 95.98 97.92 ;
    END
  END prog_clk_2_N_out
  PIN prog_clk_2_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 58.24 134.32 58.38 ;
    END
  END prog_clk_2_E_out
  PIN prog_clk_3_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 58.92 0.595 59.06 ;
    END
  END prog_clk_3_W_in
  PIN prog_clk_3_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 61.64 134.32 61.78 ;
    END
  END prog_clk_3_E_in
  PIN prog_clk_3_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.76 0 96.9 0.485 ;
    END
  END prog_clk_3_S_in
  PIN prog_clk_3_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.91 97.12 97.21 97.92 ;
    END
  END prog_clk_3_N_in
  PIN prog_clk_3_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 58.92 134.32 59.06 ;
    END
  END prog_clk_3_E_out
  PIN prog_clk_3_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 61.64 0.595 61.78 ;
    END
  END prog_clk_3_W_out
  PIN prog_clk_3_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.78 97.435 90.92 97.92 ;
    END
  END prog_clk_3_N_out
  PIN prog_clk_3_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.84 0 95.98 0.485 ;
    END
  END prog_clk_3_S_out
  PIN clk_1_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.16 97.435 92.3 97.92 ;
    END
  END clk_1_N_in
  PIN clk_1_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.54 0 70.68 0.485 ;
    END
  END clk_1_S_in
  PIN clk_1_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 23.99 134.32 24.29 ;
    END
  END clk_1_E_out
  PIN clk_1_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 23.56 0.595 23.7 ;
    END
  END clk_1_W_out
  PIN clk_2_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 87.71 97.12 88.01 97.92 ;
    END
  END clk_2_N_in
  PIN clk_2_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 63.68 134.32 63.82 ;
    END
  END clk_2_E_in
  PIN clk_2_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.96 0 83.1 0.485 ;
    END
  END clk_2_S_in
  PIN clk_2_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 64.36 0.595 64.5 ;
    END
  END clk_2_W_in
  PIN clk_2_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 63.68 0.595 63.82 ;
    END
  END clk_2_W_out
  PIN clk_2_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.68 0 97.82 0.485 ;
    END
  END clk_2_S_out
  PIN clk_2_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.68 97.435 97.82 97.92 ;
    END
  END clk_2_N_out
  PIN clk_2_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 66.06 134.32 66.2 ;
    END
  END clk_2_E_out
  PIN clk_3_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 66.06 0.595 66.2 ;
    END
  END clk_3_W_in
  PIN clk_3_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 66.74 134.32 66.88 ;
    END
  END clk_3_E_in
  PIN clk_3_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.11 0 83.41 0.8 ;
    END
  END clk_3_S_in
  PIN clk_3_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.48 97.435 88.62 97.92 ;
    END
  END clk_3_N_in
  PIN clk_3_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 64.36 134.32 64.5 ;
    END
  END clk_3_E_out
  PIN clk_3_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 66.74 0.595 66.88 ;
    END
  END clk_3_W_out
  PIN clk_3_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.6 97.435 98.74 97.92 ;
    END
  END clk_3_N_out
  PIN clk_3_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.6 0 98.74 0.485 ;
    END
  END clk_3_S_out
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 26.96 3.2 30.16 ;
        RECT 131.12 26.96 134.32 30.16 ;
        RECT 0 67.76 3.2 70.96 ;
        RECT 131.12 67.76 134.32 70.96 ;
      LAYER met4 ;
        RECT 44.78 0 45.38 0.6 ;
        RECT 74.22 0 74.82 0.6 ;
        RECT 13.5 10.88 14.1 11.48 ;
        RECT 120.22 10.88 120.82 11.48 ;
        RECT 13.5 86.44 14.1 87.04 ;
        RECT 120.22 86.44 120.82 87.04 ;
        RECT 44.78 97.32 45.38 97.92 ;
        RECT 74.22 97.32 74.82 97.92 ;
      LAYER met1 ;
        RECT 30.36 2.48 30.84 2.96 ;
        RECT 103.48 2.48 103.96 2.96 ;
        RECT 30.36 7.92 30.84 8.4 ;
        RECT 103.48 7.92 103.96 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 133.84 13.36 134.32 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 133.84 18.8 134.32 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 133.84 24.24 134.32 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 133.84 29.68 134.32 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 133.84 35.12 134.32 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 133.84 40.56 134.32 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 133.84 46 134.32 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 133.84 51.44 134.32 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 133.84 56.88 134.32 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 133.84 62.32 134.32 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 133.84 67.76 134.32 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 133.84 73.2 134.32 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 133.84 78.64 134.32 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 133.84 84.08 134.32 84.56 ;
        RECT 30.36 89.52 30.84 90 ;
        RECT 103.48 89.52 103.96 90 ;
        RECT 30.36 94.96 30.84 95.44 ;
        RECT 103.48 94.96 103.96 95.44 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 47.36 3.2 50.56 ;
        RECT 131.12 47.36 134.32 50.56 ;
      LAYER met4 ;
        RECT 59.5 0 60.1 0.6 ;
        RECT 88.94 0 89.54 0.6 ;
        RECT 59.5 97.32 60.1 97.92 ;
        RECT 88.94 97.32 89.54 97.92 ;
      LAYER met1 ;
        RECT 30.36 -0.24 30.84 0.24 ;
        RECT 103.48 -0.24 103.96 0.24 ;
        RECT 30.36 5.2 30.84 5.68 ;
        RECT 103.48 5.2 103.96 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 133.84 10.64 134.32 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 133.84 16.08 134.32 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 133.84 21.52 134.32 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 133.84 26.96 134.32 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 133.84 32.4 134.32 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 133.84 37.84 134.32 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 133.84 43.28 134.32 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 133.84 48.72 134.32 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 133.84 54.16 134.32 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 133.84 59.6 134.32 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 133.84 65.04 134.32 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 133.84 70.48 134.32 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 133.84 75.92 134.32 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 133.84 81.36 134.32 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 133.84 86.8 134.32 87.28 ;
        RECT 30.36 92.24 30.84 92.72 ;
        RECT 103.48 92.24 103.96 92.72 ;
        RECT 30.36 97.68 30.84 98.16 ;
        RECT 103.48 97.68 103.96 98.16 ;
    END
  END VSS
  OBS
    LAYER met2 ;
      RECT 89.1 97.615 89.38 97.985 ;
      RECT 59.66 97.615 59.94 97.985 ;
      POLYGON 75.28 97.82 75.28 93.26 75.14 93.26 75.14 97.68 75.1 97.68 75.1 97.82 ;
      POLYGON 31.65 97.765 31.65 97.395 31.58 97.395 31.58 87.31 31.44 87.31 31.44 97.395 31.37 97.395 31.37 97.765 ;
      RECT 98.08 96.91 98.34 97.23 ;
      RECT 72.32 96.91 72.58 97.23 ;
      RECT 41.96 96.91 42.22 97.23 ;
      POLYGON 125.95 86.885 125.95 86.515 125.88 86.515 125.88 83.91 125.74 83.91 125.74 86.515 125.67 86.515 125.67 86.885 ;
      POLYGON 26.59 86.885 26.59 86.515 26.52 86.515 26.52 71.67 26.38 71.67 26.38 86.515 26.31 86.515 26.31 86.885 ;
      POLYGON 16.01 86.885 16.01 86.515 15.94 86.515 15.94 78.3 15.8 78.3 15.8 86.515 15.73 86.515 15.73 86.885 ;
      RECT 17.12 86.03 17.38 86.35 ;
      POLYGON 24.22 38.66 24.22 11.405 24.29 11.405 24.29 11.035 24.01 11.035 24.01 11.405 24.08 11.405 24.08 38.66 ;
      POLYGON 73.9 17.24 73.9 0.24 73.94 0.24 73.94 0.1 73.76 0.1 73.76 17.24 ;
      POLYGON 82.64 15.88 82.64 0.24 82.68 0.24 82.68 0.1 82.5 0.1 82.5 15.88 ;
      POLYGON 30.66 15.37 30.66 1.77 31.58 1.77 31.58 1.63 30.52 1.63 30.52 15.37 ;
      POLYGON 103.8 11.46 103.8 5.71 102.28 5.71 102.28 5.85 103.66 5.85 103.66 11.46 ;
      RECT 89.8 0.69 90.06 1.01 ;
      RECT 56.68 0.69 56.94 1.01 ;
      RECT 41.93 0.72 42.25 0.98 ;
      RECT 64.96 0.35 65.22 0.67 ;
      RECT 89.1 -0.065 89.38 0.305 ;
      RECT 59.66 -0.065 59.94 0.305 ;
      RECT 96.26 0 96.48 0.14 ;
      POLYGON 103.68 97.64 103.68 86.76 134.04 86.76 134.04 11.16 125.24 11.16 125.24 11.645 124.54 11.645 124.54 11.16 124.32 11.16 124.32 11.645 123.62 11.645 123.62 11.16 121.56 11.16 121.56 11.645 120.86 11.645 120.86 11.16 103.68 11.16 103.68 0.28 101.78 0.28 101.78 0.765 101.08 0.765 101.08 0.28 100.86 0.28 100.86 0.765 100.16 0.765 100.16 0.28 99.94 0.28 99.94 0.765 99.24 0.765 99.24 0.28 99.02 0.28 99.02 0.765 98.32 0.765 98.32 0.28 98.1 0.28 98.1 0.765 97.4 0.765 97.4 0.28 97.18 0.28 97.18 0.765 96.48 0.765 96.48 0.28 96.26 0.28 96.26 0.765 95.56 0.765 95.56 0.28 95.34 0.28 95.34 0.765 94.64 0.765 94.64 0.28 94.42 0.28 94.42 0.765 93.72 0.765 93.72 0.28 93.5 0.28 93.5 0.765 92.8 0.765 92.8 0.28 92.58 0.28 92.58 0.765 91.88 0.765 91.88 0.28 91.66 0.28 91.66 0.765 90.96 0.765 90.96 0.28 90.74 0.28 90.74 0.765 90.04 0.765 90.04 0.28 88.9 0.28 88.9 0.765 88.2 0.765 88.2 0.28 87.98 0.28 87.98 0.765 87.28 0.765 87.28 0.28 87.06 0.28 87.06 0.765 86.36 0.765 86.36 0.28 86.14 0.28 86.14 0.765 85.44 0.765 85.44 0.28 85.22 0.28 85.22 0.765 84.52 0.765 84.52 0.28 84.3 0.28 84.3 0.765 83.6 0.765 83.6 0.28 83.38 0.28 83.38 0.765 82.68 0.765 82.68 0.28 82.46 0.28 82.46 0.765 81.76 0.765 81.76 0.28 81.54 0.28 81.54 0.765 80.84 0.765 80.84 0.28 80.62 0.28 80.62 0.765 79.92 0.765 79.92 0.28 79.24 0.28 79.24 0.765 78.54 0.765 78.54 0.28 78.32 0.28 78.32 0.765 77.62 0.765 77.62 0.28 77.4 0.28 77.4 0.765 76.7 0.765 76.7 0.28 76.48 0.28 76.48 0.765 75.78 0.765 75.78 0.28 75.56 0.28 75.56 0.765 74.86 0.765 74.86 0.28 74.64 0.28 74.64 0.765 73.94 0.765 73.94 0.28 73.72 0.28 73.72 0.765 73.02 0.765 73.02 0.28 72.8 0.28 72.8 0.765 72.1 0.765 72.1 0.28 71.88 0.28 71.88 0.765 71.18 0.765 71.18 0.28 70.96 0.28 70.96 0.765 70.26 0.765 70.26 0.28 69.58 0.28 69.58 0.765 68.88 0.765 68.88 0.28 68.66 0.28 68.66 0.765 67.96 0.765 67.96 0.28 67.74 0.28 67.74 0.765 67.04 0.765 67.04 0.28 66.82 0.28 66.82 0.765 66.12 0.765 66.12 0.28 65.9 0.28 65.9 0.765 65.2 0.765 65.2 0.28 64.98 0.28 64.98 0.765 64.28 0.765 64.28 0.28 64.06 0.28 64.06 0.765 63.36 0.765 63.36 0.28 63.14 0.28 63.14 0.765 62.44 0.765 62.44 0.28 62.22 0.28 62.22 0.765 61.52 0.765 61.52 0.28 61.3 0.28 61.3 0.765 60.6 0.765 60.6 0.28 59.46 0.28 59.46 0.765 58.76 0.765 58.76 0.28 58.54 0.28 58.54 0.765 57.84 0.765 57.84 0.28 57.62 0.28 57.62 0.765 56.92 0.765 56.92 0.28 56.7 0.28 56.7 0.765 56 0.765 56 0.28 55.78 0.28 55.78 0.765 55.08 0.765 55.08 0.28 52.56 0.28 52.56 0.765 51.86 0.765 51.86 0.28 46.12 0.28 46.12 0.765 45.42 0.765 45.42 0.28 45.2 0.28 45.2 0.765 44.5 0.765 44.5 0.28 42.9 0.28 42.9 0.765 42.2 0.765 42.2 0.28 41.98 0.28 41.98 0.765 41.28 0.765 41.28 0.28 41.06 0.28 41.06 0.765 40.36 0.765 40.36 0.28 30.64 0.28 30.64 11.16 20.36 11.16 20.36 11.645 19.66 11.645 19.66 11.16 18.52 11.16 18.52 11.645 17.82 11.645 17.82 11.16 17.14 11.16 17.14 11.645 16.44 11.645 16.44 11.16 16.22 11.16 16.22 11.645 15.52 11.645 15.52 11.16 15.3 11.16 15.3 11.645 14.6 11.645 14.6 11.16 14.38 11.16 14.38 11.645 13.68 11.645 13.68 11.16 13.46 11.16 13.46 11.645 12.76 11.645 12.76 11.16 12.54 11.16 12.54 11.645 11.84 11.645 11.84 11.16 11.62 11.16 11.62 11.645 10.92 11.645 10.92 11.16 10.7 11.16 10.7 11.645 10 11.645 10 11.16 9.78 11.16 9.78 11.645 9.08 11.645 9.08 11.16 8.86 11.16 8.86 11.645 8.16 11.645 8.16 11.16 7.94 11.16 7.94 11.645 7.24 11.645 7.24 11.16 7.02 11.16 7.02 11.645 6.32 11.645 6.32 11.16 0.28 11.16 0.28 86.76 9.54 86.76 9.54 86.275 10.24 86.275 10.24 86.76 13.68 86.76 13.68 86.275 14.38 86.275 14.38 86.76 17.36 86.76 17.36 86.275 18.06 86.275 18.06 86.76 18.28 86.76 18.28 86.275 18.98 86.275 18.98 86.76 30.64 86.76 30.64 97.64 33.46 97.64 33.46 97.155 34.16 97.155 34.16 97.64 34.38 97.64 34.38 97.155 35.08 97.155 35.08 97.64 36.68 97.64 36.68 97.155 37.38 97.155 37.38 97.64 37.6 97.64 37.6 97.155 38.3 97.155 38.3 97.64 40.82 97.64 40.82 97.155 41.52 97.155 41.52 97.64 42.2 97.64 42.2 97.155 42.9 97.155 42.9 97.64 44.04 97.64 44.04 97.155 44.74 97.155 44.74 97.64 46.34 97.64 46.34 97.155 47.04 97.155 47.04 97.64 47.72 97.64 47.72 97.155 48.42 97.155 48.42 97.64 48.64 97.64 48.64 97.155 49.34 97.155 49.34 97.64 51.4 97.64 51.4 97.155 52.1 97.155 52.1 97.64 57.84 97.64 57.84 97.155 58.54 97.155 58.54 97.64 58.76 97.64 58.76 97.155 59.46 97.155 59.46 97.64 60.6 97.64 60.6 97.155 61.3 97.155 61.3 97.64 61.52 97.64 61.52 97.155 62.22 97.155 62.22 97.64 62.9 97.64 62.9 97.155 63.6 97.155 63.6 97.64 63.82 97.64 63.82 97.155 64.52 97.155 64.52 97.64 64.74 97.64 64.74 97.155 65.44 97.155 65.44 97.64 65.66 97.64 65.66 97.155 66.36 97.155 66.36 97.64 66.58 97.64 66.58 97.155 67.28 97.155 67.28 97.64 67.5 97.64 67.5 97.155 68.2 97.155 68.2 97.64 68.42 97.64 68.42 97.155 69.12 97.155 69.12 97.64 69.34 97.64 69.34 97.155 70.04 97.155 70.04 97.64 70.72 97.64 70.72 97.155 71.42 97.155 71.42 97.64 71.64 97.64 71.64 97.155 72.34 97.155 72.34 97.64 73.02 97.64 73.02 97.155 73.72 97.155 73.72 97.64 74.4 97.64 74.4 97.155 75.1 97.155 75.1 97.64 75.32 97.64 75.32 97.155 76.02 97.155 76.02 97.64 76.24 97.64 76.24 97.155 76.94 97.155 76.94 97.64 77.16 97.64 77.16 97.155 77.86 97.155 77.86 97.64 78.08 97.64 78.08 97.155 78.78 97.155 78.78 97.64 79 97.64 79 97.155 79.7 97.155 79.7 97.64 79.92 97.64 79.92 97.155 80.62 97.155 80.62 97.64 80.84 97.64 80.84 97.155 81.54 97.155 81.54 97.64 81.76 97.64 81.76 97.155 82.46 97.155 82.46 97.64 82.68 97.64 82.68 97.155 83.38 97.155 83.38 97.64 83.6 97.64 83.6 97.155 84.3 97.155 84.3 97.64 84.52 97.64 84.52 97.155 85.22 97.155 85.22 97.64 85.44 97.64 85.44 97.155 86.14 97.155 86.14 97.64 86.36 97.64 86.36 97.155 87.06 97.155 87.06 97.64 87.28 97.64 87.28 97.155 87.98 97.155 87.98 97.64 88.2 97.64 88.2 97.155 88.9 97.155 88.9 97.64 89.58 97.64 89.58 97.155 90.28 97.155 90.28 97.64 90.5 97.64 90.5 97.155 91.2 97.155 91.2 97.64 91.88 97.64 91.88 97.155 92.58 97.155 92.58 97.64 92.8 97.64 92.8 97.155 93.5 97.155 93.5 97.64 93.72 97.64 93.72 97.155 94.42 97.155 94.42 97.64 94.64 97.64 94.64 97.155 95.34 97.155 95.34 97.64 95.56 97.64 95.56 97.155 96.26 97.155 96.26 97.64 96.48 97.64 96.48 97.155 97.18 97.155 97.18 97.64 97.4 97.64 97.4 97.155 98.1 97.155 98.1 97.64 98.32 97.64 98.32 97.155 99.02 97.155 99.02 97.64 99.24 97.64 99.24 97.155 99.94 97.155 99.94 97.64 100.16 97.64 100.16 97.155 100.86 97.155 100.86 97.64 101.08 97.64 101.08 97.155 101.78 97.155 101.78 97.64 ;
    LAYER met4 ;
      POLYGON 87.105 97.745 87.105 97.415 87.09 97.415 87.09 48.47 86.79 48.47 86.79 97.415 86.775 97.415 86.775 97.745 ;
      POLYGON 65.945 97.745 65.945 97.415 65.93 97.415 65.93 70.06 65.63 70.06 65.63 97.415 65.615 97.415 65.615 97.745 ;
      POLYGON 50.305 97.745 50.305 97.415 50.29 97.415 50.29 95.39 49.99 95.39 49.99 97.415 49.975 97.415 49.975 97.745 ;
      POLYGON 64.09 97.73 64.09 43.03 63.79 43.03 63.79 97.43 63.57 97.43 63.57 97.73 ;
      POLYGON 31.89 95.69 31.89 95.39 30.97 95.39 30.97 77.71 30.67 77.71 30.67 95.69 ;
      POLYGON 103.65 94.33 103.65 85.19 103.35 85.19 103.35 94.03 102.43 94.03 102.43 94.33 ;
      POLYGON 64.09 41.29 64.09 0.505 64.105 0.505 64.105 0.175 63.775 0.175 63.775 0.505 63.79 0.505 63.79 41.29 ;
      POLYGON 103.56 97.52 103.56 86.64 119.82 86.64 119.82 86.04 121.22 86.04 121.22 86.64 133.92 86.64 133.92 11.28 121.22 11.28 121.22 11.88 119.82 11.88 119.82 11.28 103.56 11.28 103.56 0.4 99.45 0.4 99.45 1.2 98.35 1.2 98.35 0.4 97.61 0.4 97.61 1.2 96.51 1.2 96.51 0.4 94.85 0.4 94.85 1.2 93.75 1.2 93.75 0.4 93.01 0.4 93.01 1.2 91.91 1.2 91.91 0.4 91.17 0.4 91.17 1.2 90.07 1.2 90.07 0.4 89.94 0.4 89.94 1 88.54 1 88.54 0.4 87.49 0.4 87.49 1.2 86.39 1.2 86.39 0.4 85.65 0.4 85.65 1.2 84.55 1.2 84.55 0.4 83.81 0.4 83.81 1.2 82.71 1.2 82.71 0.4 81.05 0.4 81.05 1.2 79.95 1.2 79.95 0.4 79.21 0.4 79.21 1.2 78.11 1.2 78.11 0.4 77.37 0.4 77.37 1.2 76.27 1.2 76.27 0.4 75.22 0.4 75.22 1 73.82 1 73.82 0.4 73.69 0.4 73.69 1.2 72.59 1.2 72.59 0.4 71.85 0.4 71.85 1.2 70.75 1.2 70.75 0.4 69.09 0.4 69.09 1.2 67.99 1.2 67.99 0.4 67.25 0.4 67.25 1.2 66.15 1.2 66.15 0.4 65.41 0.4 65.41 1.2 64.31 1.2 64.31 0.4 63.57 0.4 63.57 1.2 62.47 1.2 62.47 0.4 61.73 0.4 61.73 1.2 60.63 1.2 60.63 0.4 60.5 0.4 60.5 1 59.1 1 59.1 0.4 58.97 0.4 58.97 1.2 57.87 1.2 57.87 0.4 45.78 0.4 45.78 1 44.38 1 44.38 0.4 30.76 0.4 30.76 11.28 14.5 11.28 14.5 11.88 13.1 11.88 13.1 11.28 0.4 11.28 0.4 86.64 13.1 86.64 13.1 86.04 14.5 86.04 14.5 86.64 30.76 86.64 30.76 97.52 44.38 97.52 44.38 96.92 45.78 96.92 45.78 97.52 57.87 97.52 57.87 96.72 58.97 96.72 58.97 97.52 59.1 97.52 59.1 96.92 60.5 96.92 60.5 97.52 60.63 97.52 60.63 96.72 61.73 96.72 61.73 97.52 62.47 97.52 62.47 96.72 63.57 96.72 63.57 97.52 64.31 97.52 64.31 96.72 65.41 96.72 65.41 97.52 66.15 97.52 66.15 96.72 67.25 96.72 67.25 97.52 67.99 97.52 67.99 96.72 69.09 96.72 69.09 97.52 69.83 97.52 69.83 96.72 70.93 96.72 70.93 97.52 71.67 97.52 71.67 96.72 72.77 96.72 72.77 97.52 73.82 97.52 73.82 96.92 75.22 96.92 75.22 97.52 76.27 97.52 76.27 96.72 77.37 96.72 77.37 97.52 78.11 97.52 78.11 96.72 79.21 96.72 79.21 97.52 79.95 97.52 79.95 96.72 81.05 96.72 81.05 97.52 81.79 97.52 81.79 96.72 82.89 96.72 82.89 97.52 83.63 97.52 83.63 96.72 84.73 96.72 84.73 97.52 85.47 97.52 85.47 96.72 86.57 96.72 86.57 97.52 87.31 97.52 87.31 96.72 88.41 96.72 88.41 97.52 88.54 97.52 88.54 96.92 89.94 96.92 89.94 97.52 90.07 97.52 90.07 96.72 91.17 96.72 91.17 97.52 91.91 97.52 91.91 96.72 93.01 96.72 93.01 97.52 93.75 97.52 93.75 96.72 94.85 96.72 94.85 97.52 96.51 97.52 96.51 96.72 97.61 96.72 97.61 97.52 98.35 97.52 98.35 96.72 99.45 96.72 99.45 97.52 ;
    LAYER met1 ;
      POLYGON 103.2 98.16 103.2 97.68 89.4 97.68 89.4 97.67 89.08 97.67 89.08 97.68 59.96 97.68 59.96 97.67 59.64 97.67 59.64 97.68 31.12 97.68 31.12 98.16 ;
      POLYGON 37.1 90.68 37.1 90.54 30.52 90.54 30.52 90.6 31.235 90.6 31.235 90.68 ;
      RECT 72.36 86.8 133.56 87.28 ;
      RECT 0.76 86.8 71.16 87.28 ;
      POLYGON 3.98 48.52 3.98 48.38 0.76 48.38 0.76 48.12 0.62 48.12 0.62 48.52 ;
      POLYGON 133.795 37.64 133.795 37.24 133.655 37.24 133.655 37.5 128.5 37.5 128.5 37.64 ;
      RECT 72.36 10.64 133.56 11.12 ;
      RECT 0.76 10.64 71.16 11.12 ;
      POLYGON 89.4 0.25 89.4 0.24 103.2 0.24 103.2 -0.24 31.12 -0.24 31.12 0.24 59.64 0.24 59.64 0.25 59.96 0.25 59.96 0.24 89.08 0.24 89.08 0.25 ;
      POLYGON 103.2 97.64 103.2 97.4 103.68 97.4 103.68 95.72 103.2 95.72 103.2 94.68 103.68 94.68 103.68 93 103.2 93 103.2 91.96 103.68 91.96 103.68 90.28 103.2 90.28 103.2 89.24 103.68 89.24 103.68 86.76 133.56 86.76 133.56 86.52 134.04 86.52 134.04 84.84 133.56 84.84 133.56 83.8 134.04 83.8 134.04 82.12 133.56 82.12 133.56 81.08 134.04 81.08 134.04 80.08 133.445 80.08 133.445 79.38 133.56 79.38 133.56 78.36 134.04 78.36 134.04 78.04 133.445 78.04 133.445 76.66 133.56 76.66 133.56 75.64 134.04 75.64 134.04 75.32 133.445 75.32 133.445 73.94 133.56 73.94 133.56 72.92 134.04 72.92 134.04 72.6 133.445 72.6 133.445 71.22 133.56 71.22 133.56 70.2 134.04 70.2 134.04 69.88 133.445 69.88 133.445 68.5 133.56 68.5 133.56 67.48 134.04 67.48 134.04 67.16 133.445 67.16 133.445 65.78 133.56 65.78 133.56 64.78 133.445 64.78 133.445 63.4 134.04 63.4 134.04 63.08 133.56 63.08 133.56 62.06 133.445 62.06 133.445 60.68 134.04 60.68 134.04 60.36 133.56 60.36 133.56 59.34 133.445 59.34 133.445 57.96 134.04 57.96 134.04 57.64 133.56 57.64 133.56 56.62 133.445 56.62 133.445 55.24 134.04 55.24 134.04 54.92 133.56 54.92 133.56 53.88 134.04 53.88 134.04 53.56 133.445 53.56 133.445 52.18 133.56 52.18 133.56 51.16 134.04 51.16 134.04 50.84 133.445 50.84 133.445 49.46 133.56 49.46 133.56 48.44 134.04 48.44 134.04 48.12 133.445 48.12 133.445 46.74 133.56 46.74 133.56 45.72 134.04 45.72 134.04 44.72 133.445 44.72 133.445 44.02 133.56 44.02 133.56 43 134.04 43 134.04 42.68 133.445 42.68 133.445 41.3 133.56 41.3 133.56 40.28 134.04 40.28 134.04 39.96 133.445 39.96 133.445 38.58 133.56 38.58 133.56 37.56 134.04 37.56 134.04 37.24 133.445 37.24 133.445 35.86 133.56 35.86 133.56 34.86 133.445 34.86 133.445 33.48 134.04 33.48 134.04 33.16 133.56 33.16 133.56 32.14 133.445 32.14 133.445 30.76 134.04 30.76 134.04 30.44 133.56 30.44 133.56 29.42 133.445 29.42 133.445 28.72 134.04 28.72 134.04 28.4 133.445 28.4 133.445 27.7 133.56 27.7 133.56 26.68 134.04 26.68 134.04 26.36 133.445 26.36 133.445 24.98 133.56 24.98 133.56 23.96 134.04 23.96 134.04 23.64 133.445 23.64 133.445 22.26 133.56 22.26 133.56 21.24 134.04 21.24 134.04 19.56 133.56 19.56 133.56 18.52 134.04 18.52 134.04 16.84 133.56 16.84 133.56 15.82 133.445 15.82 133.445 15.12 134.04 15.12 134.04 14.8 133.445 14.8 133.445 14.1 133.56 14.1 133.56 13.1 133.445 13.1 133.445 12.4 134.04 12.4 134.04 11.4 133.56 11.4 133.56 11.16 103.68 11.16 103.68 8.68 103.2 8.68 103.2 7.64 103.68 7.64 103.68 7.32 103.085 7.32 103.085 5.94 103.2 5.94 103.2 4.92 103.68 4.92 103.68 3.24 103.2 3.24 103.2 2.22 103.085 2.22 103.085 1.52 103.68 1.52 103.68 0.52 103.2 0.52 103.2 0.28 31.12 0.28 31.12 0.52 30.64 0.52 30.64 2.2 31.12 2.2 31.12 3.24 30.64 3.24 30.64 4.92 31.12 4.92 31.12 5.94 31.235 5.94 31.235 6.64 30.64 6.64 30.64 7.64 31.12 7.64 31.12 8.68 30.64 8.68 30.64 11.16 0.76 11.16 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 19.88 0.875 19.88 0.875 20.58 0.28 20.58 0.28 21.24 0.76 21.24 0.76 22.26 0.875 22.26 0.875 22.96 0.28 22.96 0.28 23.28 0.875 23.28 0.875 23.98 0.76 23.98 0.76 24.98 0.875 24.98 0.875 26.36 0.28 26.36 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 28.04 0.875 28.04 0.875 29.42 0.76 29.42 0.76 30.44 0.28 30.44 0.28 30.76 0.875 30.76 0.875 32.14 0.76 32.14 0.76 33.16 0.28 33.16 0.28 33.48 0.875 33.48 0.875 34.86 0.76 34.86 0.76 35.86 0.875 35.86 0.875 37.24 0.28 37.24 0.28 37.56 0.76 37.56 0.76 38.58 0.875 38.58 0.875 39.96 0.28 39.96 0.28 40.28 0.76 40.28 0.76 41.3 0.875 41.3 0.875 42.68 0.28 42.68 0.28 43 0.76 43 0.76 44.02 0.875 44.02 0.875 45.4 0.28 45.4 0.28 45.72 0.76 45.72 0.76 46.74 0.875 46.74 0.875 48.12 0.28 48.12 0.28 48.44 0.76 48.44 0.76 49.46 0.875 49.46 0.875 50.84 0.28 50.84 0.28 51.16 0.76 51.16 0.76 52.18 0.875 52.18 0.875 53.56 0.28 53.56 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 55.24 0.875 55.24 0.875 56.62 0.76 56.62 0.76 57.64 0.28 57.64 0.28 57.96 0.875 57.96 0.875 59.34 0.76 59.34 0.76 60.36 0.28 60.36 0.28 60.68 0.875 60.68 0.875 62.06 0.76 62.06 0.76 63.08 0.28 63.08 0.28 63.4 0.875 63.4 0.875 64.78 0.76 64.78 0.76 65.78 0.875 65.78 0.875 67.16 0.28 67.16 0.28 67.48 0.76 67.48 0.76 68.5 0.875 68.5 0.875 69.88 0.28 69.88 0.28 70.2 0.76 70.2 0.76 71.22 0.875 71.22 0.875 72.6 0.28 72.6 0.28 72.92 0.76 72.92 0.76 73.94 0.875 73.94 0.875 75.32 0.28 75.32 0.28 75.64 0.76 75.64 0.76 76.66 0.875 76.66 0.875 78.04 0.28 78.04 0.28 78.36 0.76 78.36 0.76 79.38 0.875 79.38 0.875 80.76 0.28 80.76 0.28 81.08 0.76 81.08 0.76 82.1 0.875 82.1 0.875 83.48 0.28 83.48 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 86.76 30.64 86.76 30.64 88.56 31.235 88.56 31.235 89.26 31.12 89.26 31.12 90.28 30.64 90.28 30.64 90.6 31.235 90.6 31.235 91.98 31.12 91.98 31.12 93 30.64 93 30.64 94.68 31.12 94.68 31.12 95.72 30.64 95.72 30.64 97.4 31.12 97.4 31.12 97.64 ;
    LAYER met3 ;
      POLYGON 89.405 97.965 89.405 97.96 89.62 97.96 89.62 97.64 89.405 97.64 89.405 97.635 89.075 97.635 89.075 97.64 88.86 97.64 88.86 97.96 89.075 97.96 89.075 97.965 ;
      POLYGON 59.965 97.965 59.965 97.96 60.18 97.96 60.18 97.64 59.965 97.64 59.965 97.635 59.635 97.635 59.635 97.64 59.42 97.64 59.42 97.96 59.635 97.96 59.635 97.965 ;
      POLYGON 96.995 97.745 96.995 97.415 96.665 97.415 96.665 97.43 96.075 97.43 96.075 97.415 95.745 97.415 95.745 97.745 96.075 97.745 96.075 97.73 96.665 97.73 96.665 97.745 ;
      POLYGON 31.675 97.745 31.675 97.73 49.95 97.73 49.95 97.74 50.33 97.74 50.33 97.42 49.95 97.42 49.95 97.43 31.675 97.43 31.675 97.415 31.345 97.415 31.345 97.745 ;
      POLYGON 87.13 97.74 87.13 97.42 86.75 97.42 86.75 97.43 70.57 97.43 70.57 97.42 70.19 97.42 70.19 97.74 70.57 97.74 70.57 97.73 86.75 97.73 86.75 97.74 ;
      POLYGON 65.97 97.74 65.97 97.42 65.59 97.42 65.59 97.43 61.37 97.43 61.37 97.42 60.99 97.42 60.99 97.74 61.37 97.74 61.37 97.73 65.59 97.73 65.59 97.74 ;
      RECT 31.55 91.3 31.93 91.62 ;
      POLYGON 125.975 86.865 125.975 86.535 125.645 86.535 125.645 86.55 90.24 86.55 90.24 86.85 125.645 86.85 125.645 86.865 ;
      POLYGON 26.615 86.865 26.615 86.85 31.66 86.85 31.66 86.55 26.615 86.55 26.615 86.535 26.285 86.535 26.285 86.865 ;
      POLYGON 16.035 86.865 16.035 86.535 15.705 86.535 15.705 86.55 14.195 86.55 14.195 86.535 13.865 86.535 13.865 86.865 14.195 86.865 14.195 86.85 15.705 86.85 15.705 86.865 ;
      POLYGON 133.12 34.49 133.12 34.47 133.67 34.47 133.67 34.19 114.62 34.19 114.62 34.49 ;
      POLYGON 1.315 26.345 1.315 26.34 1.57 26.34 1.57 26.02 1.315 26.02 1.315 26.015 0.985 26.015 0.985 26.02 0.615 26.02 0.615 26.34 0.985 26.34 0.985 26.345 ;
      POLYGON 133.67 26.33 133.67 26.05 133.12 26.05 133.12 26.03 110.94 26.03 110.94 26.33 ;
      POLYGON 1.315 24.985 1.315 24.97 12.34 24.97 12.34 24.67 1.315 24.67 1.315 24.655 0.985 24.655 0.985 24.985 ;
      POLYGON 114 12.05 114 11.07 102.2 11.07 102.2 11.37 113.7 11.37 113.7 12.05 ;
      POLYGON 24.315 11.385 24.315 11.37 48.22 11.37 48.22 11.07 24.315 11.07 24.315 11.055 23.985 11.055 23.985 11.07 18.335 11.07 18.335 11.055 18.005 11.055 18.005 11.385 18.335 11.385 18.335 11.37 23.985 11.37 23.985 11.385 ;
      RECT 31.55 6.3 31.93 6.62 ;
      POLYGON 31.675 5.265 31.675 5.25 51.44 5.25 51.44 4.95 31.675 4.95 31.675 4.935 31.345 4.935 31.345 5.265 ;
      POLYGON 65.01 1.85 65.01 0.5 65.05 0.5 65.05 0.18 64.67 0.18 64.67 0.5 64.71 0.5 64.71 1.85 ;
      POLYGON 62.955 0.505 62.955 0.49 63.75 0.49 63.75 0.5 64.13 0.5 64.13 0.18 63.75 0.18 63.75 0.19 62.955 0.19 62.955 0.175 62.625 0.175 62.625 0.505 ;
      POLYGON 89.405 0.285 89.405 0.28 89.62 0.28 89.62 -0.04 89.405 -0.04 89.405 -0.045 89.075 -0.045 89.075 -0.04 88.86 -0.04 88.86 0.28 89.075 0.28 89.075 0.285 ;
      POLYGON 59.965 0.285 59.965 0.28 60.18 0.28 60.18 -0.04 59.965 -0.04 59.965 -0.045 59.635 -0.045 59.635 -0.04 59.42 -0.04 59.42 0.28 59.635 0.28 59.635 0.285 ;
      POLYGON 103.56 97.52 103.56 86.64 133.92 86.64 133.92 62.77 133.12 62.77 133.12 61.67 133.92 61.67 133.92 61.41 133.12 61.41 133.12 60.31 133.92 60.31 133.92 60.05 133.12 60.05 133.12 58.95 133.92 58.95 133.92 58.69 133.12 58.69 133.12 57.59 133.92 57.59 133.92 57.33 133.12 57.33 133.12 56.23 133.92 56.23 133.92 55.97 133.12 55.97 133.12 54.87 133.92 54.87 133.92 54.61 133.12 54.61 133.12 53.51 133.92 53.51 133.92 53.25 133.12 53.25 133.12 52.15 133.92 52.15 133.92 51.89 133.12 51.89 133.12 50.79 133.92 50.79 133.92 50.53 133.12 50.53 133.12 49.43 133.92 49.43 133.92 49.17 133.12 49.17 133.12 48.07 133.92 48.07 133.92 47.81 133.12 47.81 133.12 46.71 133.92 46.71 133.92 46.45 133.12 46.45 133.12 45.35 133.92 45.35 133.92 45.09 133.12 45.09 133.12 43.99 133.92 43.99 133.92 43.73 133.12 43.73 133.12 42.63 133.92 42.63 133.92 42.37 133.12 42.37 133.12 41.27 133.92 41.27 133.92 41.01 133.12 41.01 133.12 39.91 133.92 39.91 133.92 39.65 133.12 39.65 133.12 38.55 133.92 38.55 133.92 38.29 133.12 38.29 133.12 37.19 133.92 37.19 133.92 36.93 133.12 36.93 133.12 35.83 133.92 35.83 133.92 35.57 133.12 35.57 133.12 34.47 133.92 34.47 133.92 34.21 133.12 34.21 133.12 33.11 133.92 33.11 133.92 32.85 133.12 32.85 133.12 31.75 133.92 31.75 133.92 31.49 133.12 31.49 133.12 30.39 133.92 30.39 133.92 30.13 133.12 30.13 133.12 29.03 133.92 29.03 133.92 28.77 133.12 28.77 133.12 27.67 133.92 27.67 133.92 27.41 133.12 27.41 133.12 26.31 133.92 26.31 133.92 26.05 133.12 26.05 133.12 24.95 133.92 24.95 133.92 24.69 133.12 24.69 133.12 23.59 133.92 23.59 133.92 23.33 133.12 23.33 133.12 22.23 133.92 22.23 133.92 11.28 103.56 11.28 103.56 0.4 30.76 0.4 30.76 5.23 31.56 5.23 31.56 6.33 30.76 6.33 30.76 11.28 0.4 11.28 0.4 22.23 1.2 22.23 1.2 23.33 0.4 23.33 0.4 23.59 1.2 23.59 1.2 24.69 0.4 24.69 0.4 24.95 1.2 24.95 1.2 26.05 0.4 26.05 0.4 26.31 1.2 26.31 1.2 27.41 0.4 27.41 0.4 27.67 1.2 27.67 1.2 28.77 0.4 28.77 0.4 29.03 1.2 29.03 1.2 30.13 0.4 30.13 0.4 30.39 1.2 30.39 1.2 31.49 0.4 31.49 0.4 31.75 1.2 31.75 1.2 32.85 0.4 32.85 0.4 33.11 1.2 33.11 1.2 34.21 0.4 34.21 0.4 34.47 1.2 34.47 1.2 35.57 0.4 35.57 0.4 35.83 1.2 35.83 1.2 36.93 0.4 36.93 0.4 37.19 1.2 37.19 1.2 38.29 0.4 38.29 0.4 38.55 1.2 38.55 1.2 39.65 0.4 39.65 0.4 39.91 1.2 39.91 1.2 41.01 0.4 41.01 0.4 41.27 1.2 41.27 1.2 42.37 0.4 42.37 0.4 42.63 1.2 42.63 1.2 43.73 0.4 43.73 0.4 43.99 1.2 43.99 1.2 45.09 0.4 45.09 0.4 45.35 1.2 45.35 1.2 46.45 0.4 46.45 0.4 46.71 1.2 46.71 1.2 47.81 0.4 47.81 0.4 48.07 1.2 48.07 1.2 49.17 0.4 49.17 0.4 49.43 1.2 49.43 1.2 50.53 0.4 50.53 0.4 50.79 1.2 50.79 1.2 51.89 0.4 51.89 0.4 52.15 1.2 52.15 1.2 53.25 0.4 53.25 0.4 53.51 1.2 53.51 1.2 54.61 0.4 54.61 0.4 54.87 1.2 54.87 1.2 55.97 0.4 55.97 0.4 56.23 1.2 56.23 1.2 57.33 0.4 57.33 0.4 86.64 30.76 86.64 30.76 91.59 31.56 91.59 31.56 92.69 30.76 92.69 30.76 97.52 ;
    LAYER met5 ;
      POLYGON 102.36 96.32 102.36 85.44 132.72 85.44 132.72 72.56 129.52 72.56 129.52 66.16 132.72 66.16 132.72 52.16 129.52 52.16 129.52 45.76 132.72 45.76 132.72 31.76 129.52 31.76 129.52 25.36 132.72 25.36 132.72 12.48 102.36 12.48 102.36 1.6 31.96 1.6 31.96 12.48 1.6 12.48 1.6 25.36 4.8 25.36 4.8 31.76 1.6 31.76 1.6 45.76 4.8 45.76 4.8 52.16 1.6 52.16 1.6 66.16 4.8 66.16 4.8 72.56 1.6 72.56 1.6 85.44 31.96 85.44 31.96 96.32 ;
    LAYER li1 ;
      POLYGON 103.96 98.005 103.96 97.835 100.265 97.835 100.265 97.035 99.935 97.035 99.935 97.835 99.425 97.835 99.425 97.355 99.095 97.355 99.095 97.835 98.585 97.835 98.585 97.355 98.255 97.355 98.255 97.835 97.745 97.835 97.745 97.355 97.415 97.355 97.415 97.835 96.905 97.835 96.905 97.355 96.575 97.355 96.575 97.835 96.065 97.835 96.065 97.355 95.735 97.355 95.735 97.835 94.705 97.835 94.705 97.355 94.375 97.355 94.375 97.835 93.865 97.835 93.865 97.355 93.535 97.355 93.535 97.835 93.025 97.835 93.025 97.355 92.695 97.355 92.695 97.835 92.185 97.835 92.185 97.355 91.855 97.355 91.855 97.835 91.345 97.835 91.345 97.355 91.015 97.355 91.015 97.835 90.505 97.835 90.505 97.035 90.175 97.035 90.175 97.835 89.225 97.835 89.225 97.035 88.895 97.035 88.895 97.835 88.385 97.835 88.385 97.355 88.055 97.355 88.055 97.835 87.545 97.835 87.545 97.355 87.215 97.355 87.215 97.835 86.705 97.835 86.705 97.355 86.375 97.355 86.375 97.835 85.865 97.835 85.865 97.355 85.535 97.355 85.535 97.835 85.025 97.835 85.025 97.355 84.695 97.355 84.695 97.835 83.705 97.835 83.705 97.035 83.375 97.035 83.375 97.835 82.865 97.835 82.865 97.355 82.535 97.355 82.535 97.835 82.025 97.835 82.025 97.355 81.695 97.355 81.695 97.835 81.185 97.835 81.185 97.355 80.855 97.355 80.855 97.835 80.345 97.835 80.345 97.355 80.015 97.355 80.015 97.835 79.505 97.835 79.505 97.355 79.175 97.355 79.175 97.835 77.485 97.835 77.485 97.375 77.23 97.375 77.23 97.835 76.56 97.835 76.56 97.375 76.39 97.375 76.39 97.835 75.72 97.835 75.72 97.375 75.55 97.375 75.55 97.835 74.88 97.835 74.88 97.375 74.71 97.375 74.71 97.835 74.04 97.835 74.04 97.375 73.735 97.375 73.735 97.835 73.165 97.835 73.165 97.355 72.995 97.355 72.995 97.835 72.325 97.835 72.325 97.355 72.155 97.355 72.155 97.835 71.565 97.835 71.565 97.355 71.235 97.355 71.235 97.835 70.725 97.835 70.725 97.355 70.395 97.355 70.395 97.835 69.885 97.835 69.885 97.035 69.555 97.035 69.555 97.835 67.565 97.835 67.565 97.355 67.235 97.355 67.235 97.835 66.725 97.835 66.725 97.355 66.395 97.355 66.395 97.835 65.885 97.835 65.885 97.355 65.555 97.355 65.555 97.835 65.045 97.835 65.045 97.355 64.715 97.355 64.715 97.835 64.205 97.835 64.205 97.355 63.875 97.355 63.875 97.835 63.365 97.835 63.365 97.035 63.035 97.035 63.035 97.835 62.305 97.835 62.305 97.375 62.05 97.375 62.05 97.835 61.38 97.835 61.38 97.375 61.21 97.375 61.21 97.835 60.54 97.835 60.54 97.375 60.37 97.375 60.37 97.835 59.7 97.835 59.7 97.375 59.53 97.375 59.53 97.835 58.86 97.835 58.86 97.375 58.555 97.375 58.555 97.835 56.945 97.835 56.945 97.035 56.615 97.035 56.615 97.835 56.105 97.835 56.105 97.355 55.775 97.355 55.775 97.835 55.265 97.835 55.265 97.355 54.935 97.355 54.935 97.835 54.345 97.835 54.345 97.355 54.175 97.355 54.175 97.835 53.505 97.835 53.505 97.355 53.335 97.355 53.335 97.835 51.465 97.835 51.465 97.375 51.16 97.375 51.16 97.835 49.675 97.835 49.675 97.395 49.485 97.395 49.485 97.835 47.585 97.835 47.585 97.375 47.255 97.375 47.255 97.835 44.655 97.835 44.655 97.475 44.325 97.475 44.325 97.835 43.625 97.835 43.625 97.455 43.295 97.455 43.295 97.835 41.885 97.835 41.885 97.355 41.715 97.355 41.715 97.835 41.045 97.835 41.045 97.355 40.875 97.355 40.875 97.835 40.285 97.835 40.285 97.355 39.955 97.355 39.955 97.835 39.445 97.835 39.445 97.355 39.115 97.355 39.115 97.835 38.605 97.835 38.605 97.035 38.275 97.035 38.275 97.835 37.585 97.835 37.585 97.375 37.28 97.375 37.28 97.835 36.61 97.835 36.61 97.375 36.44 97.375 36.44 97.835 35.77 97.835 35.77 97.375 35.6 97.375 35.6 97.835 34.93 97.835 34.93 97.375 34.76 97.375 34.76 97.835 34.09 97.835 34.09 97.375 33.835 97.375 33.835 97.835 30.36 97.835 30.36 98.005 ;
      RECT 103.04 95.115 103.96 95.285 ;
      RECT 30.36 95.115 32.2 95.285 ;
      RECT 103.04 92.395 103.96 92.565 ;
      RECT 30.36 92.395 32.2 92.565 ;
      RECT 103.04 89.675 103.96 89.845 ;
      RECT 30.36 89.675 32.2 89.845 ;
      POLYGON 134.32 87.125 134.32 86.955 130.085 86.955 130.085 86.155 129.755 86.155 129.755 86.955 129.245 86.955 129.245 86.475 128.915 86.475 128.915 86.955 128.405 86.955 128.405 86.475 128.075 86.475 128.075 86.955 127.485 86.955 127.485 86.475 127.315 86.475 127.315 86.955 126.645 86.955 126.645 86.475 126.475 86.475 126.475 86.955 125.565 86.955 125.565 86.155 125.235 86.155 125.235 86.955 124.725 86.955 124.725 86.475 124.395 86.475 124.395 86.955 123.885 86.955 123.885 86.475 123.555 86.475 123.555 86.955 123.045 86.955 123.045 86.475 122.715 86.475 122.715 86.955 122.205 86.955 122.205 86.475 121.875 86.475 121.875 86.955 121.365 86.955 121.365 86.475 121.035 86.475 121.035 86.955 120.005 86.955 120.005 86.495 119.7 86.495 119.7 86.955 118.215 86.955 118.215 86.515 118.025 86.515 118.025 86.955 116.125 86.955 116.125 86.495 115.795 86.495 115.795 86.955 113.195 86.955 113.195 86.595 112.865 86.595 112.865 86.955 112.165 86.955 112.165 86.575 111.835 86.575 111.835 86.955 110.805 86.955 110.805 86.495 110.5 86.495 110.5 86.955 109.015 86.955 109.015 86.515 108.825 86.515 108.825 86.955 106.925 86.955 106.925 86.495 106.595 86.495 106.595 86.955 103.995 86.955 103.995 86.595 103.665 86.595 103.665 86.955 102.965 86.955 102.965 86.575 102.635 86.575 102.635 86.955 102.12 86.955 102.12 87.125 ;
      POLYGON 32.2 87.125 32.2 86.955 31.685 86.955 31.685 86.495 31.38 86.495 31.38 86.955 29.895 86.955 29.895 86.515 29.705 86.515 29.705 86.955 27.805 86.955 27.805 86.495 27.475 86.495 27.475 86.955 24.875 86.955 24.875 86.595 24.545 86.595 24.545 86.955 23.845 86.955 23.845 86.575 23.515 86.575 23.515 86.955 22.17 86.955 22.17 86.135 21.94 86.135 21.94 86.955 21.105 86.955 21.105 86.555 20.775 86.555 20.775 86.955 18.815 86.955 18.815 86.42 18.305 86.42 18.305 86.955 16.965 86.955 16.965 86.495 16.66 86.495 16.66 86.955 15.175 86.955 15.175 86.515 14.985 86.515 14.985 86.955 13.085 86.955 13.085 86.495 12.755 86.495 12.755 86.955 10.155 86.955 10.155 86.595 9.825 86.595 9.825 86.955 9.125 86.955 9.125 86.575 8.795 86.575 8.795 86.955 7.805 86.955 7.805 86.155 7.475 86.155 7.475 86.955 6.965 86.955 6.965 86.475 6.635 86.475 6.635 86.955 6.125 86.955 6.125 86.475 5.795 86.475 5.795 86.955 5.285 86.955 5.285 86.475 4.955 86.475 4.955 86.955 4.445 86.955 4.445 86.475 4.115 86.475 4.115 86.955 3.605 86.955 3.605 86.475 3.275 86.475 3.275 86.955 0 86.955 0 87.125 ;
      RECT 133.4 84.235 134.32 84.405 ;
      RECT 0 84.235 1.84 84.405 ;
      RECT 133.4 81.515 134.32 81.685 ;
      RECT 0 81.515 1.84 81.685 ;
      RECT 133.4 78.795 134.32 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 133.4 76.075 134.32 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 133.4 73.355 134.32 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 133.4 70.635 134.32 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 133.4 67.915 134.32 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 133.4 65.195 134.32 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 133.4 62.475 134.32 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 133.4 59.755 134.32 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 133.4 57.035 134.32 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 133.4 54.315 134.32 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 133.4 51.595 134.32 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 133.4 48.875 134.32 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 133.4 46.155 134.32 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 133.4 43.435 134.32 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 133.4 40.715 134.32 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 133.4 37.995 134.32 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 133.4 35.275 134.32 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 133.4 32.555 134.32 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 132.48 29.835 134.32 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 132.48 27.115 134.32 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 133.4 24.395 134.32 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 133.4 21.675 134.32 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 133.4 18.955 134.32 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 133.4 16.235 134.32 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 133.4 13.515 134.32 13.685 ;
      RECT 0 13.515 1.84 13.685 ;
      POLYGON 8.42 11.785 8.42 10.965 9.565 10.965 9.565 11.5 10.075 11.5 10.075 10.965 12.035 10.965 12.035 11.365 12.365 11.365 12.365 10.965 13.395 10.965 13.395 11.365 13.725 11.365 13.725 10.965 15.685 10.965 15.685 11.5 16.195 11.5 16.195 10.965 17.535 10.965 17.535 11.345 17.865 11.345 17.865 10.965 18.565 10.965 18.565 11.325 18.895 11.325 18.895 10.965 21.495 10.965 21.495 11.425 21.825 11.425 21.825 10.965 23.725 10.965 23.725 11.405 23.915 11.405 23.915 10.965 25.4 10.965 25.4 11.425 25.705 11.425 25.705 10.965 26.745 10.965 26.745 11.345 27.075 11.345 27.075 10.965 28.115 10.965 28.115 11.345 28.445 11.345 28.445 10.965 29.145 10.965 29.145 11.325 29.475 11.325 29.475 10.965 32.075 10.965 32.075 11.425 32.405 11.425 32.405 10.965 34.305 10.965 34.305 11.405 34.495 11.405 34.495 10.965 35.98 10.965 35.98 11.425 36.285 11.425 36.285 10.965 36.8 10.965 36.8 10.795 0 10.795 0 10.965 3.315 10.965 3.315 11.765 3.645 11.765 3.645 10.965 4.155 10.965 4.155 11.445 4.485 11.445 4.485 10.965 4.995 10.965 4.995 11.445 5.325 11.445 5.325 10.965 5.915 10.965 5.915 11.445 6.085 11.445 6.085 10.965 6.755 10.965 6.755 11.445 6.925 11.445 6.925 10.965 8.19 10.965 8.19 11.785 ;
      POLYGON 118.635 11.5 118.635 10.965 120.595 10.965 120.595 11.365 120.925 11.365 120.925 10.965 122.415 10.965 122.415 11.345 122.745 11.345 122.745 10.965 123.445 10.965 123.445 11.325 123.775 11.325 123.775 10.965 126.375 10.965 126.375 11.425 126.705 11.425 126.705 10.965 128.605 10.965 128.605 11.405 128.795 11.405 128.795 10.965 130.28 10.965 130.28 11.425 130.585 11.425 130.585 10.965 134.32 10.965 134.32 10.795 102.58 10.795 102.58 10.965 103.405 10.965 103.405 11.5 103.915 11.5 103.915 10.965 105.875 10.965 105.875 11.365 106.205 11.365 106.205 10.965 107.235 10.965 107.235 11.345 107.565 11.345 107.565 10.965 108.265 10.965 108.265 11.325 108.595 11.325 108.595 10.965 111.195 10.965 111.195 11.425 111.525 11.425 111.525 10.965 113.425 10.965 113.425 11.405 113.615 11.405 113.615 10.965 115.1 10.965 115.1 11.425 115.405 11.425 115.405 10.965 116.445 10.965 116.445 11.345 116.775 11.345 116.775 10.965 118.125 10.965 118.125 11.5 ;
      RECT 100.28 8.075 103.96 8.245 ;
      RECT 30.36 8.075 32.2 8.245 ;
      RECT 100.28 5.355 103.96 5.525 ;
      RECT 30.36 5.355 32.2 5.525 ;
      RECT 102.12 2.635 103.96 2.805 ;
      RECT 30.36 2.635 34.04 2.805 ;
      POLYGON 97.965 0.885 97.965 0.085 103.96 0.085 103.96 -0.085 30.36 -0.085 30.36 0.085 34.515 0.085 34.515 0.885 34.845 0.885 34.845 0.085 35.355 0.085 35.355 0.565 35.685 0.565 35.685 0.085 36.195 0.085 36.195 0.565 36.525 0.565 36.525 0.085 37.035 0.085 37.035 0.565 37.365 0.565 37.365 0.085 37.875 0.085 37.875 0.565 38.205 0.565 38.205 0.085 38.715 0.085 38.715 0.565 39.045 0.565 39.045 0.085 40.075 0.085 40.075 0.485 40.405 0.485 40.405 0.085 42.365 0.085 42.365 0.62 42.875 0.62 42.875 0.085 44.215 0.085 44.215 0.465 44.545 0.465 44.545 0.085 45.245 0.085 45.245 0.445 45.575 0.445 45.575 0.085 48.175 0.085 48.175 0.545 48.505 0.545 48.505 0.085 50.405 0.085 50.405 0.525 50.595 0.525 50.595 0.085 52.08 0.085 52.08 0.545 52.385 0.545 52.385 0.085 53.425 0.085 53.425 0.465 53.755 0.465 53.755 0.085 54.755 0.085 54.755 0.885 55.085 0.885 55.085 0.085 55.595 0.085 55.595 0.565 55.925 0.565 55.925 0.085 56.435 0.085 56.435 0.565 56.765 0.565 56.765 0.085 57.275 0.085 57.275 0.565 57.605 0.565 57.605 0.085 58.115 0.085 58.115 0.565 58.445 0.565 58.445 0.085 58.955 0.085 58.955 0.565 59.285 0.565 59.285 0.085 60.325 0.085 60.325 0.565 60.565 0.565 60.565 0.085 61.155 0.085 61.155 0.565 61.485 0.565 61.485 0.085 61.995 0.085 61.995 0.885 62.325 0.885 62.325 0.085 62.815 0.085 62.815 0.545 63.07 0.545 63.07 0.085 63.74 0.085 63.74 0.545 63.91 0.545 63.91 0.085 64.58 0.085 64.58 0.545 64.75 0.545 64.75 0.085 65.42 0.085 65.42 0.545 65.59 0.545 65.59 0.085 66.26 0.085 66.26 0.545 66.565 0.545 66.565 0.085 67.215 0.085 67.215 0.565 67.545 0.565 67.545 0.085 68.055 0.085 68.055 0.565 68.385 0.565 68.385 0.085 68.895 0.085 68.895 0.565 69.225 0.565 69.225 0.085 69.735 0.085 69.735 0.565 70.065 0.565 70.065 0.085 70.575 0.085 70.575 0.565 70.905 0.565 70.905 0.085 71.415 0.085 71.415 0.885 71.745 0.885 71.745 0.085 72.735 0.085 72.735 0.565 73.065 0.565 73.065 0.085 73.575 0.085 73.575 0.565 73.905 0.565 73.905 0.085 74.415 0.085 74.415 0.565 74.745 0.565 74.745 0.085 75.255 0.085 75.255 0.565 75.585 0.565 75.585 0.085 76.095 0.085 76.095 0.565 76.425 0.565 76.425 0.085 76.935 0.085 76.935 0.885 77.265 0.885 77.265 0.085 78.255 0.085 78.255 0.565 78.585 0.565 78.585 0.085 79.095 0.085 79.095 0.565 79.425 0.565 79.425 0.085 79.935 0.085 79.935 0.565 80.265 0.565 80.265 0.085 80.775 0.085 80.775 0.565 81.105 0.565 81.105 0.085 81.615 0.085 81.615 0.565 81.945 0.565 81.945 0.085 82.455 0.085 82.455 0.885 82.785 0.885 82.785 0.085 83.395 0.085 83.395 0.545 83.7 0.545 83.7 0.085 84.37 0.085 84.37 0.545 84.54 0.545 84.54 0.085 85.21 0.085 85.21 0.545 85.38 0.545 85.38 0.085 86.05 0.085 86.05 0.545 86.22 0.545 86.22 0.085 86.89 0.085 86.89 0.545 87.145 0.545 87.145 0.085 87.875 0.085 87.875 0.885 88.205 0.885 88.205 0.085 88.715 0.085 88.715 0.565 89.045 0.565 89.045 0.085 89.555 0.085 89.555 0.565 89.885 0.565 89.885 0.085 90.395 0.085 90.395 0.565 90.725 0.565 90.725 0.085 91.235 0.085 91.235 0.565 91.565 0.565 91.565 0.085 92.075 0.085 92.075 0.565 92.405 0.565 92.405 0.085 93.435 0.085 93.435 0.565 93.765 0.565 93.765 0.085 94.275 0.085 94.275 0.565 94.605 0.565 94.605 0.085 95.115 0.085 95.115 0.565 95.445 0.565 95.445 0.085 95.955 0.085 95.955 0.565 96.285 0.565 96.285 0.085 96.795 0.085 96.795 0.565 97.125 0.565 97.125 0.085 97.635 0.085 97.635 0.885 ;
      POLYGON 103.79 97.75 103.79 86.87 134.15 86.87 134.15 11.05 103.79 11.05 103.79 0.17 30.53 0.17 30.53 11.05 0.17 11.05 0.17 86.87 30.53 86.87 30.53 97.75 ;
    LAYER via ;
      RECT 89.165 97.725 89.315 97.875 ;
      RECT 59.725 97.725 59.875 97.875 ;
      RECT 80.195 97.335 80.345 97.485 ;
      RECT 61.795 97.335 61.945 97.485 ;
      RECT 123.895 11.315 124.045 11.465 ;
      RECT 75.135 0.435 75.285 0.585 ;
      RECT 68.235 0.435 68.385 0.585 ;
      RECT 57.195 0.435 57.345 0.585 ;
      RECT 89.165 0.045 89.315 0.195 ;
      RECT 59.725 0.045 59.875 0.195 ;
    LAYER via2 ;
      RECT 89.14 97.7 89.34 97.9 ;
      RECT 59.7 97.7 59.9 97.9 ;
      RECT 96.73 97.48 96.93 97.68 ;
      RECT 95.81 97.48 96.01 97.68 ;
      RECT 31.41 97.48 31.61 97.68 ;
      RECT 125.71 86.6 125.91 86.8 ;
      RECT 26.35 86.6 26.55 86.8 ;
      RECT 15.77 86.6 15.97 86.8 ;
      RECT 13.93 86.6 14.13 86.8 ;
      RECT 133.07 62.12 133.27 62.32 ;
      RECT 1.05 52.6 1.25 52.8 ;
      RECT 133.07 45.8 133.27 46 ;
      RECT 1.05 44.44 1.25 44.64 ;
      RECT 133.07 41.72 133.27 41.92 ;
      RECT 24.05 11.12 24.25 11.32 ;
      RECT 18.07 11.12 18.27 11.32 ;
      RECT 62.69 0.24 62.89 0.44 ;
      RECT 89.14 0.02 89.34 0.22 ;
      RECT 59.7 0.02 59.9 0.22 ;
    LAYER via3 ;
      RECT 89.14 97.7 89.34 97.9 ;
      RECT 59.7 97.7 59.9 97.9 ;
      RECT 86.84 97.48 87.04 97.68 ;
      RECT 70.28 97.48 70.48 97.68 ;
      RECT 65.68 97.48 65.88 97.68 ;
      RECT 61.08 97.48 61.28 97.68 ;
      RECT 50.04 97.48 50.24 97.68 ;
      RECT 92.36 0.92 92.56 1.12 ;
      RECT 78.56 0.92 78.76 1.12 ;
      RECT 64.76 0.24 64.96 0.44 ;
      RECT 63.84 0.24 64.04 0.44 ;
      RECT 89.14 0.02 89.34 0.22 ;
      RECT 59.7 0.02 59.9 0.22 ;
    LAYER OVERLAP ;
      POLYGON 30.36 0 30.36 10.88 0 10.88 0 87.04 30.36 87.04 30.36 97.92 103.96 97.92 103.96 87.04 134.32 87.04 134.32 10.88 103.96 10.88 103.96 0 ;
  END
END sb_1__1_

END LIBRARY
