VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO cbx_1__0_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 75.44 BY 119.68 ;
  SYMMETRY X Y ;
  PIN pReset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 66.06 0.595 66.2 ;
    END
  END pReset[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 44.64 0.595 44.78 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 77.96 0.595 78.1 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 63.34 0.595 63.48 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 115.02 0.595 115.16 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 115.7 0.595 115.84 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 29 0.595 29.14 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 102.19 0.8 102.49 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 101.42 0.595 101.56 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 80 0.595 80.14 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 113.32 0.595 113.46 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 117.74 0.595 117.88 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 88.16 0.595 88.3 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 94.28 0.595 94.42 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 99.72 0.595 99.86 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 72.52 0.595 72.66 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 97 0.595 97.14 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 95.98 0.595 96.12 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 91.22 0.595 91.36 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 103.55 0.8 103.85 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 104.91 0.8 105.21 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 80.68 0.595 80.82 ;
    END
  END chanx_left_in[20]
  PIN chanx_left_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 104.14 0.595 104.28 ;
    END
  END chanx_left_in[21]
  PIN chanx_left_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 106.27 0.8 106.57 ;
    END
  END chanx_left_in[22]
  PIN chanx_left_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 90.54 0.595 90.68 ;
    END
  END chanx_left_in[23]
  PIN chanx_left_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 96.07 0.8 96.37 ;
    END
  END chanx_left_in[24]
  PIN chanx_left_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 108.31 0.8 108.61 ;
    END
  END chanx_left_in[25]
  PIN chanx_left_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 85.78 0.595 85.92 ;
    END
  END chanx_left_in[26]
  PIN chanx_left_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 112.3 0.595 112.44 ;
    END
  END chanx_left_in[27]
  PIN chanx_left_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 111.71 0.8 112.01 ;
    END
  END chanx_left_in[28]
  PIN chanx_left_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 88.84 0.595 88.98 ;
    END
  END chanx_left_in[29]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 85.19 75.44 85.49 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 55.52 75.44 55.66 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 60.96 75.44 61.1 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 83.83 75.44 84.13 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 115.7 75.44 115.84 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 61.64 75.44 61.78 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 87.82 75.44 87.96 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 94.28 75.44 94.42 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 82.72 75.44 82.86 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 99.04 75.44 99.18 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 117.74 75.44 117.88 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 93.6 75.44 93.74 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 99.72 75.44 99.86 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 91.22 75.44 91.36 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 80.68 75.44 80.82 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 112.98 75.44 113.12 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 101.76 75.44 101.9 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 90.54 75.44 90.68 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 110.26 75.44 110.4 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 109.67 75.44 109.97 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 82.47 75.44 82.77 ;
    END
  END chanx_right_in[20]
  PIN chanx_right_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 97 75.44 97.14 ;
    END
  END chanx_right_in[21]
  PIN chanx_right_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 79.75 75.44 80.05 ;
    END
  END chanx_right_in[22]
  PIN chanx_right_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 83.4 75.44 83.54 ;
    END
  END chanx_right_in[23]
  PIN chanx_right_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 107.54 75.44 107.68 ;
    END
  END chanx_right_in[24]
  PIN chanx_right_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 109.58 75.44 109.72 ;
    END
  END chanx_right_in[25]
  PIN chanx_right_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 80 75.44 80.14 ;
    END
  END chanx_right_in[26]
  PIN chanx_right_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 112.3 75.44 112.44 ;
    END
  END chanx_right_in[27]
  PIN chanx_right_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 105.16 75.44 105.3 ;
    END
  END chanx_right_in[28]
  PIN chanx_right_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 106.86 75.44 107 ;
    END
  END chanx_right_in[29]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 85.78 75.44 85.92 ;
    END
  END ccff_head[0]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 23.56 0.595 23.7 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 109.67 0.8 109.97 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 28.32 0.595 28.46 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 69.12 0.595 69.26 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 110.26 0.595 110.4 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 48.04 0.595 48.18 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 42.6 0.595 42.74 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 109.58 0.595 109.72 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 60.96 0.595 61.1 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 105.16 0.595 105.3 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 102.44 0.595 102.58 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 85.1 0.595 85.24 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 26.28 0.595 26.42 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 106.86 0.595 107 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 50.76 0.595 50.9 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 83.83 0.8 84.13 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 64.02 0.595 64.16 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 47.36 0.595 47.5 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 25.6 0.595 25.74 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 71.84 0.595 71.98 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 98.7 0.595 98.84 ;
    END
  END chanx_left_out[20]
  PIN chanx_left_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 93.6 0.595 93.74 ;
    END
  END chanx_left_out[21]
  PIN chanx_left_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 85.19 0.8 85.49 ;
    END
  END chanx_left_out[22]
  PIN chanx_left_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 82.72 0.595 82.86 ;
    END
  END chanx_left_out[23]
  PIN chanx_left_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 45.32 0.595 45.46 ;
    END
  END chanx_left_out[24]
  PIN chanx_left_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 107.54 0.595 107.68 ;
    END
  END chanx_left_out[25]
  PIN chanx_left_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 97.43 0.8 97.73 ;
    END
  END chanx_left_out[26]
  PIN chanx_left_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 50.08 0.595 50.22 ;
    END
  END chanx_left_out[27]
  PIN chanx_left_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 69.8 0.595 69.94 ;
    END
  END chanx_left_out[28]
  PIN chanx_left_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 83.4 0.595 83.54 ;
    END
  END chanx_left_out[29]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 69.8 75.44 69.94 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 106.95 75.44 107.25 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 115.02 75.44 115.16 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 47.36 75.44 47.5 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 72.52 75.44 72.66 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 63.34 75.44 63.48 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 48.04 75.44 48.18 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 71.84 75.44 71.98 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 45.32 75.44 45.46 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 101.51 75.44 101.81 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 50.08 75.44 50.22 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 58.92 75.44 59.06 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 85.1 75.44 85.24 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 105.59 75.44 105.89 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 95.39 75.44 95.69 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 102.44 75.44 102.58 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 104.48 75.44 104.62 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 98.79 75.44 99.09 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 111.03 75.44 111.33 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 87.91 75.44 88.21 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 88.5 75.44 88.64 ;
    END
  END chanx_right_out[20]
  PIN chanx_right_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 102.87 75.44 103.17 ;
    END
  END chanx_right_out[21]
  PIN chanx_right_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 81.11 75.44 81.41 ;
    END
  END chanx_right_out[22]
  PIN chanx_right_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 58.24 75.44 58.38 ;
    END
  END chanx_right_out[23]
  PIN chanx_right_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 56.2 75.44 56.34 ;
    END
  END chanx_right_out[24]
  PIN chanx_right_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 108.31 75.44 108.61 ;
    END
  END chanx_right_out[25]
  PIN chanx_right_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 86.55 75.44 86.85 ;
    END
  END chanx_right_out[26]
  PIN chanx_right_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 112.39 75.44 112.69 ;
    END
  END chanx_right_out[27]
  PIN chanx_right_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 100.15 75.44 100.45 ;
    END
  END chanx_right_out[28]
  PIN chanx_right_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 104.23 75.44 104.53 ;
    END
  END chanx_right_out[29]
  PIN bottom_grid_pin_0_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 41.92 75.44 42.06 ;
    END
  END bottom_grid_pin_0_[0]
  PIN bottom_grid_pin_2_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 36.82 75.44 36.96 ;
    END
  END bottom_grid_pin_2_[0]
  PIN bottom_grid_pin_4_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 0 39.4 0.485 ;
    END
  END bottom_grid_pin_4_[0]
  PIN bottom_grid_pin_6_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 53.14 0.595 53.28 ;
    END
  END bottom_grid_pin_6_[0]
  PIN bottom_grid_pin_8_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 30.7 75.44 30.84 ;
    END
  END bottom_grid_pin_8_[0]
  PIN bottom_grid_pin_10_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.7 0 45.84 0.485 ;
    END
  END bottom_grid_pin_10_[0]
  PIN bottom_grid_pin_12_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.86 0 44 0.485 ;
    END
  END bottom_grid_pin_12_[0]
  PIN bottom_grid_pin_14_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 31.38 0.595 31.52 ;
    END
  END bottom_grid_pin_14_[0]
  PIN bottom_grid_pin_16_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 34.1 0.595 34.24 ;
    END
  END bottom_grid_pin_16_[0]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 61.64 0.595 61.78 ;
    END
  END ccff_tail[0]
  PIN IO_ISOL_N[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 90.63 0.8 90.93 ;
    END
  END IO_ISOL_N[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 0 41.24 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.9 0 55.04 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.7 0 68.84 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.62 0 69.76 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 0 62.4 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.62 0 23.76 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.8 0 15.94 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.88 0 15.02 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.84 0 3.98 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48 0 48.14 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 0 65.16 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.46 0 71.6 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.38 0 72.52 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.4 0 66.54 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.86 0 21 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.96 0 14.1 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.72 0 16.86 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.52 0 7.66 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.94 0 43.08 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 0 56.42 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 0 64.24 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.32 0 67.46 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.88 0 61.02 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.24 0 22.38 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.04 0 13.18 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.66 0 11.8 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.92 0 3.06 0.485 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
  PIN top_width_0_height_0__pin_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 42.6 75.44 42.74 ;
    END
  END top_width_0_height_0__pin_0_[0]
  PIN top_width_0_height_0__pin_2_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 36.14 75.44 36.28 ;
    END
  END top_width_0_height_0__pin_2_[0]
  PIN top_width_0_height_0__pin_4_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.18 0 40.32 0.485 ;
    END
  END top_width_0_height_0__pin_4_[0]
  PIN top_width_0_height_0__pin_6_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 41.92 0.595 42.06 ;
    END
  END top_width_0_height_0__pin_6_[0]
  PIN top_width_0_height_0__pin_8_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 31.38 75.44 31.52 ;
    END
  END top_width_0_height_0__pin_8_[0]
  PIN top_width_0_height_0__pin_10_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.62 0 46.76 0.485 ;
    END
  END top_width_0_height_0__pin_10_[0]
  PIN top_width_0_height_0__pin_12_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.02 0 42.16 0.485 ;
    END
  END top_width_0_height_0__pin_12_[0]
  PIN top_width_0_height_0__pin_14_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 30.7 0.595 30.84 ;
    END
  END top_width_0_height_0__pin_14_[0]
  PIN top_width_0_height_0__pin_16_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 33.42 0.595 33.56 ;
    END
  END top_width_0_height_0__pin_16_[0]
  PIN top_width_0_height_0__pin_1_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 98.79 0.8 99.09 ;
    END
  END top_width_0_height_0__pin_1_upper[0]
  PIN top_width_0_height_0__pin_1_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 66.06 75.44 66.2 ;
    END
  END top_width_0_height_0__pin_1_lower[0]
  PIN top_width_0_height_0__pin_3_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 58.92 0.595 59.06 ;
    END
  END top_width_0_height_0__pin_3_upper[0]
  PIN top_width_0_height_0__pin_3_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 94.03 75.44 94.33 ;
    END
  END top_width_0_height_0__pin_3_lower[0]
  PIN top_width_0_height_0__pin_5_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 93.35 0.8 93.65 ;
    END
  END top_width_0_height_0__pin_5_upper[0]
  PIN top_width_0_height_0__pin_5_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 113.75 75.44 114.05 ;
    END
  END top_width_0_height_0__pin_5_lower[0]
  PIN top_width_0_height_0__pin_7_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 39.88 0.595 40.02 ;
    END
  END top_width_0_height_0__pin_7_upper[0]
  PIN top_width_0_height_0__pin_7_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 97.43 75.44 97.73 ;
    END
  END top_width_0_height_0__pin_7_lower[0]
  PIN top_width_0_height_0__pin_9_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 115.79 0.8 116.09 ;
    END
  END top_width_0_height_0__pin_9_upper[0]
  PIN top_width_0_height_0__pin_9_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 64.02 75.44 64.16 ;
    END
  END top_width_0_height_0__pin_9_lower[0]
  PIN top_width_0_height_0__pin_11_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 114.43 0.8 114.73 ;
    END
  END top_width_0_height_0__pin_11_upper[0]
  PIN top_width_0_height_0__pin_11_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 92.67 75.44 92.97 ;
    END
  END top_width_0_height_0__pin_11_lower[0]
  PIN top_width_0_height_0__pin_13_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 113.07 0.8 113.37 ;
    END
  END top_width_0_height_0__pin_13_upper[0]
  PIN top_width_0_height_0__pin_13_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 68.78 75.44 68.92 ;
    END
  END top_width_0_height_0__pin_13_lower[0]
  PIN top_width_0_height_0__pin_15_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 94.71 0.8 95.01 ;
    END
  END top_width_0_height_0__pin_15_upper[0]
  PIN top_width_0_height_0__pin_15_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 89.27 75.44 89.57 ;
    END
  END top_width_0_height_0__pin_15_lower[0]
  PIN top_width_0_height_0__pin_17_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 100.83 0.8 101.13 ;
    END
  END top_width_0_height_0__pin_17_upper[0]
  PIN top_width_0_height_0__pin_17_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 67.08 75.44 67.22 ;
    END
  END top_width_0_height_0__pin_17_lower[0]
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.5 119.195 36.64 119.68 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 115.79 75.44 116.09 ;
    END
  END SC_OUT_BOT
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 91.99 0.8 92.29 ;
    END
  END SC_IN_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.14 119.195 29.28 119.68 ;
    END
  END SC_OUT_TOP
  PIN pReset_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 50.76 75.44 50.9 ;
    END
  END pReset_E_in
  PIN pReset_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 52.46 0.595 52.6 ;
    END
  END pReset_W_in
  PIN pReset_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 36.14 0.595 36.28 ;
    END
  END pReset_W_out
  PIN pReset_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 95.98 75.44 96.12 ;
    END
  END pReset_E_out
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 2.92 119.195 3.06 119.68 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 0 7.24 0.595 7.38 ;
    END
  END prog_clk_0_W_out
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 17.44 3.2 20.64 ;
        RECT 72.24 17.44 75.44 20.64 ;
        RECT 0 58.24 3.2 61.44 ;
        RECT 72.24 58.24 75.44 61.44 ;
        RECT 0 99.04 3.2 102.24 ;
        RECT 72.24 99.04 75.44 102.24 ;
      LAYER met4 ;
        RECT 7.98 0 8.58 0.6 ;
        RECT 37.42 0 38.02 0.6 ;
        RECT 66.86 0 67.46 0.6 ;
        RECT 7.98 119.08 8.58 119.68 ;
        RECT 37.42 119.08 38.02 119.68 ;
        RECT 66.86 119.08 67.46 119.68 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 74.96 2.48 75.44 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 74.96 7.92 75.44 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 74.96 13.36 75.44 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 74.96 18.8 75.44 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 74.96 24.24 75.44 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 74.96 29.68 75.44 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 74.96 35.12 75.44 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 74.96 40.56 75.44 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 74.96 46 75.44 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 74.96 51.44 75.44 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 74.96 56.88 75.44 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 74.96 62.32 75.44 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 74.96 67.76 75.44 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 74.96 73.2 75.44 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 74.96 78.64 75.44 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 74.96 84.08 75.44 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 74.96 89.52 75.44 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 74.96 94.96 75.44 95.44 ;
        RECT 0 100.4 0.48 100.88 ;
        RECT 74.96 100.4 75.44 100.88 ;
        RECT 0 105.84 0.48 106.32 ;
        RECT 74.96 105.84 75.44 106.32 ;
        RECT 0 111.28 0.48 111.76 ;
        RECT 74.96 111.28 75.44 111.76 ;
        RECT 0 116.72 0.48 117.2 ;
        RECT 74.96 116.72 75.44 117.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 37.84 3.2 41.04 ;
        RECT 72.24 37.84 75.44 41.04 ;
        RECT 0 78.64 3.2 81.84 ;
        RECT 72.24 78.64 75.44 81.84 ;
      LAYER met4 ;
        RECT 22.7 0 23.3 0.6 ;
        RECT 52.14 0 52.74 0.6 ;
        RECT 22.7 119.08 23.3 119.68 ;
        RECT 52.14 119.08 52.74 119.68 ;
      LAYER met1 ;
        RECT 0 -0.24 0.48 0.24 ;
        RECT 74.96 -0.24 75.44 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 74.96 5.2 75.44 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 74.96 10.64 75.44 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 74.96 16.08 75.44 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 74.96 21.52 75.44 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 74.96 26.96 75.44 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 74.96 32.4 75.44 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 74.96 37.84 75.44 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 74.96 43.28 75.44 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 74.96 48.72 75.44 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 74.96 54.16 75.44 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 74.96 59.6 75.44 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 74.96 65.04 75.44 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 74.96 70.48 75.44 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 74.96 75.92 75.44 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 74.96 81.36 75.44 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 74.96 86.8 75.44 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 74.96 92.24 75.44 92.72 ;
        RECT 0 97.68 0.48 98.16 ;
        RECT 74.96 97.68 75.44 98.16 ;
        RECT 0 103.12 0.48 103.6 ;
        RECT 74.96 103.12 75.44 103.6 ;
        RECT 0 108.56 0.48 109.04 ;
        RECT 74.96 108.56 75.44 109.04 ;
        RECT 0 114 0.48 114.48 ;
        RECT 74.96 114 75.44 114.48 ;
        RECT 0 119.44 0.48 119.92 ;
        RECT 74.96 119.44 75.44 119.92 ;
    END
  END VSS
  OBS
    LAYER met1 ;
      POLYGON 74.68 119.92 74.68 119.44 52.6 119.44 52.6 119.43 52.28 119.43 52.28 119.44 23.16 119.44 23.16 119.43 22.84 119.43 22.84 119.44 0.76 119.44 0.76 119.92 ;
      POLYGON 74.915 98.76 74.915 98.36 71 98.36 71 98.5 74.775 98.5 74.775 98.76 ;
      POLYGON 4.44 92.04 4.44 91.9 0.665 91.9 0.665 91.64 0.525 91.64 0.525 92.04 ;
      POLYGON 52.6 0.25 52.6 0.24 74.68 0.24 74.68 -0.24 0.76 -0.24 0.76 0.24 22.84 0.24 22.84 0.25 23.16 0.25 23.16 0.24 52.28 0.24 52.28 0.25 ;
      POLYGON 74.68 119.4 74.68 119.16 75.16 119.16 75.16 118.16 74.565 118.16 74.565 117.46 74.68 117.46 74.68 116.44 75.16 116.44 75.16 116.12 74.565 116.12 74.565 114.74 74.68 114.74 74.68 113.72 75.16 113.72 75.16 113.4 74.565 113.4 74.565 112.02 74.68 112.02 74.68 111 75.16 111 75.16 110.68 74.565 110.68 74.565 109.3 74.68 109.3 74.68 108.28 75.16 108.28 75.16 107.96 74.565 107.96 74.565 106.58 74.68 106.58 74.68 105.58 74.565 105.58 74.565 104.2 75.16 104.2 75.16 103.88 74.68 103.88 74.68 102.86 74.565 102.86 74.565 101.48 75.16 101.48 75.16 101.16 74.68 101.16 74.68 100.14 74.565 100.14 74.565 98.76 75.16 98.76 75.16 98.44 74.68 98.44 74.68 97.42 74.565 97.42 74.565 96.72 75.16 96.72 75.16 96.4 74.565 96.4 74.565 95.7 74.68 95.7 74.68 94.7 74.565 94.7 74.565 93.32 75.16 93.32 75.16 93 74.68 93 74.68 91.96 75.16 91.96 75.16 91.64 74.565 91.64 74.565 90.26 74.68 90.26 74.68 89.24 75.16 89.24 75.16 88.92 74.565 88.92 74.565 87.54 74.68 87.54 74.68 86.52 75.16 86.52 75.16 86.2 74.565 86.2 74.565 84.82 74.68 84.82 74.68 83.82 74.565 83.82 74.565 82.44 75.16 82.44 75.16 82.12 74.68 82.12 74.68 81.1 74.565 81.1 74.565 79.72 75.16 79.72 75.16 79.4 74.68 79.4 74.68 78.36 75.16 78.36 75.16 76.68 74.68 76.68 74.68 75.64 75.16 75.64 75.16 73.96 74.68 73.96 74.68 72.94 74.565 72.94 74.565 71.56 75.16 71.56 75.16 71.24 74.68 71.24 74.68 70.22 74.565 70.22 74.565 69.52 75.16 69.52 75.16 69.2 74.565 69.2 74.565 68.5 74.68 68.5 74.68 67.5 74.565 67.5 74.565 66.8 75.16 66.8 75.16 66.48 74.565 66.48 74.565 65.78 74.68 65.78 74.68 64.76 75.16 64.76 75.16 64.44 74.565 64.44 74.565 63.06 74.68 63.06 74.68 62.06 74.565 62.06 74.565 60.68 75.16 60.68 75.16 60.36 74.68 60.36 74.68 59.34 74.565 59.34 74.565 57.96 75.16 57.96 75.16 57.64 74.68 57.64 74.68 56.62 74.565 56.62 74.565 55.24 75.16 55.24 75.16 54.92 74.68 54.92 74.68 53.88 75.16 53.88 75.16 52.2 74.68 52.2 74.68 51.18 74.565 51.18 74.565 49.8 75.16 49.8 75.16 49.48 74.68 49.48 74.68 48.46 74.565 48.46 74.565 47.08 75.16 47.08 75.16 46.76 74.68 46.76 74.68 45.74 74.565 45.74 74.565 45.04 75.16 45.04 75.16 44.04 74.68 44.04 74.68 43.02 74.565 43.02 74.565 41.64 75.16 41.64 75.16 41.32 74.68 41.32 74.68 40.28 75.16 40.28 75.16 38.6 74.68 38.6 74.68 37.56 75.16 37.56 75.16 37.24 74.565 37.24 74.565 35.86 74.68 35.86 74.68 34.84 75.16 34.84 75.16 33.16 74.68 33.16 74.68 32.12 75.16 32.12 75.16 31.8 74.565 31.8 74.565 30.42 74.68 30.42 74.68 29.4 75.16 29.4 75.16 27.72 74.68 27.72 74.68 26.68 75.16 26.68 75.16 25 74.68 25 74.68 23.96 75.16 23.96 75.16 22.28 74.68 22.28 74.68 21.24 75.16 21.24 75.16 19.56 74.68 19.56 74.68 18.52 75.16 18.52 75.16 16.84 74.68 16.84 74.68 15.8 75.16 15.8 75.16 14.12 74.68 14.12 74.68 13.08 75.16 13.08 75.16 11.4 74.68 11.4 74.68 10.36 75.16 10.36 75.16 8.68 74.68 8.68 74.68 7.64 75.16 7.64 75.16 5.96 74.68 5.96 74.68 4.92 75.16 4.92 75.16 3.24 74.68 3.24 74.68 2.2 75.16 2.2 75.16 0.52 74.68 0.52 74.68 0.28 0.76 0.28 0.76 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 6.96 0.875 6.96 0.875 7.66 0.76 7.66 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.28 0.875 23.28 0.875 23.98 0.76 23.98 0.76 25 0.28 25 0.28 25.32 0.875 25.32 0.875 26.7 0.76 26.7 0.76 27.72 0.28 27.72 0.28 28.04 0.875 28.04 0.875 29.42 0.76 29.42 0.76 30.42 0.875 30.42 0.875 31.8 0.28 31.8 0.28 32.12 0.76 32.12 0.76 33.14 0.875 33.14 0.875 34.52 0.28 34.52 0.28 34.84 0.76 34.84 0.76 35.86 0.875 35.86 0.875 36.56 0.28 36.56 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 39.6 0.875 39.6 0.875 40.3 0.76 40.3 0.76 41.32 0.28 41.32 0.28 41.64 0.875 41.64 0.875 43.02 0.76 43.02 0.76 44.04 0.28 44.04 0.28 44.36 0.875 44.36 0.875 45.74 0.76 45.74 0.76 46.76 0.28 46.76 0.28 47.08 0.875 47.08 0.875 48.46 0.76 48.46 0.76 49.48 0.28 49.48 0.28 49.8 0.875 49.8 0.875 51.18 0.76 51.18 0.76 52.18 0.875 52.18 0.875 53.56 0.28 53.56 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 58.64 0.875 58.64 0.875 59.34 0.76 59.34 0.76 60.36 0.28 60.36 0.28 60.68 0.875 60.68 0.875 62.06 0.76 62.06 0.76 63.06 0.875 63.06 0.875 64.44 0.28 64.44 0.28 64.76 0.76 64.76 0.76 65.78 0.875 65.78 0.875 66.48 0.28 66.48 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 68.84 0.875 68.84 0.875 70.22 0.76 70.22 0.76 71.24 0.28 71.24 0.28 71.56 0.875 71.56 0.875 72.94 0.76 72.94 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 77.68 0.875 77.68 0.875 78.38 0.76 78.38 0.76 79.4 0.28 79.4 0.28 79.72 0.875 79.72 0.875 81.1 0.76 81.1 0.76 82.12 0.28 82.12 0.28 82.44 0.875 82.44 0.875 83.82 0.76 83.82 0.76 84.82 0.875 84.82 0.875 86.2 0.28 86.2 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 87.88 0.875 87.88 0.875 89.26 0.76 89.26 0.76 90.26 0.875 90.26 0.875 91.64 0.28 91.64 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 93.32 0.875 93.32 0.875 94.7 0.76 94.7 0.76 95.7 0.875 95.7 0.875 96.4 0.28 96.4 0.28 96.72 0.875 96.72 0.875 97.42 0.76 97.42 0.76 98.42 0.875 98.42 0.875 99.12 0.28 99.12 0.28 99.44 0.875 99.44 0.875 100.14 0.76 100.14 0.76 101.14 0.875 101.14 0.875 101.84 0.28 101.84 0.28 102.16 0.875 102.16 0.875 102.86 0.76 102.86 0.76 103.86 0.875 103.86 0.875 104.56 0.28 104.56 0.28 104.88 0.875 104.88 0.875 105.58 0.76 105.58 0.76 106.58 0.875 106.58 0.875 107.96 0.28 107.96 0.28 108.28 0.76 108.28 0.76 109.3 0.875 109.3 0.875 110.68 0.28 110.68 0.28 111 0.76 111 0.76 112.02 0.875 112.02 0.875 112.72 0.28 112.72 0.28 113.04 0.875 113.04 0.875 113.74 0.76 113.74 0.76 114.74 0.875 114.74 0.875 116.12 0.28 116.12 0.28 116.44 0.76 116.44 0.76 117.46 0.875 117.46 0.875 118.16 0.28 118.16 0.28 119.16 0.76 119.16 0.76 119.4 ;
    LAYER met3 ;
      POLYGON 52.605 119.725 52.605 119.72 52.82 119.72 52.82 119.4 52.605 119.4 52.605 119.395 52.275 119.395 52.275 119.4 52.06 119.4 52.06 119.72 52.275 119.72 52.275 119.725 ;
      POLYGON 23.165 119.725 23.165 119.72 23.38 119.72 23.38 119.4 23.165 119.4 23.165 119.395 22.835 119.395 22.835 119.4 22.62 119.4 22.62 119.72 22.835 119.72 22.835 119.725 ;
      POLYGON 52.605 0.285 52.605 0.28 52.82 0.28 52.82 -0.04 52.605 -0.04 52.605 -0.045 52.275 -0.045 52.275 -0.04 52.06 -0.04 52.06 0.28 52.275 0.28 52.275 0.285 ;
      POLYGON 23.165 0.285 23.165 0.28 23.38 0.28 23.38 -0.04 23.165 -0.04 23.165 -0.045 22.835 -0.045 22.835 -0.04 22.62 -0.04 22.62 0.28 22.835 0.28 22.835 0.285 ;
      POLYGON 75.04 119.28 75.04 116.49 74.24 116.49 74.24 115.39 75.04 115.39 75.04 114.45 74.24 114.45 74.24 113.35 75.04 113.35 75.04 113.09 74.24 113.09 74.24 111.99 75.04 111.99 75.04 111.73 74.24 111.73 74.24 110.63 75.04 110.63 75.04 110.37 74.24 110.37 74.24 109.27 75.04 109.27 75.04 109.01 74.24 109.01 74.24 107.91 75.04 107.91 75.04 107.65 74.24 107.65 74.24 106.55 75.04 106.55 75.04 106.29 74.24 106.29 74.24 105.19 75.04 105.19 75.04 104.93 74.24 104.93 74.24 103.83 75.04 103.83 75.04 103.57 74.24 103.57 74.24 102.47 75.04 102.47 75.04 102.21 74.24 102.21 74.24 101.11 75.04 101.11 75.04 100.85 74.24 100.85 74.24 99.75 75.04 99.75 75.04 99.49 74.24 99.49 74.24 98.39 75.04 98.39 75.04 98.13 74.24 98.13 74.24 97.03 75.04 97.03 75.04 96.09 74.24 96.09 74.24 94.99 75.04 94.99 75.04 94.73 74.24 94.73 74.24 93.63 75.04 93.63 75.04 93.37 74.24 93.37 74.24 92.27 75.04 92.27 75.04 89.97 74.24 89.97 74.24 88.87 75.04 88.87 75.04 88.61 74.24 88.61 74.24 87.51 75.04 87.51 75.04 87.25 74.24 87.25 74.24 86.15 75.04 86.15 75.04 85.89 74.24 85.89 74.24 84.79 75.04 84.79 75.04 84.53 74.24 84.53 74.24 83.43 75.04 83.43 75.04 83.17 74.24 83.17 74.24 82.07 75.04 82.07 75.04 81.81 74.24 81.81 74.24 80.71 75.04 80.71 75.04 80.45 74.24 80.45 74.24 79.35 75.04 79.35 75.04 0.4 0.4 0.4 0.4 83.43 1.2 83.43 1.2 84.53 0.4 84.53 0.4 84.79 1.2 84.79 1.2 85.89 0.4 85.89 0.4 90.23 1.2 90.23 1.2 91.33 0.4 91.33 0.4 91.59 1.2 91.59 1.2 92.69 0.4 92.69 0.4 92.95 1.2 92.95 1.2 94.05 0.4 94.05 0.4 94.31 1.2 94.31 1.2 95.41 0.4 95.41 0.4 95.67 1.2 95.67 1.2 96.77 0.4 96.77 0.4 97.03 1.2 97.03 1.2 98.13 0.4 98.13 0.4 98.39 1.2 98.39 1.2 99.49 0.4 99.49 0.4 100.43 1.2 100.43 1.2 101.53 0.4 101.53 0.4 101.79 1.2 101.79 1.2 102.89 0.4 102.89 0.4 103.15 1.2 103.15 1.2 104.25 0.4 104.25 0.4 104.51 1.2 104.51 1.2 105.61 0.4 105.61 0.4 105.87 1.2 105.87 1.2 106.97 0.4 106.97 0.4 107.91 1.2 107.91 1.2 109.01 0.4 109.01 0.4 109.27 1.2 109.27 1.2 110.37 0.4 110.37 0.4 111.31 1.2 111.31 1.2 112.41 0.4 112.41 0.4 112.67 1.2 112.67 1.2 113.77 0.4 113.77 0.4 114.03 1.2 114.03 1.2 115.13 0.4 115.13 0.4 115.39 1.2 115.39 1.2 116.49 0.4 116.49 0.4 119.28 ;
    LAYER met2 ;
      RECT 52.3 119.375 52.58 119.745 ;
      RECT 22.86 119.375 23.14 119.745 ;
      POLYGON 67.92 9.08 67.92 0.1 67.74 0.1 67.74 0.24 67.78 0.24 67.78 9.08 ;
      RECT 20.34 0.69 20.6 1.01 ;
      RECT 52.3 -0.065 52.58 0.305 ;
      RECT 22.86 -0.065 23.14 0.305 ;
      POLYGON 75.16 119.4 75.16 0.28 72.8 0.28 72.8 0.765 72.1 0.765 72.1 0.28 71.88 0.28 71.88 0.765 71.18 0.765 71.18 0.28 70.04 0.28 70.04 0.765 69.34 0.765 69.34 0.28 69.12 0.28 69.12 0.765 68.42 0.765 68.42 0.28 67.74 0.28 67.74 0.765 67.04 0.765 67.04 0.28 66.82 0.28 66.82 0.765 66.12 0.765 66.12 0.28 65.44 0.28 65.44 0.765 64.74 0.765 64.74 0.28 64.52 0.28 64.52 0.765 63.82 0.765 63.82 0.28 62.68 0.28 62.68 0.765 61.98 0.765 61.98 0.28 61.3 0.28 61.3 0.765 60.6 0.765 60.6 0.28 56.7 0.28 56.7 0.765 56 0.765 56 0.28 55.32 0.28 55.32 0.765 54.62 0.765 54.62 0.28 48.42 0.28 48.42 0.765 47.72 0.765 47.72 0.28 47.04 0.28 47.04 0.765 46.34 0.765 46.34 0.28 46.12 0.28 46.12 0.765 45.42 0.765 45.42 0.28 44.28 0.28 44.28 0.765 43.58 0.765 43.58 0.28 43.36 0.28 43.36 0.765 42.66 0.765 42.66 0.28 42.44 0.28 42.44 0.765 41.74 0.765 41.74 0.28 41.52 0.28 41.52 0.765 40.82 0.765 40.82 0.28 40.6 0.28 40.6 0.765 39.9 0.765 39.9 0.28 39.68 0.28 39.68 0.765 38.98 0.765 38.98 0.28 24.04 0.28 24.04 0.765 23.34 0.765 23.34 0.28 22.66 0.28 22.66 0.765 21.96 0.765 21.96 0.28 21.28 0.28 21.28 0.765 20.58 0.765 20.58 0.28 17.14 0.28 17.14 0.765 16.44 0.765 16.44 0.28 16.22 0.28 16.22 0.765 15.52 0.765 15.52 0.28 15.3 0.28 15.3 0.765 14.6 0.765 14.6 0.28 14.38 0.28 14.38 0.765 13.68 0.765 13.68 0.28 13.46 0.28 13.46 0.765 12.76 0.765 12.76 0.28 12.08 0.28 12.08 0.765 11.38 0.765 11.38 0.28 7.94 0.28 7.94 0.765 7.24 0.765 7.24 0.28 4.26 0.28 4.26 0.765 3.56 0.765 3.56 0.28 3.34 0.28 3.34 0.765 2.64 0.765 2.64 0.28 0.28 0.28 0.28 119.4 2.64 119.4 2.64 118.915 3.34 118.915 3.34 119.4 28.86 119.4 28.86 118.915 29.56 118.915 29.56 119.4 36.22 119.4 36.22 118.915 36.92 118.915 36.92 119.4 ;
    LAYER met4 ;
      POLYGON 75.04 119.28 75.04 0.4 67.86 0.4 67.86 1 66.46 1 66.46 0.4 53.14 0.4 53.14 1 51.74 1 51.74 0.4 38.42 0.4 38.42 1 37.02 1 37.02 0.4 23.7 0.4 23.7 1 22.3 1 22.3 0.4 8.98 0.4 8.98 1 7.58 1 7.58 0.4 0.4 0.4 0.4 119.28 7.58 119.28 7.58 118.68 8.98 118.68 8.98 119.28 22.3 119.28 22.3 118.68 23.7 118.68 23.7 119.28 37.02 119.28 37.02 118.68 38.42 118.68 38.42 119.28 51.74 119.28 51.74 118.68 53.14 118.68 53.14 119.28 66.46 119.28 66.46 118.68 67.86 118.68 67.86 119.28 ;
    LAYER met5 ;
      POLYGON 73.84 118.08 73.84 103.84 70.64 103.84 70.64 97.44 73.84 97.44 73.84 83.44 70.64 83.44 70.64 77.04 73.84 77.04 73.84 63.04 70.64 63.04 70.64 56.64 73.84 56.64 73.84 42.64 70.64 42.64 70.64 36.24 73.84 36.24 73.84 22.24 70.64 22.24 70.64 15.84 73.84 15.84 73.84 1.6 1.6 1.6 1.6 15.84 4.8 15.84 4.8 22.24 1.6 22.24 1.6 36.24 4.8 36.24 4.8 42.64 1.6 42.64 1.6 56.64 4.8 56.64 4.8 63.04 1.6 63.04 1.6 77.04 4.8 77.04 4.8 83.44 1.6 83.44 1.6 97.44 4.8 97.44 4.8 103.84 1.6 103.84 1.6 118.08 ;
    LAYER li1 ;
      POLYGON 75.44 119.765 75.44 119.595 71.705 119.595 71.705 119.115 71.375 119.115 71.375 119.595 70.865 119.595 70.865 119.115 70.535 119.115 70.535 119.595 70.025 119.595 70.025 119.115 69.695 119.115 69.695 119.595 69.185 119.595 69.185 119.115 68.855 119.115 68.855 119.595 68.345 119.595 68.345 119.115 68.015 119.115 68.015 119.595 67.505 119.595 67.505 118.795 67.175 118.795 67.175 119.595 63.885 119.595 63.885 119.115 63.555 119.115 63.555 119.595 63.045 119.595 63.045 119.115 62.715 119.115 62.715 119.595 62.205 119.595 62.205 119.115 61.875 119.115 61.875 119.595 61.365 119.595 61.365 119.115 61.035 119.115 61.035 119.595 60.525 119.595 60.525 119.115 60.195 119.115 60.195 119.595 59.685 119.595 59.685 118.795 59.355 118.795 59.355 119.595 55.445 119.595 55.445 118.86 55.105 118.86 55.105 119.595 50.685 119.595 50.685 118.86 50.355 118.86 50.355 119.595 42.685 119.595 42.685 118.795 42.355 118.795 42.355 119.595 41.845 119.595 41.845 119.115 41.515 119.115 41.515 119.595 41.005 119.595 41.005 119.115 40.675 119.115 40.675 119.595 40.085 119.595 40.085 119.115 39.915 119.115 39.915 119.595 39.245 119.595 39.245 119.115 39.075 119.115 39.075 119.595 31.195 119.595 31.195 119.09 30.91 119.09 30.91 119.595 27.125 119.595 27.125 118.795 26.795 118.795 26.795 119.595 26.285 119.595 26.285 119.115 25.955 119.115 25.955 119.595 25.445 119.595 25.445 119.115 25.115 119.115 25.115 119.595 24.605 119.595 24.605 119.115 24.275 119.115 24.275 119.595 23.765 119.595 23.765 119.115 23.435 119.115 23.435 119.595 22.925 119.595 22.925 119.115 22.595 119.115 22.595 119.595 15.205 119.595 15.205 119.115 15.035 119.115 15.035 119.595 14.365 119.595 14.365 119.115 14.195 119.115 14.195 119.595 13.605 119.595 13.605 119.115 13.275 119.115 13.275 119.595 12.765 119.595 12.765 119.115 12.435 119.115 12.435 119.595 11.925 119.595 11.925 118.795 11.595 118.795 11.595 119.595 8.725 119.595 8.725 118.795 8.395 118.795 8.395 119.595 7.885 119.595 7.885 119.115 7.555 119.115 7.555 119.595 7.045 119.595 7.045 119.115 6.715 119.115 6.715 119.595 6.205 119.595 6.205 119.115 5.875 119.115 5.875 119.595 5.365 119.595 5.365 119.115 5.035 119.115 5.035 119.595 4.525 119.595 4.525 119.115 4.195 119.115 4.195 119.595 0 119.595 0 119.765 ;
      RECT 74.52 116.875 75.44 117.045 ;
      RECT 0 116.875 3.68 117.045 ;
      RECT 74.52 114.155 75.44 114.325 ;
      RECT 0 114.155 3.68 114.325 ;
      RECT 74.52 111.435 75.44 111.605 ;
      RECT 0 111.435 1.84 111.605 ;
      RECT 74.52 108.715 75.44 108.885 ;
      RECT 0 108.715 3.68 108.885 ;
      RECT 74.98 105.995 75.44 106.165 ;
      RECT 0 105.995 3.68 106.165 ;
      RECT 71.76 103.275 75.44 103.445 ;
      RECT 0 103.275 1.84 103.445 ;
      RECT 71.76 100.555 75.44 100.725 ;
      RECT 0 100.555 3.68 100.725 ;
      RECT 74.98 97.835 75.44 98.005 ;
      RECT 0 97.835 3.68 98.005 ;
      RECT 74.98 95.115 75.44 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 74.98 92.395 75.44 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 74.52 89.675 75.44 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 73.6 86.955 75.44 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 73.6 84.235 75.44 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 74.52 81.515 75.44 81.685 ;
      RECT 0 81.515 1.84 81.685 ;
      RECT 74.52 78.795 75.44 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 74.52 76.075 75.44 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 74.52 73.355 75.44 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 71.76 70.635 75.44 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 71.76 67.915 75.44 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 74.98 65.195 75.44 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 74.98 62.475 75.44 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 74.98 59.755 75.44 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 74.98 57.035 75.44 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 74.98 54.315 75.44 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 74.98 51.595 75.44 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 74.98 48.875 75.44 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 74.98 46.155 75.44 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 74.52 43.435 75.44 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 74.52 40.715 75.44 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 74.52 37.995 75.44 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 71.76 35.275 75.44 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 71.76 32.555 75.44 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 74.52 29.835 75.44 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 74.98 27.115 75.44 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 74.98 24.395 75.44 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 71.76 21.675 75.44 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 71.76 18.955 75.44 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 74.52 16.235 75.44 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 71.76 13.515 75.44 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 71.76 10.795 75.44 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 74.52 8.075 75.44 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 74.52 5.355 75.44 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 71.76 2.635 75.44 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      POLYGON 63.57 0.905 63.57 0.085 66.295 0.085 66.295 0.595 66.71 0.595 66.71 0.085 68.125 0.085 68.125 0.485 68.455 0.485 68.455 0.085 68.965 0.085 68.965 0.485 69.295 0.485 69.295 0.085 75.44 0.085 75.44 -0.085 0 -0.085 0 0.085 8.075 0.085 8.075 0.545 8.33 0.545 8.33 0.085 9 0.085 9 0.545 9.17 0.545 9.17 0.085 9.84 0.085 9.84 0.545 10.01 0.545 10.01 0.085 10.68 0.085 10.68 0.545 10.85 0.545 10.85 0.085 11.52 0.085 11.52 0.545 11.825 0.545 11.825 0.085 12.215 0.085 12.215 0.545 12.47 0.545 12.47 0.085 13.14 0.085 13.14 0.545 13.31 0.545 13.31 0.085 13.98 0.085 13.98 0.545 14.15 0.545 14.15 0.085 14.82 0.085 14.82 0.545 14.99 0.545 14.99 0.085 15.66 0.085 15.66 0.545 15.965 0.545 15.965 0.085 19.025 0.085 19.025 0.485 19.355 0.485 19.355 0.085 19.865 0.085 19.865 0.485 20.195 0.485 20.195 0.085 21.61 0.085 21.61 0.595 22.025 0.595 22.025 0.085 25.005 0.085 25.005 0.485 25.335 0.485 25.335 0.085 25.845 0.085 25.845 0.485 26.175 0.485 26.175 0.085 27.59 0.085 27.59 0.595 28.005 0.595 28.005 0.085 41.99 0.085 41.99 0.545 42.255 0.545 42.255 0.085 42.925 0.085 42.925 0.545 43.095 0.545 43.095 0.085 43.765 0.085 43.765 0.55 44.015 0.55 44.015 0.085 44.795 0.085 44.795 0.565 44.965 0.565 44.965 0.085 45.635 0.085 45.635 0.565 45.805 0.565 45.805 0.085 46.475 0.085 46.475 0.565 46.645 0.565 46.645 0.085 47.315 0.085 47.315 0.565 47.485 0.565 47.485 0.085 48.155 0.085 48.155 0.565 48.325 0.565 48.325 0.085 48.995 0.085 48.995 0.565 49.165 0.565 49.165 0.085 49.835 0.085 49.835 0.565 50.005 0.565 50.005 0.085 50.675 0.085 50.675 0.565 50.845 0.565 50.845 0.085 51.515 0.085 51.515 0.565 51.685 0.565 51.685 0.085 52.355 0.085 52.355 0.565 52.525 0.565 52.525 0.085 53.195 0.085 53.195 0.565 53.365 0.565 53.365 0.085 54.035 0.085 54.035 0.565 54.205 0.565 54.205 0.085 54.875 0.085 54.875 0.565 55.045 0.565 55.045 0.085 56.235 0.085 56.235 0.905 56.405 0.905 56.405 0.085 59.045 0.085 59.045 0.485 59.375 0.485 59.375 0.085 59.885 0.085 59.885 0.485 60.215 0.485 60.215 0.085 61.63 0.085 61.63 0.595 62.045 0.595 62.045 0.085 63.34 0.085 63.34 0.905 ;
      RECT 0.17 0.17 75.27 119.51 ;
    LAYER mcon ;
      RECT 55.345 119.595 55.515 119.765 ;
      RECT 54.885 119.595 55.055 119.765 ;
      RECT 54.425 119.595 54.595 119.765 ;
      RECT 53.965 119.595 54.135 119.765 ;
      RECT 53.505 119.595 53.675 119.765 ;
      RECT 53.045 119.595 53.215 119.765 ;
      RECT 52.585 119.595 52.755 119.765 ;
      RECT 52.125 119.595 52.295 119.765 ;
      RECT 51.665 119.595 51.835 119.765 ;
      RECT 51.205 119.595 51.375 119.765 ;
      RECT 50.745 119.595 50.915 119.765 ;
      RECT 50.285 119.595 50.455 119.765 ;
    LAYER via ;
      RECT 52.365 119.485 52.515 119.635 ;
      RECT 22.925 119.485 23.075 119.635 ;
      RECT 42.015 0.435 42.165 0.585 ;
      RECT 11.655 0.435 11.805 0.585 ;
      RECT 52.365 0.045 52.515 0.195 ;
      RECT 22.925 0.045 23.075 0.195 ;
    LAYER via2 ;
      RECT 52.34 119.46 52.54 119.66 ;
      RECT 22.9 119.46 23.1 119.66 ;
      RECT 1.05 106.32 1.25 106.52 ;
      RECT 52.34 0.02 52.54 0.22 ;
      RECT 22.9 0.02 23.1 0.22 ;
    LAYER via3 ;
      RECT 52.34 119.46 52.54 119.66 ;
      RECT 22.9 119.46 23.1 119.66 ;
      RECT 52.34 0.02 52.54 0.22 ;
      RECT 22.9 0.02 23.1 0.22 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 119.68 75.44 119.68 75.44 0 ;
  END
END cbx_1__0_

END LIBRARY
