VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER fieldpoly
  TYPE MASTERSLICE ;
END fieldpoly

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER diff
  TYPE MASTERSLICE ;
END diff

LAYER licon1
  TYPE MASTERSLICE ;
END licon1

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO cbx_1__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 104.88 BY 76.16 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 3.15 0 3.29 1.36 ;
    END
  END prog_clk[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.97 1.38 57.27 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 55.61 1.38 55.91 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 35.21 1.38 35.51 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 46.77 1.38 47.07 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.89 1.38 53.19 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.73 1.38 45.03 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.13 1.38 31.43 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 8.01 1.38 8.31 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 18.89 1.38 19.19 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.57 1.38 36.87 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.85 1.38 34.15 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 51.53 1.38 51.83 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 14.81 1.38 15.11 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 58.33 1.38 58.63 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 20.25 1.38 20.55 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 40.65 1.38 40.95 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 13.45 1.38 13.75 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.29 1.38 39.59 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.01 1.38 25.31 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 62.41 1.38 62.71 ;
    END
  END chanx_left_in[19]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 33.85 104.88 34.15 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 54.25 104.88 54.55 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 55.61 104.88 55.91 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 47.45 104.88 47.75 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 52.89 104.88 53.19 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 20.25 104.88 20.55 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 22.97 104.88 23.27 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 38.61 104.88 38.91 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 21.61 104.88 21.91 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 42.01 104.88 42.31 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 25.69 104.88 25.99 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 69.21 104.88 69.51 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 17.53 104.88 17.83 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 71.93 104.88 72.23 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 27.05 104.88 27.35 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.51 0 102.65 1.36 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 4.61 104.88 4.91 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 61.05 104.88 61.35 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 43.37 104.88 43.67 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 63.77 104.88 64.07 ;
    END
  END chanx_right_in[19]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 37.25 104.88 37.55 ;
    END
  END ccff_head[0]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 4.45 0 4.75 1.36 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 71.93 1.38 72.23 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 28.41 1.38 28.71 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.53 0 4.67 1.36 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 66.49 1.38 66.79 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 67.85 1.38 68.15 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.17 1.38 50.47 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.01 1.38 42.31 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 17.53 1.38 17.83 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 23.65 1.38 23.95 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 9.37 1.38 9.67 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.45 0 5.59 1.36 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.21 1.38 69.51 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.37 0 6.51 1.36 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 63.77 1.38 64.07 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.77 1.38 30.07 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 12.09 1.38 12.39 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 6.65 1.38 6.95 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.15 74.8 3.29 76.16 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 3.93 1.38 4.23 ;
    END
  END chanx_left_out[19]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 48.81 104.88 49.11 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 10.73 104.88 11.03 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.67 0 100.81 1.36 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 12.09 104.88 12.39 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 58.33 104.88 58.63 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 59.69 104.88 59.99 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 6.65 104.88 6.95 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 14.81 104.88 15.11 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 16.17 104.88 16.47 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 44.73 104.88 45.03 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 31.81 104.88 32.11 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 9.37 104.88 9.67 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 70.57 104.88 70.87 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 66.49 104.88 66.79 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 65.13 104.88 65.43 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 50.17 104.88 50.47 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.59 0 101.73 1.36 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.5 28.41 104.88 28.71 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.51 74.8 102.65 76.16 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 100.13 0 100.43 1.36 ;
    END
  END chanx_right_out[19]
  PIN top_grid_pin_16_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.97 74.8 34.11 76.16 ;
    END
  END top_grid_pin_16_[0]
  PIN top_grid_pin_17_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.81 74.8 35.95 76.16 ;
    END
  END top_grid_pin_17_[0]
  PIN top_grid_pin_18_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.89 74.8 35.03 76.16 ;
    END
  END top_grid_pin_18_[0]
  PIN top_grid_pin_19_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.73 74.8 36.87 76.16 ;
    END
  END top_grid_pin_19_[0]
  PIN top_grid_pin_20_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 74.8 57.57 76.16 ;
    END
  END top_grid_pin_20_[0]
  PIN top_grid_pin_21_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.03 74.8 16.17 76.16 ;
    END
  END top_grid_pin_21_[0]
  PIN top_grid_pin_22_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.05 74.8 33.19 76.16 ;
    END
  END top_grid_pin_22_[0]
  PIN top_grid_pin_23_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.11 74.8 15.25 76.16 ;
    END
  END top_grid_pin_23_[0]
  PIN top_grid_pin_24_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.23 74.8 2.37 76.16 ;
    END
  END top_grid_pin_24_[0]
  PIN top_grid_pin_25_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.35 74.8 12.49 76.16 ;
    END
  END top_grid_pin_25_[0]
  PIN top_grid_pin_26_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.27 74.8 13.41 76.16 ;
    END
  END top_grid_pin_26_[0]
  PIN top_grid_pin_27_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.19 74.8 14.33 76.16 ;
    END
  END top_grid_pin_27_[0]
  PIN top_grid_pin_28_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.53 74.8 73.67 76.16 ;
    END
  END top_grid_pin_28_[0]
  PIN top_grid_pin_29_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.45 74.8 74.59 76.16 ;
    END
  END top_grid_pin_29_[0]
  PIN top_grid_pin_30_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.29 74.8 76.43 76.16 ;
    END
  END top_grid_pin_30_[0]
  PIN top_grid_pin_31_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.37 74.8 75.51 76.16 ;
    END
  END top_grid_pin_31_[0]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 61.05 1.38 61.35 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.34 0 15.94 0.6 ;
        RECT 44.78 0 45.38 0.6 ;
        RECT 74.22 0 74.82 0.6 ;
        RECT 103.66 0 104.26 0.6 ;
        RECT 15.34 75.56 15.94 76.16 ;
        RECT 44.78 75.56 45.38 76.16 ;
        RECT 74.22 75.56 74.82 76.16 ;
        RECT 103.66 75.56 104.26 76.16 ;
      LAYER met5 ;
        RECT 0 16.08 3.2 19.28 ;
        RECT 101.68 16.08 104.88 19.28 ;
        RECT 0 56.88 3.2 60.08 ;
        RECT 101.68 56.88 104.88 60.08 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 104.4 2.48 104.88 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 104.4 7.92 104.88 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 104.4 13.36 104.88 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 104.4 18.8 104.88 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 104.4 24.24 104.88 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 104.4 29.68 104.88 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 104.4 35.12 104.88 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 104.4 40.56 104.88 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 104.4 46 104.88 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 104.4 51.44 104.88 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 104.4 56.88 104.88 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 104.4 62.32 104.88 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 104.4 67.76 104.88 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 104.4 73.2 104.88 73.68 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.62 0 1.22 0.6 ;
        RECT 30.06 0 30.66 0.6 ;
        RECT 59.5 0 60.1 0.6 ;
        RECT 88.94 0 89.54 0.6 ;
        RECT 0.62 75.56 1.22 76.16 ;
        RECT 30.06 75.56 30.66 76.16 ;
        RECT 59.5 75.56 60.1 76.16 ;
        RECT 88.94 75.56 89.54 76.16 ;
      LAYER met5 ;
        RECT 0 36.48 3.2 39.68 ;
        RECT 101.68 36.48 104.88 39.68 ;
      LAYER met1 ;
        RECT 0 0 104.88 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 104.4 5.2 104.88 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 104.4 10.64 104.88 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 104.4 16.08 104.88 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 104.4 21.52 104.88 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 104.4 26.96 104.88 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 104.4 32.4 104.88 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 104.4 37.84 104.88 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 104.4 43.28 104.88 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 104.4 48.72 104.88 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 104.4 54.16 104.88 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 104.4 59.6 104.88 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 104.4 65.04 104.88 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 104.4 70.48 104.88 70.96 ;
        RECT 0 75.92 104.88 76.16 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 0 76.075 104.88 76.245 ;
      RECT 103.04 73.355 104.88 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 103.96 70.635 104.88 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 103.96 67.915 104.88 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 103.96 65.195 104.88 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 103.96 62.475 104.88 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 103.96 59.755 104.88 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 103.96 57.035 104.88 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 103.96 54.315 104.88 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 103.96 51.595 104.88 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 103.96 48.875 104.88 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 103.96 46.155 104.88 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 103.96 43.435 104.88 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 103.96 40.715 104.88 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 103.96 37.995 104.88 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 103.96 35.275 104.88 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 104.42 32.555 104.88 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 103.96 29.835 104.88 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 103.96 27.115 104.88 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 103.04 24.395 104.88 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 103.04 21.675 104.88 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 103.96 18.955 104.88 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 103.96 16.235 104.88 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 103.96 13.515 104.88 13.685 ;
      RECT 0 13.515 1.84 13.685 ;
      RECT 103.96 10.795 104.88 10.965 ;
      RECT 0 10.795 1.84 10.965 ;
      RECT 103.96 8.075 104.88 8.245 ;
      RECT 0 8.075 1.84 8.245 ;
      RECT 103.96 5.355 104.88 5.525 ;
      RECT 0 5.355 1.84 5.525 ;
      RECT 103.04 2.635 104.88 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 104.88 0.085 ;
    LAYER met2 ;
      RECT 89.1 75.975 89.38 76.345 ;
      RECT 59.66 75.975 59.94 76.345 ;
      RECT 30.22 75.975 30.5 76.345 ;
      RECT 0.78 75.975 1.06 76.345 ;
      RECT 89.1 -0.185 89.38 0.185 ;
      RECT 59.66 -0.185 59.94 0.185 ;
      RECT 30.22 -0.185 30.5 0.185 ;
      RECT 0.78 -0.185 1.06 0.185 ;
      POLYGON 104.6 75.88 104.6 0.28 102.93 0.28 102.93 1.64 102.23 1.64 102.23 0.28 102.01 0.28 102.01 1.64 101.31 1.64 101.31 0.28 101.09 0.28 101.09 1.64 100.39 1.64 100.39 0.28 6.79 0.28 6.79 1.64 6.09 1.64 6.09 0.28 5.87 0.28 5.87 1.64 5.17 1.64 5.17 0.28 4.95 0.28 4.95 1.64 4.25 1.64 4.25 0.28 3.57 0.28 3.57 1.64 2.87 1.64 2.87 0.28 0.28 0.28 0.28 75.88 1.95 75.88 1.95 74.52 2.65 74.52 2.65 75.88 2.87 75.88 2.87 74.52 3.57 74.52 3.57 75.88 12.07 75.88 12.07 74.52 12.77 74.52 12.77 75.88 12.99 75.88 12.99 74.52 13.69 74.52 13.69 75.88 13.91 75.88 13.91 74.52 14.61 74.52 14.61 75.88 14.83 75.88 14.83 74.52 15.53 74.52 15.53 75.88 15.75 75.88 15.75 74.52 16.45 74.52 16.45 75.88 32.77 75.88 32.77 74.52 33.47 74.52 33.47 75.88 33.69 75.88 33.69 74.52 34.39 74.52 34.39 75.88 34.61 75.88 34.61 74.52 35.31 74.52 35.31 75.88 35.53 75.88 35.53 74.52 36.23 74.52 36.23 75.88 36.45 75.88 36.45 74.52 37.15 74.52 37.15 75.88 57.15 75.88 57.15 74.52 57.85 74.52 57.85 75.88 73.25 75.88 73.25 74.52 73.95 74.52 73.95 75.88 74.17 75.88 74.17 74.52 74.87 74.52 74.87 75.88 75.09 75.88 75.09 74.52 75.79 74.52 75.79 75.88 76.01 75.88 76.01 74.52 76.71 74.52 76.71 75.88 102.23 75.88 102.23 74.52 102.93 74.52 102.93 75.88 ;
    LAYER met3 ;
      POLYGON 89.405 76.325 89.405 76.32 89.62 76.32 89.62 76 89.405 76 89.405 75.995 89.075 75.995 89.075 76 88.86 76 88.86 76.32 89.075 76.32 89.075 76.325 ;
      POLYGON 59.965 76.325 59.965 76.32 60.18 76.32 60.18 76 59.965 76 59.965 75.995 59.635 75.995 59.635 76 59.42 76 59.42 76.32 59.635 76.32 59.635 76.325 ;
      POLYGON 30.525 76.325 30.525 76.32 30.74 76.32 30.74 76 30.525 76 30.525 75.995 30.195 75.995 30.195 76 29.98 76 29.98 76.32 30.195 76.32 30.195 76.325 ;
      POLYGON 1.085 76.325 1.085 76.32 1.3 76.32 1.3 76 1.085 76 1.085 75.995 0.755 75.995 0.755 76 0.54 76 0.54 76.32 0.755 76.32 0.755 76.325 ;
      POLYGON 2.91 68.83 2.91 68.53 1.23 68.53 1.23 68.81 1.78 68.81 1.78 68.83 ;
      POLYGON 103.1 66.79 103.1 66.09 103.19 66.09 103.19 65.81 100.13 65.81 100.13 66.11 102.89 66.11 102.89 66.79 ;
      POLYGON 8.89 7.63 8.89 7.33 1.99 7.33 1.99 6.65 1.78 6.65 1.78 7.35 1.69 7.35 1.69 7.63 ;
      POLYGON 89.405 0.165 89.405 0.16 89.62 0.16 89.62 -0.16 89.405 -0.16 89.405 -0.165 89.075 -0.165 89.075 -0.16 88.86 -0.16 88.86 0.16 89.075 0.16 89.075 0.165 ;
      POLYGON 59.965 0.165 59.965 0.16 60.18 0.16 60.18 -0.16 59.965 -0.16 59.965 -0.165 59.635 -0.165 59.635 -0.16 59.42 -0.16 59.42 0.16 59.635 0.16 59.635 0.165 ;
      POLYGON 30.525 0.165 30.525 0.16 30.74 0.16 30.74 -0.16 30.525 -0.16 30.525 -0.165 30.195 -0.165 30.195 -0.16 29.98 -0.16 29.98 0.16 30.195 0.16 30.195 0.165 ;
      POLYGON 1.085 0.165 1.085 0.16 1.3 0.16 1.3 -0.16 1.085 -0.16 1.085 -0.165 0.755 -0.165 0.755 -0.16 0.54 -0.16 0.54 0.16 0.755 0.16 0.755 0.165 ;
      POLYGON 104.48 75.76 104.48 72.63 103.1 72.63 103.1 71.53 104.48 71.53 104.48 71.27 103.1 71.27 103.1 70.17 104.48 70.17 104.48 69.91 103.1 69.91 103.1 68.81 104.48 68.81 104.48 67.19 103.1 67.19 103.1 66.09 104.48 66.09 104.48 65.83 103.1 65.83 103.1 64.73 104.48 64.73 104.48 64.47 103.1 64.47 103.1 63.37 104.48 63.37 104.48 61.75 103.1 61.75 103.1 60.65 104.48 60.65 104.48 60.39 103.1 60.39 103.1 59.29 104.48 59.29 104.48 59.03 103.1 59.03 103.1 57.93 104.48 57.93 104.48 56.31 103.1 56.31 103.1 55.21 104.48 55.21 104.48 54.95 103.1 54.95 103.1 53.85 104.48 53.85 104.48 53.59 103.1 53.59 103.1 52.49 104.48 52.49 104.48 50.87 103.1 50.87 103.1 49.77 104.48 49.77 104.48 49.51 103.1 49.51 103.1 48.41 104.48 48.41 104.48 48.15 103.1 48.15 103.1 47.05 104.48 47.05 104.48 45.43 103.1 45.43 103.1 44.33 104.48 44.33 104.48 44.07 103.1 44.07 103.1 42.97 104.48 42.97 104.48 42.71 103.1 42.71 103.1 41.61 104.48 41.61 104.48 39.31 103.1 39.31 103.1 38.21 104.48 38.21 104.48 37.95 103.1 37.95 103.1 36.85 104.48 36.85 104.48 34.55 103.1 34.55 103.1 33.45 104.48 33.45 104.48 32.51 103.1 32.51 103.1 31.41 104.48 31.41 104.48 29.11 103.1 29.11 103.1 28.01 104.48 28.01 104.48 27.75 103.1 27.75 103.1 26.65 104.48 26.65 104.48 26.39 103.1 26.39 103.1 25.29 104.48 25.29 104.48 23.67 103.1 23.67 103.1 22.57 104.48 22.57 104.48 22.31 103.1 22.31 103.1 21.21 104.48 21.21 104.48 20.95 103.1 20.95 103.1 19.85 104.48 19.85 104.48 18.23 103.1 18.23 103.1 17.13 104.48 17.13 104.48 16.87 103.1 16.87 103.1 15.77 104.48 15.77 104.48 15.51 103.1 15.51 103.1 14.41 104.48 14.41 104.48 12.79 103.1 12.79 103.1 11.69 104.48 11.69 104.48 11.43 103.1 11.43 103.1 10.33 104.48 10.33 104.48 10.07 103.1 10.07 103.1 8.97 104.48 8.97 104.48 7.35 103.1 7.35 103.1 6.25 104.48 6.25 104.48 5.31 103.1 5.31 103.1 4.21 104.48 4.21 104.48 0.4 0.4 0.4 0.4 3.53 1.78 3.53 1.78 4.63 0.4 4.63 0.4 6.25 1.78 6.25 1.78 7.35 0.4 7.35 0.4 7.61 1.78 7.61 1.78 8.71 0.4 8.71 0.4 8.97 1.78 8.97 1.78 10.07 0.4 10.07 0.4 11.69 1.78 11.69 1.78 12.79 0.4 12.79 0.4 13.05 1.78 13.05 1.78 14.15 0.4 14.15 0.4 14.41 1.78 14.41 1.78 15.51 0.4 15.51 0.4 17.13 1.78 17.13 1.78 18.23 0.4 18.23 0.4 18.49 1.78 18.49 1.78 19.59 0.4 19.59 0.4 19.85 1.78 19.85 1.78 20.95 0.4 20.95 0.4 23.25 1.78 23.25 1.78 24.35 0.4 24.35 0.4 24.61 1.78 24.61 1.78 25.71 0.4 25.71 0.4 28.01 1.78 28.01 1.78 29.11 0.4 29.11 0.4 29.37 1.78 29.37 1.78 30.47 0.4 30.47 0.4 30.73 1.78 30.73 1.78 31.83 0.4 31.83 0.4 33.45 1.78 33.45 1.78 34.55 0.4 34.55 0.4 34.81 1.78 34.81 1.78 35.91 0.4 35.91 0.4 36.17 1.78 36.17 1.78 37.27 0.4 37.27 0.4 38.89 1.78 38.89 1.78 39.99 0.4 39.99 0.4 40.25 1.78 40.25 1.78 41.35 0.4 41.35 0.4 41.61 1.78 41.61 1.78 42.71 0.4 42.71 0.4 44.33 1.78 44.33 1.78 45.43 0.4 45.43 0.4 46.37 1.78 46.37 1.78 47.47 0.4 47.47 0.4 49.77 1.78 49.77 1.78 50.87 0.4 50.87 0.4 51.13 1.78 51.13 1.78 52.23 0.4 52.23 0.4 52.49 1.78 52.49 1.78 53.59 0.4 53.59 0.4 55.21 1.78 55.21 1.78 56.31 0.4 56.31 0.4 56.57 1.78 56.57 1.78 57.67 0.4 57.67 0.4 57.93 1.78 57.93 1.78 59.03 0.4 59.03 0.4 60.65 1.78 60.65 1.78 61.75 0.4 61.75 0.4 62.01 1.78 62.01 1.78 63.11 0.4 63.11 0.4 63.37 1.78 63.37 1.78 64.47 0.4 64.47 0.4 66.09 1.78 66.09 1.78 67.19 0.4 67.19 0.4 67.45 1.78 67.45 1.78 68.55 0.4 68.55 0.4 68.81 1.78 68.81 1.78 69.91 0.4 69.91 0.4 71.53 1.78 71.53 1.78 72.63 0.4 72.63 0.4 75.76 ;
    LAYER met4 ;
      POLYGON 104.26 75.16 104.26 59.87 104.55 59.87 104.55 57.09 104.26 57.09 104.26 19.07 104.55 19.07 104.55 16.29 104.26 16.29 104.26 1 103.66 1 103.66 16.29 103.37 16.29 103.37 19.07 103.66 19.07 103.66 57.09 103.37 57.09 103.37 59.87 103.66 59.87 103.66 75.16 ;
      POLYGON 1.22 75.16 1.22 39.47 1.51 39.47 1.51 36.69 1.22 36.69 1.22 1 0.62 1 0.62 36.69 0.33 36.69 0.33 39.47 0.62 39.47 0.62 75.16 ;
      POLYGON 103.26 75.76 103.26 75.16 104.48 75.16 104.48 1 103.26 1 103.26 0.4 100.83 0.4 100.83 1.76 99.73 1.76 99.73 0.4 89.94 0.4 89.94 1 88.54 1 88.54 0.4 75.22 0.4 75.22 1 73.82 1 73.82 0.4 60.5 0.4 60.5 1 59.1 1 59.1 0.4 45.78 0.4 45.78 1 44.38 1 44.38 0.4 31.06 0.4 31.06 1 29.66 1 29.66 0.4 16.34 0.4 16.34 1 14.94 1 14.94 0.4 5.15 0.4 5.15 1.76 4.05 1.76 4.05 0.4 1.62 0.4 1.62 1 0.4 1 0.4 75.16 1.62 75.16 1.62 75.76 14.94 75.76 14.94 75.16 16.34 75.16 16.34 75.76 29.66 75.76 29.66 75.16 31.06 75.16 31.06 75.76 44.38 75.76 44.38 75.16 45.78 75.16 45.78 75.76 59.1 75.76 59.1 75.16 60.5 75.16 60.5 75.76 73.82 75.76 73.82 75.16 75.22 75.16 75.22 75.76 88.54 75.76 88.54 75.16 89.94 75.16 89.94 75.76 ;
    LAYER met1 ;
      POLYGON 104.6 75.64 104.6 73.96 104.12 73.96 104.12 72.92 104.6 72.92 104.6 71.24 104.12 71.24 104.12 70.2 104.6 70.2 104.6 68.52 104.12 68.52 104.12 67.48 104.6 67.48 104.6 65.8 104.12 65.8 104.12 64.76 104.6 64.76 104.6 63.08 104.12 63.08 104.12 62.04 104.6 62.04 104.6 60.36 104.12 60.36 104.12 59.32 104.6 59.32 104.6 57.64 104.12 57.64 104.12 56.6 104.6 56.6 104.6 54.92 104.12 54.92 104.12 53.88 104.6 53.88 104.6 52.2 104.12 52.2 104.12 51.16 104.6 51.16 104.6 49.48 104.12 49.48 104.12 48.44 104.6 48.44 104.6 46.76 104.12 46.76 104.12 45.72 104.6 45.72 104.6 44.04 104.12 44.04 104.12 43 104.6 43 104.6 41.32 104.12 41.32 104.12 40.28 104.6 40.28 104.6 38.6 104.12 38.6 104.12 37.56 104.6 37.56 104.6 35.88 104.12 35.88 104.12 34.84 104.6 34.84 104.6 33.16 104.12 33.16 104.12 32.12 104.6 32.12 104.6 30.44 104.12 30.44 104.12 29.4 104.6 29.4 104.6 27.72 104.12 27.72 104.12 26.68 104.6 26.68 104.6 25 104.12 25 104.12 23.96 104.6 23.96 104.6 22.28 104.12 22.28 104.12 21.24 104.6 21.24 104.6 19.56 104.12 19.56 104.12 18.52 104.6 18.52 104.6 16.84 104.12 16.84 104.12 15.8 104.6 15.8 104.6 14.12 104.12 14.12 104.12 13.08 104.6 13.08 104.6 11.4 104.12 11.4 104.12 10.36 104.6 10.36 104.6 8.68 104.12 8.68 104.12 7.64 104.6 7.64 104.6 5.96 104.12 5.96 104.12 4.92 104.6 4.92 104.6 3.24 104.12 3.24 104.12 2.2 104.6 2.2 104.6 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 ;
    LAYER met5 ;
      POLYGON 101.68 72.96 101.68 63.28 98.48 63.28 98.48 53.68 101.68 53.68 101.68 42.88 98.48 42.88 98.48 33.28 101.68 33.28 101.68 22.48 98.48 22.48 98.48 12.88 101.68 12.88 101.68 3.2 3.2 3.2 3.2 12.88 6.4 12.88 6.4 22.48 3.2 22.48 3.2 33.28 6.4 33.28 6.4 42.88 3.2 42.88 3.2 53.68 6.4 53.68 6.4 63.28 3.2 63.28 3.2 72.96 ;
    LAYER li1 ;
      RECT 0.34 0.34 104.54 75.82 ;
    LAYER mcon ;
      RECT 104.565 76.075 104.735 76.245 ;
      RECT 104.105 76.075 104.275 76.245 ;
      RECT 103.645 76.075 103.815 76.245 ;
      RECT 103.185 76.075 103.355 76.245 ;
      RECT 102.725 76.075 102.895 76.245 ;
      RECT 102.265 76.075 102.435 76.245 ;
      RECT 101.805 76.075 101.975 76.245 ;
      RECT 101.345 76.075 101.515 76.245 ;
      RECT 100.885 76.075 101.055 76.245 ;
      RECT 100.425 76.075 100.595 76.245 ;
      RECT 99.965 76.075 100.135 76.245 ;
      RECT 99.505 76.075 99.675 76.245 ;
      RECT 99.045 76.075 99.215 76.245 ;
      RECT 98.585 76.075 98.755 76.245 ;
      RECT 98.125 76.075 98.295 76.245 ;
      RECT 97.665 76.075 97.835 76.245 ;
      RECT 97.205 76.075 97.375 76.245 ;
      RECT 96.745 76.075 96.915 76.245 ;
      RECT 96.285 76.075 96.455 76.245 ;
      RECT 95.825 76.075 95.995 76.245 ;
      RECT 95.365 76.075 95.535 76.245 ;
      RECT 94.905 76.075 95.075 76.245 ;
      RECT 94.445 76.075 94.615 76.245 ;
      RECT 93.985 76.075 94.155 76.245 ;
      RECT 93.525 76.075 93.695 76.245 ;
      RECT 93.065 76.075 93.235 76.245 ;
      RECT 92.605 76.075 92.775 76.245 ;
      RECT 92.145 76.075 92.315 76.245 ;
      RECT 91.685 76.075 91.855 76.245 ;
      RECT 91.225 76.075 91.395 76.245 ;
      RECT 90.765 76.075 90.935 76.245 ;
      RECT 90.305 76.075 90.475 76.245 ;
      RECT 89.845 76.075 90.015 76.245 ;
      RECT 89.385 76.075 89.555 76.245 ;
      RECT 88.925 76.075 89.095 76.245 ;
      RECT 88.465 76.075 88.635 76.245 ;
      RECT 88.005 76.075 88.175 76.245 ;
      RECT 87.545 76.075 87.715 76.245 ;
      RECT 87.085 76.075 87.255 76.245 ;
      RECT 86.625 76.075 86.795 76.245 ;
      RECT 86.165 76.075 86.335 76.245 ;
      RECT 85.705 76.075 85.875 76.245 ;
      RECT 85.245 76.075 85.415 76.245 ;
      RECT 84.785 76.075 84.955 76.245 ;
      RECT 84.325 76.075 84.495 76.245 ;
      RECT 83.865 76.075 84.035 76.245 ;
      RECT 83.405 76.075 83.575 76.245 ;
      RECT 82.945 76.075 83.115 76.245 ;
      RECT 82.485 76.075 82.655 76.245 ;
      RECT 82.025 76.075 82.195 76.245 ;
      RECT 81.565 76.075 81.735 76.245 ;
      RECT 81.105 76.075 81.275 76.245 ;
      RECT 80.645 76.075 80.815 76.245 ;
      RECT 80.185 76.075 80.355 76.245 ;
      RECT 79.725 76.075 79.895 76.245 ;
      RECT 79.265 76.075 79.435 76.245 ;
      RECT 78.805 76.075 78.975 76.245 ;
      RECT 78.345 76.075 78.515 76.245 ;
      RECT 77.885 76.075 78.055 76.245 ;
      RECT 77.425 76.075 77.595 76.245 ;
      RECT 76.965 76.075 77.135 76.245 ;
      RECT 76.505 76.075 76.675 76.245 ;
      RECT 76.045 76.075 76.215 76.245 ;
      RECT 75.585 76.075 75.755 76.245 ;
      RECT 75.125 76.075 75.295 76.245 ;
      RECT 74.665 76.075 74.835 76.245 ;
      RECT 74.205 76.075 74.375 76.245 ;
      RECT 73.745 76.075 73.915 76.245 ;
      RECT 73.285 76.075 73.455 76.245 ;
      RECT 72.825 76.075 72.995 76.245 ;
      RECT 72.365 76.075 72.535 76.245 ;
      RECT 71.905 76.075 72.075 76.245 ;
      RECT 71.445 76.075 71.615 76.245 ;
      RECT 70.985 76.075 71.155 76.245 ;
      RECT 70.525 76.075 70.695 76.245 ;
      RECT 70.065 76.075 70.235 76.245 ;
      RECT 69.605 76.075 69.775 76.245 ;
      RECT 69.145 76.075 69.315 76.245 ;
      RECT 68.685 76.075 68.855 76.245 ;
      RECT 68.225 76.075 68.395 76.245 ;
      RECT 67.765 76.075 67.935 76.245 ;
      RECT 67.305 76.075 67.475 76.245 ;
      RECT 66.845 76.075 67.015 76.245 ;
      RECT 66.385 76.075 66.555 76.245 ;
      RECT 65.925 76.075 66.095 76.245 ;
      RECT 65.465 76.075 65.635 76.245 ;
      RECT 65.005 76.075 65.175 76.245 ;
      RECT 64.545 76.075 64.715 76.245 ;
      RECT 64.085 76.075 64.255 76.245 ;
      RECT 63.625 76.075 63.795 76.245 ;
      RECT 63.165 76.075 63.335 76.245 ;
      RECT 62.705 76.075 62.875 76.245 ;
      RECT 62.245 76.075 62.415 76.245 ;
      RECT 61.785 76.075 61.955 76.245 ;
      RECT 61.325 76.075 61.495 76.245 ;
      RECT 60.865 76.075 61.035 76.245 ;
      RECT 60.405 76.075 60.575 76.245 ;
      RECT 59.945 76.075 60.115 76.245 ;
      RECT 59.485 76.075 59.655 76.245 ;
      RECT 59.025 76.075 59.195 76.245 ;
      RECT 58.565 76.075 58.735 76.245 ;
      RECT 58.105 76.075 58.275 76.245 ;
      RECT 57.645 76.075 57.815 76.245 ;
      RECT 57.185 76.075 57.355 76.245 ;
      RECT 56.725 76.075 56.895 76.245 ;
      RECT 56.265 76.075 56.435 76.245 ;
      RECT 55.805 76.075 55.975 76.245 ;
      RECT 55.345 76.075 55.515 76.245 ;
      RECT 54.885 76.075 55.055 76.245 ;
      RECT 54.425 76.075 54.595 76.245 ;
      RECT 53.965 76.075 54.135 76.245 ;
      RECT 53.505 76.075 53.675 76.245 ;
      RECT 53.045 76.075 53.215 76.245 ;
      RECT 52.585 76.075 52.755 76.245 ;
      RECT 52.125 76.075 52.295 76.245 ;
      RECT 51.665 76.075 51.835 76.245 ;
      RECT 51.205 76.075 51.375 76.245 ;
      RECT 50.745 76.075 50.915 76.245 ;
      RECT 50.285 76.075 50.455 76.245 ;
      RECT 49.825 76.075 49.995 76.245 ;
      RECT 49.365 76.075 49.535 76.245 ;
      RECT 48.905 76.075 49.075 76.245 ;
      RECT 48.445 76.075 48.615 76.245 ;
      RECT 47.985 76.075 48.155 76.245 ;
      RECT 47.525 76.075 47.695 76.245 ;
      RECT 47.065 76.075 47.235 76.245 ;
      RECT 46.605 76.075 46.775 76.245 ;
      RECT 46.145 76.075 46.315 76.245 ;
      RECT 45.685 76.075 45.855 76.245 ;
      RECT 45.225 76.075 45.395 76.245 ;
      RECT 44.765 76.075 44.935 76.245 ;
      RECT 44.305 76.075 44.475 76.245 ;
      RECT 43.845 76.075 44.015 76.245 ;
      RECT 43.385 76.075 43.555 76.245 ;
      RECT 42.925 76.075 43.095 76.245 ;
      RECT 42.465 76.075 42.635 76.245 ;
      RECT 42.005 76.075 42.175 76.245 ;
      RECT 41.545 76.075 41.715 76.245 ;
      RECT 41.085 76.075 41.255 76.245 ;
      RECT 40.625 76.075 40.795 76.245 ;
      RECT 40.165 76.075 40.335 76.245 ;
      RECT 39.705 76.075 39.875 76.245 ;
      RECT 39.245 76.075 39.415 76.245 ;
      RECT 38.785 76.075 38.955 76.245 ;
      RECT 38.325 76.075 38.495 76.245 ;
      RECT 37.865 76.075 38.035 76.245 ;
      RECT 37.405 76.075 37.575 76.245 ;
      RECT 36.945 76.075 37.115 76.245 ;
      RECT 36.485 76.075 36.655 76.245 ;
      RECT 36.025 76.075 36.195 76.245 ;
      RECT 35.565 76.075 35.735 76.245 ;
      RECT 35.105 76.075 35.275 76.245 ;
      RECT 34.645 76.075 34.815 76.245 ;
      RECT 34.185 76.075 34.355 76.245 ;
      RECT 33.725 76.075 33.895 76.245 ;
      RECT 33.265 76.075 33.435 76.245 ;
      RECT 32.805 76.075 32.975 76.245 ;
      RECT 32.345 76.075 32.515 76.245 ;
      RECT 31.885 76.075 32.055 76.245 ;
      RECT 31.425 76.075 31.595 76.245 ;
      RECT 30.965 76.075 31.135 76.245 ;
      RECT 30.505 76.075 30.675 76.245 ;
      RECT 30.045 76.075 30.215 76.245 ;
      RECT 29.585 76.075 29.755 76.245 ;
      RECT 29.125 76.075 29.295 76.245 ;
      RECT 28.665 76.075 28.835 76.245 ;
      RECT 28.205 76.075 28.375 76.245 ;
      RECT 27.745 76.075 27.915 76.245 ;
      RECT 27.285 76.075 27.455 76.245 ;
      RECT 26.825 76.075 26.995 76.245 ;
      RECT 26.365 76.075 26.535 76.245 ;
      RECT 25.905 76.075 26.075 76.245 ;
      RECT 25.445 76.075 25.615 76.245 ;
      RECT 24.985 76.075 25.155 76.245 ;
      RECT 24.525 76.075 24.695 76.245 ;
      RECT 24.065 76.075 24.235 76.245 ;
      RECT 23.605 76.075 23.775 76.245 ;
      RECT 23.145 76.075 23.315 76.245 ;
      RECT 22.685 76.075 22.855 76.245 ;
      RECT 22.225 76.075 22.395 76.245 ;
      RECT 21.765 76.075 21.935 76.245 ;
      RECT 21.305 76.075 21.475 76.245 ;
      RECT 20.845 76.075 21.015 76.245 ;
      RECT 20.385 76.075 20.555 76.245 ;
      RECT 19.925 76.075 20.095 76.245 ;
      RECT 19.465 76.075 19.635 76.245 ;
      RECT 19.005 76.075 19.175 76.245 ;
      RECT 18.545 76.075 18.715 76.245 ;
      RECT 18.085 76.075 18.255 76.245 ;
      RECT 17.625 76.075 17.795 76.245 ;
      RECT 17.165 76.075 17.335 76.245 ;
      RECT 16.705 76.075 16.875 76.245 ;
      RECT 16.245 76.075 16.415 76.245 ;
      RECT 15.785 76.075 15.955 76.245 ;
      RECT 15.325 76.075 15.495 76.245 ;
      RECT 14.865 76.075 15.035 76.245 ;
      RECT 14.405 76.075 14.575 76.245 ;
      RECT 13.945 76.075 14.115 76.245 ;
      RECT 13.485 76.075 13.655 76.245 ;
      RECT 13.025 76.075 13.195 76.245 ;
      RECT 12.565 76.075 12.735 76.245 ;
      RECT 12.105 76.075 12.275 76.245 ;
      RECT 11.645 76.075 11.815 76.245 ;
      RECT 11.185 76.075 11.355 76.245 ;
      RECT 10.725 76.075 10.895 76.245 ;
      RECT 10.265 76.075 10.435 76.245 ;
      RECT 9.805 76.075 9.975 76.245 ;
      RECT 9.345 76.075 9.515 76.245 ;
      RECT 8.885 76.075 9.055 76.245 ;
      RECT 8.425 76.075 8.595 76.245 ;
      RECT 7.965 76.075 8.135 76.245 ;
      RECT 7.505 76.075 7.675 76.245 ;
      RECT 7.045 76.075 7.215 76.245 ;
      RECT 6.585 76.075 6.755 76.245 ;
      RECT 6.125 76.075 6.295 76.245 ;
      RECT 5.665 76.075 5.835 76.245 ;
      RECT 5.205 76.075 5.375 76.245 ;
      RECT 4.745 76.075 4.915 76.245 ;
      RECT 4.285 76.075 4.455 76.245 ;
      RECT 3.825 76.075 3.995 76.245 ;
      RECT 3.365 76.075 3.535 76.245 ;
      RECT 2.905 76.075 3.075 76.245 ;
      RECT 2.445 76.075 2.615 76.245 ;
      RECT 1.985 76.075 2.155 76.245 ;
      RECT 1.525 76.075 1.695 76.245 ;
      RECT 1.065 76.075 1.235 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 104.565 73.355 104.735 73.525 ;
      RECT 104.105 73.355 104.275 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 104.565 70.635 104.735 70.805 ;
      RECT 104.105 70.635 104.275 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 104.565 67.915 104.735 68.085 ;
      RECT 104.105 67.915 104.275 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 104.565 65.195 104.735 65.365 ;
      RECT 104.105 65.195 104.275 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 104.565 62.475 104.735 62.645 ;
      RECT 104.105 62.475 104.275 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 104.565 59.755 104.735 59.925 ;
      RECT 104.105 59.755 104.275 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 104.565 57.035 104.735 57.205 ;
      RECT 104.105 57.035 104.275 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 104.565 54.315 104.735 54.485 ;
      RECT 104.105 54.315 104.275 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 104.565 51.595 104.735 51.765 ;
      RECT 104.105 51.595 104.275 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 104.565 48.875 104.735 49.045 ;
      RECT 104.105 48.875 104.275 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 104.565 46.155 104.735 46.325 ;
      RECT 104.105 46.155 104.275 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 104.565 43.435 104.735 43.605 ;
      RECT 104.105 43.435 104.275 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 104.565 40.715 104.735 40.885 ;
      RECT 104.105 40.715 104.275 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 104.565 37.995 104.735 38.165 ;
      RECT 104.105 37.995 104.275 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 104.565 35.275 104.735 35.445 ;
      RECT 104.105 35.275 104.275 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 104.565 32.555 104.735 32.725 ;
      RECT 104.105 32.555 104.275 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 104.565 29.835 104.735 30.005 ;
      RECT 104.105 29.835 104.275 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 104.565 27.115 104.735 27.285 ;
      RECT 104.105 27.115 104.275 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 104.565 24.395 104.735 24.565 ;
      RECT 104.105 24.395 104.275 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 104.565 21.675 104.735 21.845 ;
      RECT 104.105 21.675 104.275 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 104.565 18.955 104.735 19.125 ;
      RECT 104.105 18.955 104.275 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 104.565 16.235 104.735 16.405 ;
      RECT 104.105 16.235 104.275 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 104.565 13.515 104.735 13.685 ;
      RECT 104.105 13.515 104.275 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 104.565 10.795 104.735 10.965 ;
      RECT 104.105 10.795 104.275 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 104.565 8.075 104.735 8.245 ;
      RECT 104.105 8.075 104.275 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 104.565 5.355 104.735 5.525 ;
      RECT 104.105 5.355 104.275 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 104.565 2.635 104.735 2.805 ;
      RECT 104.105 2.635 104.275 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 104.565 -0.085 104.735 0.085 ;
      RECT 104.105 -0.085 104.275 0.085 ;
      RECT 103.645 -0.085 103.815 0.085 ;
      RECT 103.185 -0.085 103.355 0.085 ;
      RECT 102.725 -0.085 102.895 0.085 ;
      RECT 102.265 -0.085 102.435 0.085 ;
      RECT 101.805 -0.085 101.975 0.085 ;
      RECT 101.345 -0.085 101.515 0.085 ;
      RECT 100.885 -0.085 101.055 0.085 ;
      RECT 100.425 -0.085 100.595 0.085 ;
      RECT 99.965 -0.085 100.135 0.085 ;
      RECT 99.505 -0.085 99.675 0.085 ;
      RECT 99.045 -0.085 99.215 0.085 ;
      RECT 98.585 -0.085 98.755 0.085 ;
      RECT 98.125 -0.085 98.295 0.085 ;
      RECT 97.665 -0.085 97.835 0.085 ;
      RECT 97.205 -0.085 97.375 0.085 ;
      RECT 96.745 -0.085 96.915 0.085 ;
      RECT 96.285 -0.085 96.455 0.085 ;
      RECT 95.825 -0.085 95.995 0.085 ;
      RECT 95.365 -0.085 95.535 0.085 ;
      RECT 94.905 -0.085 95.075 0.085 ;
      RECT 94.445 -0.085 94.615 0.085 ;
      RECT 93.985 -0.085 94.155 0.085 ;
      RECT 93.525 -0.085 93.695 0.085 ;
      RECT 93.065 -0.085 93.235 0.085 ;
      RECT 92.605 -0.085 92.775 0.085 ;
      RECT 92.145 -0.085 92.315 0.085 ;
      RECT 91.685 -0.085 91.855 0.085 ;
      RECT 91.225 -0.085 91.395 0.085 ;
      RECT 90.765 -0.085 90.935 0.085 ;
      RECT 90.305 -0.085 90.475 0.085 ;
      RECT 89.845 -0.085 90.015 0.085 ;
      RECT 89.385 -0.085 89.555 0.085 ;
      RECT 88.925 -0.085 89.095 0.085 ;
      RECT 88.465 -0.085 88.635 0.085 ;
      RECT 88.005 -0.085 88.175 0.085 ;
      RECT 87.545 -0.085 87.715 0.085 ;
      RECT 87.085 -0.085 87.255 0.085 ;
      RECT 86.625 -0.085 86.795 0.085 ;
      RECT 86.165 -0.085 86.335 0.085 ;
      RECT 85.705 -0.085 85.875 0.085 ;
      RECT 85.245 -0.085 85.415 0.085 ;
      RECT 84.785 -0.085 84.955 0.085 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 89.165 76.085 89.315 76.235 ;
      RECT 59.725 76.085 59.875 76.235 ;
      RECT 30.285 76.085 30.435 76.235 ;
      RECT 0.845 76.085 0.995 76.235 ;
      RECT 16.025 74.385 16.175 74.535 ;
      RECT 100.665 1.625 100.815 1.775 ;
      RECT 89.165 -0.075 89.315 0.075 ;
      RECT 59.725 -0.075 59.875 0.075 ;
      RECT 30.285 -0.075 30.435 0.075 ;
      RECT 0.845 -0.075 0.995 0.075 ;
    LAYER via2 ;
      RECT 89.14 76.06 89.34 76.26 ;
      RECT 59.7 76.06 59.9 76.26 ;
      RECT 30.26 76.06 30.46 76.26 ;
      RECT 0.82 76.06 1.02 76.26 ;
      RECT 1.28 61.1 1.48 61.3 ;
      RECT 103.4 59.74 103.6 59.94 ;
      RECT 103.4 50.22 103.6 50.42 ;
      RECT 1.28 17.58 1.48 17.78 ;
      RECT 102.94 16.22 103.14 16.42 ;
      RECT 1.74 12.14 1.94 12.34 ;
      RECT 102.94 9.42 103.14 9.62 ;
      RECT 103.4 6.7 103.6 6.9 ;
      RECT 89.14 -0.1 89.34 0.1 ;
      RECT 59.7 -0.1 59.9 0.1 ;
      RECT 30.26 -0.1 30.46 0.1 ;
      RECT 0.82 -0.1 1.02 0.1 ;
    LAYER via3 ;
      RECT 89.14 76.06 89.34 76.26 ;
      RECT 59.7 76.06 59.9 76.26 ;
      RECT 30.26 76.06 30.46 76.26 ;
      RECT 0.82 76.06 1.02 76.26 ;
      RECT 89.14 -0.1 89.34 0.1 ;
      RECT 59.7 -0.1 59.9 0.1 ;
      RECT 30.26 -0.1 30.46 0.1 ;
      RECT 0.82 -0.1 1.02 0.1 ;
    LAYER via4 ;
      RECT 103.56 58.88 104.36 59.68 ;
      RECT 103.56 57.28 104.36 58.08 ;
      RECT 0.52 38.48 1.32 39.28 ;
      RECT 0.52 36.88 1.32 37.68 ;
      RECT 103.56 18.08 104.36 18.88 ;
      RECT 103.56 16.48 104.36 17.28 ;
    LAYER fieldpoly ;
      RECT 0.14 0.14 104.74 76.02 ;
    LAYER diff ;
      RECT 0 0 104.88 76.16 ;
    LAYER nwell ;
      POLYGON 105.07 74.855 105.07 72.025 103.77 72.025 103.77 73.25 102.85 73.25 102.85 74.855 ;
      POLYGON 3.87 74.855 3.87 73.25 2.03 73.25 2.03 72.025 -0.19 72.025 -0.19 74.855 ;
      RECT 103.77 66.585 105.07 69.415 ;
      RECT -0.19 66.585 2.03 69.415 ;
      RECT 103.77 61.145 105.07 63.975 ;
      RECT -0.19 61.145 2.03 63.975 ;
      RECT 103.77 55.705 105.07 58.535 ;
      RECT -0.19 55.705 2.03 58.535 ;
      RECT 103.77 50.265 105.07 53.095 ;
      RECT -0.19 50.265 2.03 53.095 ;
      RECT 103.77 44.825 105.07 47.655 ;
      RECT -0.19 44.825 2.03 47.655 ;
      RECT 103.77 39.385 105.07 42.215 ;
      POLYGON 2.03 42.215 2.03 40.99 3.87 40.99 3.87 39.385 -0.19 39.385 -0.19 42.215 ;
      POLYGON 105.07 36.775 105.07 33.945 104.23 33.945 104.23 35.17 103.77 35.17 103.77 36.775 ;
      RECT -0.19 33.945 2.03 36.775 ;
      POLYGON 105.07 31.335 105.07 28.505 103.77 28.505 103.77 30.11 104.23 30.11 104.23 31.335 ;
      RECT -0.19 28.505 2.03 31.335 ;
      POLYGON 105.07 25.895 105.07 23.065 102.85 23.065 102.85 24.67 103.77 24.67 103.77 25.895 ;
      RECT -0.19 23.065 2.03 25.895 ;
      RECT 103.77 17.625 105.07 20.455 ;
      RECT -0.19 17.625 2.03 20.455 ;
      RECT 103.77 12.185 105.07 15.015 ;
      RECT -0.19 12.185 2.03 15.015 ;
      RECT 103.77 6.745 105.07 9.575 ;
      RECT -0.19 6.745 2.03 9.575 ;
      POLYGON 105.07 4.135 105.07 1.305 102.85 1.305 102.85 2.91 103.77 2.91 103.77 4.135 ;
      POLYGON 2.03 4.135 2.03 2.91 3.87 2.91 3.87 1.305 -0.19 1.305 -0.19 4.135 ;
      RECT 0 0 104.88 76.16 ;
    LAYER pwell ;
      RECT 99.49 76.11 99.71 76.28 ;
      RECT 95.81 76.11 96.03 76.28 ;
      RECT 92.13 76.11 92.35 76.28 ;
      RECT 88.45 76.11 88.67 76.28 ;
      RECT 84.77 76.11 84.99 76.28 ;
      RECT 81.09 76.11 81.31 76.28 ;
      RECT 77.41 76.11 77.63 76.28 ;
      RECT 73.73 76.11 73.95 76.28 ;
      RECT 70.05 76.11 70.27 76.28 ;
      RECT 66.37 76.11 66.59 76.28 ;
      RECT 62.69 76.11 62.91 76.28 ;
      RECT 59.01 76.11 59.23 76.28 ;
      RECT 55.33 76.11 55.55 76.28 ;
      RECT 51.65 76.11 51.87 76.28 ;
      RECT 47.97 76.11 48.19 76.28 ;
      RECT 44.29 76.11 44.51 76.28 ;
      RECT 40.61 76.11 40.83 76.28 ;
      RECT 36.93 76.11 37.15 76.28 ;
      RECT 33.25 76.11 33.47 76.28 ;
      RECT 29.57 76.11 29.79 76.28 ;
      RECT 25.89 76.11 26.11 76.28 ;
      RECT 22.21 76.11 22.43 76.28 ;
      RECT 18.53 76.11 18.75 76.28 ;
      RECT 14.85 76.11 15.07 76.28 ;
      RECT 11.17 76.11 11.39 76.28 ;
      RECT 7.49 76.11 7.71 76.28 ;
      RECT 3.81 76.11 4.03 76.28 ;
      RECT 0.13 76.11 0.35 76.28 ;
      RECT 103.215 76.1 103.325 76.22 ;
      RECT 103.215 -0.06 103.325 0.06 ;
      RECT 99.49 -0.12 99.71 0.05 ;
      RECT 95.81 -0.12 96.03 0.05 ;
      RECT 92.13 -0.12 92.35 0.05 ;
      RECT 88.45 -0.12 88.67 0.05 ;
      RECT 84.77 -0.12 84.99 0.05 ;
      RECT 81.09 -0.12 81.31 0.05 ;
      RECT 77.41 -0.12 77.63 0.05 ;
      RECT 73.73 -0.12 73.95 0.05 ;
      RECT 70.05 -0.12 70.27 0.05 ;
      RECT 66.37 -0.12 66.59 0.05 ;
      RECT 62.69 -0.12 62.91 0.05 ;
      RECT 59.01 -0.12 59.23 0.05 ;
      RECT 55.33 -0.12 55.55 0.05 ;
      RECT 51.65 -0.12 51.87 0.05 ;
      RECT 47.97 -0.12 48.19 0.05 ;
      RECT 44.29 -0.12 44.51 0.05 ;
      RECT 40.61 -0.12 40.83 0.05 ;
      RECT 36.93 -0.12 37.15 0.05 ;
      RECT 33.25 -0.12 33.47 0.05 ;
      RECT 29.57 -0.12 29.79 0.05 ;
      RECT 25.89 -0.12 26.11 0.05 ;
      RECT 22.21 -0.12 22.43 0.05 ;
      RECT 18.53 -0.12 18.75 0.05 ;
      RECT 14.85 -0.12 15.07 0.05 ;
      RECT 11.17 -0.12 11.39 0.05 ;
      RECT 7.49 -0.12 7.71 0.05 ;
      RECT 3.81 -0.12 4.03 0.05 ;
      RECT 0.13 -0.12 0.35 0.05 ;
      RECT 0 0 104.88 76.16 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 76.16 104.88 76.16 104.88 0 ;
  END
END cbx_1__1_

END LIBRARY
