

module fpga_core
( prog_clk, Test_en, IO_ISOL_N, clk, gfpga_pad_EMBEDDED_IO_HD_SOC_IN, gfpga_pad_EMBEDDED_IO_HD_SOC_OUT, gfpga_pad_EMBEDDED_IO_HD_SOC_DIR, ccff_head, ccff_tail, sc_head, sc_tail ); 
  input [0:0] prog_clk;
  input [0:0] Test_en;
  input [0:0] IO_ISOL_N;
  input [0:0] clk;
  input [0:143] gfpga_pad_EMBEDDED_IO_HD_SOC_IN;
  output [0:143] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT;
  output [0:143] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR;
  input [0:0] ccff_head;
  output [0:0] ccff_tail;
  input sc_head;
  output sc_tail;

  wire [0:0] cbx_1__0__0_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__0_ccff_tail;
  wire [0:19] cbx_1__0__0_chanx_left_out;
  wire [0:19] cbx_1__0__0_chanx_right_out;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__10_ccff_tail;
  wire [0:19] cbx_1__0__10_chanx_left_out;
  wire [0:19] cbx_1__0__10_chanx_right_out;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__11_ccff_tail;
  wire [0:19] cbx_1__0__11_chanx_left_out;
  wire [0:19] cbx_1__0__11_chanx_right_out;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__1_ccff_tail;
  wire [0:19] cbx_1__0__1_chanx_left_out;
  wire [0:19] cbx_1__0__1_chanx_right_out;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__2_ccff_tail;
  wire [0:19] cbx_1__0__2_chanx_left_out;
  wire [0:19] cbx_1__0__2_chanx_right_out;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__3_ccff_tail;
  wire [0:19] cbx_1__0__3_chanx_left_out;
  wire [0:19] cbx_1__0__3_chanx_right_out;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__4_ccff_tail;
  wire [0:19] cbx_1__0__4_chanx_left_out;
  wire [0:19] cbx_1__0__4_chanx_right_out;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__5_ccff_tail;
  wire [0:19] cbx_1__0__5_chanx_left_out;
  wire [0:19] cbx_1__0__5_chanx_right_out;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__6_ccff_tail;
  wire [0:19] cbx_1__0__6_chanx_left_out;
  wire [0:19] cbx_1__0__6_chanx_right_out;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__7_ccff_tail;
  wire [0:19] cbx_1__0__7_chanx_left_out;
  wire [0:19] cbx_1__0__7_chanx_right_out;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__8_ccff_tail;
  wire [0:19] cbx_1__0__8_chanx_left_out;
  wire [0:19] cbx_1__0__8_chanx_right_out;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__9_ccff_tail;
  wire [0:19] cbx_1__0__9_chanx_left_out;
  wire [0:19] cbx_1__0__9_chanx_right_out;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__0_ccff_tail;
  wire [0:19] cbx_1__12__0_chanx_left_out;
  wire [0:19] cbx_1__12__0_chanx_right_out;
  wire [0:0] cbx_1__12__0_top_grid_pin_0_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__10_ccff_tail;
  wire [0:19] cbx_1__12__10_chanx_left_out;
  wire [0:19] cbx_1__12__10_chanx_right_out;
  wire [0:0] cbx_1__12__10_top_grid_pin_0_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__11_ccff_tail;
  wire [0:19] cbx_1__12__11_chanx_left_out;
  wire [0:19] cbx_1__12__11_chanx_right_out;
  wire [0:0] cbx_1__12__11_top_grid_pin_0_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__1_ccff_tail;
  wire [0:19] cbx_1__12__1_chanx_left_out;
  wire [0:19] cbx_1__12__1_chanx_right_out;
  wire [0:0] cbx_1__12__1_top_grid_pin_0_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__2_ccff_tail;
  wire [0:19] cbx_1__12__2_chanx_left_out;
  wire [0:19] cbx_1__12__2_chanx_right_out;
  wire [0:0] cbx_1__12__2_top_grid_pin_0_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__3_ccff_tail;
  wire [0:19] cbx_1__12__3_chanx_left_out;
  wire [0:19] cbx_1__12__3_chanx_right_out;
  wire [0:0] cbx_1__12__3_top_grid_pin_0_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__4_ccff_tail;
  wire [0:19] cbx_1__12__4_chanx_left_out;
  wire [0:19] cbx_1__12__4_chanx_right_out;
  wire [0:0] cbx_1__12__4_top_grid_pin_0_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__5_ccff_tail;
  wire [0:19] cbx_1__12__5_chanx_left_out;
  wire [0:19] cbx_1__12__5_chanx_right_out;
  wire [0:0] cbx_1__12__5_top_grid_pin_0_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__6_ccff_tail;
  wire [0:19] cbx_1__12__6_chanx_left_out;
  wire [0:19] cbx_1__12__6_chanx_right_out;
  wire [0:0] cbx_1__12__6_top_grid_pin_0_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__7_ccff_tail;
  wire [0:19] cbx_1__12__7_chanx_left_out;
  wire [0:19] cbx_1__12__7_chanx_right_out;
  wire [0:0] cbx_1__12__7_top_grid_pin_0_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__8_ccff_tail;
  wire [0:19] cbx_1__12__8_chanx_left_out;
  wire [0:19] cbx_1__12__8_chanx_right_out;
  wire [0:0] cbx_1__12__8_top_grid_pin_0_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__9_ccff_tail;
  wire [0:19] cbx_1__12__9_chanx_left_out;
  wire [0:19] cbx_1__12__9_chanx_right_out;
  wire [0:0] cbx_1__12__9_top_grid_pin_0_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__0_ccff_tail;
  wire [0:19] cbx_1__1__0_chanx_left_out;
  wire [0:19] cbx_1__1__0_chanx_right_out;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__100_ccff_tail;
  wire [0:19] cbx_1__1__100_chanx_left_out;
  wire [0:19] cbx_1__1__100_chanx_right_out;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__101_ccff_tail;
  wire [0:19] cbx_1__1__101_chanx_left_out;
  wire [0:19] cbx_1__1__101_chanx_right_out;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__102_ccff_tail;
  wire [0:19] cbx_1__1__102_chanx_left_out;
  wire [0:19] cbx_1__1__102_chanx_right_out;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__103_ccff_tail;
  wire [0:19] cbx_1__1__103_chanx_left_out;
  wire [0:19] cbx_1__1__103_chanx_right_out;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__104_ccff_tail;
  wire [0:19] cbx_1__1__104_chanx_left_out;
  wire [0:19] cbx_1__1__104_chanx_right_out;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__105_ccff_tail;
  wire [0:19] cbx_1__1__105_chanx_left_out;
  wire [0:19] cbx_1__1__105_chanx_right_out;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__106_ccff_tail;
  wire [0:19] cbx_1__1__106_chanx_left_out;
  wire [0:19] cbx_1__1__106_chanx_right_out;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__107_ccff_tail;
  wire [0:19] cbx_1__1__107_chanx_left_out;
  wire [0:19] cbx_1__1__107_chanx_right_out;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__108_ccff_tail;
  wire [0:19] cbx_1__1__108_chanx_left_out;
  wire [0:19] cbx_1__1__108_chanx_right_out;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__109_ccff_tail;
  wire [0:19] cbx_1__1__109_chanx_left_out;
  wire [0:19] cbx_1__1__109_chanx_right_out;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__10_ccff_tail;
  wire [0:19] cbx_1__1__10_chanx_left_out;
  wire [0:19] cbx_1__1__10_chanx_right_out;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__110_ccff_tail;
  wire [0:19] cbx_1__1__110_chanx_left_out;
  wire [0:19] cbx_1__1__110_chanx_right_out;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__111_ccff_tail;
  wire [0:19] cbx_1__1__111_chanx_left_out;
  wire [0:19] cbx_1__1__111_chanx_right_out;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__112_ccff_tail;
  wire [0:19] cbx_1__1__112_chanx_left_out;
  wire [0:19] cbx_1__1__112_chanx_right_out;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__113_ccff_tail;
  wire [0:19] cbx_1__1__113_chanx_left_out;
  wire [0:19] cbx_1__1__113_chanx_right_out;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__114_ccff_tail;
  wire [0:19] cbx_1__1__114_chanx_left_out;
  wire [0:19] cbx_1__1__114_chanx_right_out;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__115_ccff_tail;
  wire [0:19] cbx_1__1__115_chanx_left_out;
  wire [0:19] cbx_1__1__115_chanx_right_out;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__116_ccff_tail;
  wire [0:19] cbx_1__1__116_chanx_left_out;
  wire [0:19] cbx_1__1__116_chanx_right_out;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__117_ccff_tail;
  wire [0:19] cbx_1__1__117_chanx_left_out;
  wire [0:19] cbx_1__1__117_chanx_right_out;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__118_ccff_tail;
  wire [0:19] cbx_1__1__118_chanx_left_out;
  wire [0:19] cbx_1__1__118_chanx_right_out;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__119_ccff_tail;
  wire [0:19] cbx_1__1__119_chanx_left_out;
  wire [0:19] cbx_1__1__119_chanx_right_out;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__11_ccff_tail;
  wire [0:19] cbx_1__1__11_chanx_left_out;
  wire [0:19] cbx_1__1__11_chanx_right_out;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__120_ccff_tail;
  wire [0:19] cbx_1__1__120_chanx_left_out;
  wire [0:19] cbx_1__1__120_chanx_right_out;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__121_ccff_tail;
  wire [0:19] cbx_1__1__121_chanx_left_out;
  wire [0:19] cbx_1__1__121_chanx_right_out;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__122_ccff_tail;
  wire [0:19] cbx_1__1__122_chanx_left_out;
  wire [0:19] cbx_1__1__122_chanx_right_out;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__123_ccff_tail;
  wire [0:19] cbx_1__1__123_chanx_left_out;
  wire [0:19] cbx_1__1__123_chanx_right_out;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__124_ccff_tail;
  wire [0:19] cbx_1__1__124_chanx_left_out;
  wire [0:19] cbx_1__1__124_chanx_right_out;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__125_ccff_tail;
  wire [0:19] cbx_1__1__125_chanx_left_out;
  wire [0:19] cbx_1__1__125_chanx_right_out;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__126_ccff_tail;
  wire [0:19] cbx_1__1__126_chanx_left_out;
  wire [0:19] cbx_1__1__126_chanx_right_out;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__127_ccff_tail;
  wire [0:19] cbx_1__1__127_chanx_left_out;
  wire [0:19] cbx_1__1__127_chanx_right_out;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__128_ccff_tail;
  wire [0:19] cbx_1__1__128_chanx_left_out;
  wire [0:19] cbx_1__1__128_chanx_right_out;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__129_ccff_tail;
  wire [0:19] cbx_1__1__129_chanx_left_out;
  wire [0:19] cbx_1__1__129_chanx_right_out;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__12_ccff_tail;
  wire [0:19] cbx_1__1__12_chanx_left_out;
  wire [0:19] cbx_1__1__12_chanx_right_out;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__130_ccff_tail;
  wire [0:19] cbx_1__1__130_chanx_left_out;
  wire [0:19] cbx_1__1__130_chanx_right_out;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__131_ccff_tail;
  wire [0:19] cbx_1__1__131_chanx_left_out;
  wire [0:19] cbx_1__1__131_chanx_right_out;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__13_ccff_tail;
  wire [0:19] cbx_1__1__13_chanx_left_out;
  wire [0:19] cbx_1__1__13_chanx_right_out;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__14_ccff_tail;
  wire [0:19] cbx_1__1__14_chanx_left_out;
  wire [0:19] cbx_1__1__14_chanx_right_out;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__15_ccff_tail;
  wire [0:19] cbx_1__1__15_chanx_left_out;
  wire [0:19] cbx_1__1__15_chanx_right_out;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__16_ccff_tail;
  wire [0:19] cbx_1__1__16_chanx_left_out;
  wire [0:19] cbx_1__1__16_chanx_right_out;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__17_ccff_tail;
  wire [0:19] cbx_1__1__17_chanx_left_out;
  wire [0:19] cbx_1__1__17_chanx_right_out;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__18_ccff_tail;
  wire [0:19] cbx_1__1__18_chanx_left_out;
  wire [0:19] cbx_1__1__18_chanx_right_out;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__19_ccff_tail;
  wire [0:19] cbx_1__1__19_chanx_left_out;
  wire [0:19] cbx_1__1__19_chanx_right_out;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__1_ccff_tail;
  wire [0:19] cbx_1__1__1_chanx_left_out;
  wire [0:19] cbx_1__1__1_chanx_right_out;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__20_ccff_tail;
  wire [0:19] cbx_1__1__20_chanx_left_out;
  wire [0:19] cbx_1__1__20_chanx_right_out;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__21_ccff_tail;
  wire [0:19] cbx_1__1__21_chanx_left_out;
  wire [0:19] cbx_1__1__21_chanx_right_out;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__22_ccff_tail;
  wire [0:19] cbx_1__1__22_chanx_left_out;
  wire [0:19] cbx_1__1__22_chanx_right_out;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__23_ccff_tail;
  wire [0:19] cbx_1__1__23_chanx_left_out;
  wire [0:19] cbx_1__1__23_chanx_right_out;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__24_ccff_tail;
  wire [0:19] cbx_1__1__24_chanx_left_out;
  wire [0:19] cbx_1__1__24_chanx_right_out;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__25_ccff_tail;
  wire [0:19] cbx_1__1__25_chanx_left_out;
  wire [0:19] cbx_1__1__25_chanx_right_out;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__26_ccff_tail;
  wire [0:19] cbx_1__1__26_chanx_left_out;
  wire [0:19] cbx_1__1__26_chanx_right_out;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__27_ccff_tail;
  wire [0:19] cbx_1__1__27_chanx_left_out;
  wire [0:19] cbx_1__1__27_chanx_right_out;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__28_ccff_tail;
  wire [0:19] cbx_1__1__28_chanx_left_out;
  wire [0:19] cbx_1__1__28_chanx_right_out;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__29_ccff_tail;
  wire [0:19] cbx_1__1__29_chanx_left_out;
  wire [0:19] cbx_1__1__29_chanx_right_out;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__2_ccff_tail;
  wire [0:19] cbx_1__1__2_chanx_left_out;
  wire [0:19] cbx_1__1__2_chanx_right_out;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__30_ccff_tail;
  wire [0:19] cbx_1__1__30_chanx_left_out;
  wire [0:19] cbx_1__1__30_chanx_right_out;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__31_ccff_tail;
  wire [0:19] cbx_1__1__31_chanx_left_out;
  wire [0:19] cbx_1__1__31_chanx_right_out;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__32_ccff_tail;
  wire [0:19] cbx_1__1__32_chanx_left_out;
  wire [0:19] cbx_1__1__32_chanx_right_out;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__33_ccff_tail;
  wire [0:19] cbx_1__1__33_chanx_left_out;
  wire [0:19] cbx_1__1__33_chanx_right_out;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__34_ccff_tail;
  wire [0:19] cbx_1__1__34_chanx_left_out;
  wire [0:19] cbx_1__1__34_chanx_right_out;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__35_ccff_tail;
  wire [0:19] cbx_1__1__35_chanx_left_out;
  wire [0:19] cbx_1__1__35_chanx_right_out;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__36_ccff_tail;
  wire [0:19] cbx_1__1__36_chanx_left_out;
  wire [0:19] cbx_1__1__36_chanx_right_out;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__37_ccff_tail;
  wire [0:19] cbx_1__1__37_chanx_left_out;
  wire [0:19] cbx_1__1__37_chanx_right_out;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__38_ccff_tail;
  wire [0:19] cbx_1__1__38_chanx_left_out;
  wire [0:19] cbx_1__1__38_chanx_right_out;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__39_ccff_tail;
  wire [0:19] cbx_1__1__39_chanx_left_out;
  wire [0:19] cbx_1__1__39_chanx_right_out;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__3_ccff_tail;
  wire [0:19] cbx_1__1__3_chanx_left_out;
  wire [0:19] cbx_1__1__3_chanx_right_out;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__40_ccff_tail;
  wire [0:19] cbx_1__1__40_chanx_left_out;
  wire [0:19] cbx_1__1__40_chanx_right_out;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__41_ccff_tail;
  wire [0:19] cbx_1__1__41_chanx_left_out;
  wire [0:19] cbx_1__1__41_chanx_right_out;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__42_ccff_tail;
  wire [0:19] cbx_1__1__42_chanx_left_out;
  wire [0:19] cbx_1__1__42_chanx_right_out;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__43_ccff_tail;
  wire [0:19] cbx_1__1__43_chanx_left_out;
  wire [0:19] cbx_1__1__43_chanx_right_out;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__44_ccff_tail;
  wire [0:19] cbx_1__1__44_chanx_left_out;
  wire [0:19] cbx_1__1__44_chanx_right_out;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__45_ccff_tail;
  wire [0:19] cbx_1__1__45_chanx_left_out;
  wire [0:19] cbx_1__1__45_chanx_right_out;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__46_ccff_tail;
  wire [0:19] cbx_1__1__46_chanx_left_out;
  wire [0:19] cbx_1__1__46_chanx_right_out;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__47_ccff_tail;
  wire [0:19] cbx_1__1__47_chanx_left_out;
  wire [0:19] cbx_1__1__47_chanx_right_out;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__48_ccff_tail;
  wire [0:19] cbx_1__1__48_chanx_left_out;
  wire [0:19] cbx_1__1__48_chanx_right_out;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__49_ccff_tail;
  wire [0:19] cbx_1__1__49_chanx_left_out;
  wire [0:19] cbx_1__1__49_chanx_right_out;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__4_ccff_tail;
  wire [0:19] cbx_1__1__4_chanx_left_out;
  wire [0:19] cbx_1__1__4_chanx_right_out;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__50_ccff_tail;
  wire [0:19] cbx_1__1__50_chanx_left_out;
  wire [0:19] cbx_1__1__50_chanx_right_out;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__51_ccff_tail;
  wire [0:19] cbx_1__1__51_chanx_left_out;
  wire [0:19] cbx_1__1__51_chanx_right_out;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__52_ccff_tail;
  wire [0:19] cbx_1__1__52_chanx_left_out;
  wire [0:19] cbx_1__1__52_chanx_right_out;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__53_ccff_tail;
  wire [0:19] cbx_1__1__53_chanx_left_out;
  wire [0:19] cbx_1__1__53_chanx_right_out;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__54_ccff_tail;
  wire [0:19] cbx_1__1__54_chanx_left_out;
  wire [0:19] cbx_1__1__54_chanx_right_out;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__55_ccff_tail;
  wire [0:19] cbx_1__1__55_chanx_left_out;
  wire [0:19] cbx_1__1__55_chanx_right_out;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__56_ccff_tail;
  wire [0:19] cbx_1__1__56_chanx_left_out;
  wire [0:19] cbx_1__1__56_chanx_right_out;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__57_ccff_tail;
  wire [0:19] cbx_1__1__57_chanx_left_out;
  wire [0:19] cbx_1__1__57_chanx_right_out;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__58_ccff_tail;
  wire [0:19] cbx_1__1__58_chanx_left_out;
  wire [0:19] cbx_1__1__58_chanx_right_out;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__59_ccff_tail;
  wire [0:19] cbx_1__1__59_chanx_left_out;
  wire [0:19] cbx_1__1__59_chanx_right_out;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__5_ccff_tail;
  wire [0:19] cbx_1__1__5_chanx_left_out;
  wire [0:19] cbx_1__1__5_chanx_right_out;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__60_ccff_tail;
  wire [0:19] cbx_1__1__60_chanx_left_out;
  wire [0:19] cbx_1__1__60_chanx_right_out;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__61_ccff_tail;
  wire [0:19] cbx_1__1__61_chanx_left_out;
  wire [0:19] cbx_1__1__61_chanx_right_out;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__62_ccff_tail;
  wire [0:19] cbx_1__1__62_chanx_left_out;
  wire [0:19] cbx_1__1__62_chanx_right_out;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__63_ccff_tail;
  wire [0:19] cbx_1__1__63_chanx_left_out;
  wire [0:19] cbx_1__1__63_chanx_right_out;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__64_ccff_tail;
  wire [0:19] cbx_1__1__64_chanx_left_out;
  wire [0:19] cbx_1__1__64_chanx_right_out;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__65_ccff_tail;
  wire [0:19] cbx_1__1__65_chanx_left_out;
  wire [0:19] cbx_1__1__65_chanx_right_out;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__66_ccff_tail;
  wire [0:19] cbx_1__1__66_chanx_left_out;
  wire [0:19] cbx_1__1__66_chanx_right_out;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__67_ccff_tail;
  wire [0:19] cbx_1__1__67_chanx_left_out;
  wire [0:19] cbx_1__1__67_chanx_right_out;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__68_ccff_tail;
  wire [0:19] cbx_1__1__68_chanx_left_out;
  wire [0:19] cbx_1__1__68_chanx_right_out;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__69_ccff_tail;
  wire [0:19] cbx_1__1__69_chanx_left_out;
  wire [0:19] cbx_1__1__69_chanx_right_out;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__6_ccff_tail;
  wire [0:19] cbx_1__1__6_chanx_left_out;
  wire [0:19] cbx_1__1__6_chanx_right_out;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__70_ccff_tail;
  wire [0:19] cbx_1__1__70_chanx_left_out;
  wire [0:19] cbx_1__1__70_chanx_right_out;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__71_ccff_tail;
  wire [0:19] cbx_1__1__71_chanx_left_out;
  wire [0:19] cbx_1__1__71_chanx_right_out;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__72_ccff_tail;
  wire [0:19] cbx_1__1__72_chanx_left_out;
  wire [0:19] cbx_1__1__72_chanx_right_out;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__73_ccff_tail;
  wire [0:19] cbx_1__1__73_chanx_left_out;
  wire [0:19] cbx_1__1__73_chanx_right_out;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__74_ccff_tail;
  wire [0:19] cbx_1__1__74_chanx_left_out;
  wire [0:19] cbx_1__1__74_chanx_right_out;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__75_ccff_tail;
  wire [0:19] cbx_1__1__75_chanx_left_out;
  wire [0:19] cbx_1__1__75_chanx_right_out;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__76_ccff_tail;
  wire [0:19] cbx_1__1__76_chanx_left_out;
  wire [0:19] cbx_1__1__76_chanx_right_out;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__77_ccff_tail;
  wire [0:19] cbx_1__1__77_chanx_left_out;
  wire [0:19] cbx_1__1__77_chanx_right_out;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__78_ccff_tail;
  wire [0:19] cbx_1__1__78_chanx_left_out;
  wire [0:19] cbx_1__1__78_chanx_right_out;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__79_ccff_tail;
  wire [0:19] cbx_1__1__79_chanx_left_out;
  wire [0:19] cbx_1__1__79_chanx_right_out;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__7_ccff_tail;
  wire [0:19] cbx_1__1__7_chanx_left_out;
  wire [0:19] cbx_1__1__7_chanx_right_out;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__80_ccff_tail;
  wire [0:19] cbx_1__1__80_chanx_left_out;
  wire [0:19] cbx_1__1__80_chanx_right_out;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__81_ccff_tail;
  wire [0:19] cbx_1__1__81_chanx_left_out;
  wire [0:19] cbx_1__1__81_chanx_right_out;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__82_ccff_tail;
  wire [0:19] cbx_1__1__82_chanx_left_out;
  wire [0:19] cbx_1__1__82_chanx_right_out;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__83_ccff_tail;
  wire [0:19] cbx_1__1__83_chanx_left_out;
  wire [0:19] cbx_1__1__83_chanx_right_out;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__84_ccff_tail;
  wire [0:19] cbx_1__1__84_chanx_left_out;
  wire [0:19] cbx_1__1__84_chanx_right_out;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__85_ccff_tail;
  wire [0:19] cbx_1__1__85_chanx_left_out;
  wire [0:19] cbx_1__1__85_chanx_right_out;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__86_ccff_tail;
  wire [0:19] cbx_1__1__86_chanx_left_out;
  wire [0:19] cbx_1__1__86_chanx_right_out;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__87_ccff_tail;
  wire [0:19] cbx_1__1__87_chanx_left_out;
  wire [0:19] cbx_1__1__87_chanx_right_out;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__88_ccff_tail;
  wire [0:19] cbx_1__1__88_chanx_left_out;
  wire [0:19] cbx_1__1__88_chanx_right_out;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__89_ccff_tail;
  wire [0:19] cbx_1__1__89_chanx_left_out;
  wire [0:19] cbx_1__1__89_chanx_right_out;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__8_ccff_tail;
  wire [0:19] cbx_1__1__8_chanx_left_out;
  wire [0:19] cbx_1__1__8_chanx_right_out;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__90_ccff_tail;
  wire [0:19] cbx_1__1__90_chanx_left_out;
  wire [0:19] cbx_1__1__90_chanx_right_out;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__91_ccff_tail;
  wire [0:19] cbx_1__1__91_chanx_left_out;
  wire [0:19] cbx_1__1__91_chanx_right_out;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__92_ccff_tail;
  wire [0:19] cbx_1__1__92_chanx_left_out;
  wire [0:19] cbx_1__1__92_chanx_right_out;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__93_ccff_tail;
  wire [0:19] cbx_1__1__93_chanx_left_out;
  wire [0:19] cbx_1__1__93_chanx_right_out;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__94_ccff_tail;
  wire [0:19] cbx_1__1__94_chanx_left_out;
  wire [0:19] cbx_1__1__94_chanx_right_out;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__95_ccff_tail;
  wire [0:19] cbx_1__1__95_chanx_left_out;
  wire [0:19] cbx_1__1__95_chanx_right_out;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__96_ccff_tail;
  wire [0:19] cbx_1__1__96_chanx_left_out;
  wire [0:19] cbx_1__1__96_chanx_right_out;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__97_ccff_tail;
  wire [0:19] cbx_1__1__97_chanx_left_out;
  wire [0:19] cbx_1__1__97_chanx_right_out;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__98_ccff_tail;
  wire [0:19] cbx_1__1__98_chanx_left_out;
  wire [0:19] cbx_1__1__98_chanx_right_out;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__99_ccff_tail;
  wire [0:19] cbx_1__1__99_chanx_left_out;
  wire [0:19] cbx_1__1__99_chanx_right_out;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__9_ccff_tail;
  wire [0:19] cbx_1__1__9_chanx_left_out;
  wire [0:19] cbx_1__1__9_chanx_right_out;
  wire [0:0] cby_0__1__0_ccff_tail;
  wire [0:19] cby_0__1__0_chany_bottom_out;
  wire [0:19] cby_0__1__0_chany_top_out;
  wire [0:0] cby_0__1__0_left_grid_pin_0_;
  wire [0:0] cby_0__1__10_ccff_tail;
  wire [0:19] cby_0__1__10_chany_bottom_out;
  wire [0:19] cby_0__1__10_chany_top_out;
  wire [0:0] cby_0__1__10_left_grid_pin_0_;
  wire [0:0] cby_0__1__11_ccff_tail;
  wire [0:19] cby_0__1__11_chany_bottom_out;
  wire [0:19] cby_0__1__11_chany_top_out;
  wire [0:0] cby_0__1__11_left_grid_pin_0_;
  wire [0:0] cby_0__1__1_ccff_tail;
  wire [0:19] cby_0__1__1_chany_bottom_out;
  wire [0:19] cby_0__1__1_chany_top_out;
  wire [0:0] cby_0__1__1_left_grid_pin_0_;
  wire [0:0] cby_0__1__2_ccff_tail;
  wire [0:19] cby_0__1__2_chany_bottom_out;
  wire [0:19] cby_0__1__2_chany_top_out;
  wire [0:0] cby_0__1__2_left_grid_pin_0_;
  wire [0:0] cby_0__1__3_ccff_tail;
  wire [0:19] cby_0__1__3_chany_bottom_out;
  wire [0:19] cby_0__1__3_chany_top_out;
  wire [0:0] cby_0__1__3_left_grid_pin_0_;
  wire [0:0] cby_0__1__4_ccff_tail;
  wire [0:19] cby_0__1__4_chany_bottom_out;
  wire [0:19] cby_0__1__4_chany_top_out;
  wire [0:0] cby_0__1__4_left_grid_pin_0_;
  wire [0:0] cby_0__1__5_ccff_tail;
  wire [0:19] cby_0__1__5_chany_bottom_out;
  wire [0:19] cby_0__1__5_chany_top_out;
  wire [0:0] cby_0__1__5_left_grid_pin_0_;
  wire [0:0] cby_0__1__6_ccff_tail;
  wire [0:19] cby_0__1__6_chany_bottom_out;
  wire [0:19] cby_0__1__6_chany_top_out;
  wire [0:0] cby_0__1__6_left_grid_pin_0_;
  wire [0:0] cby_0__1__7_ccff_tail;
  wire [0:19] cby_0__1__7_chany_bottom_out;
  wire [0:19] cby_0__1__7_chany_top_out;
  wire [0:0] cby_0__1__7_left_grid_pin_0_;
  wire [0:0] cby_0__1__8_ccff_tail;
  wire [0:19] cby_0__1__8_chany_bottom_out;
  wire [0:19] cby_0__1__8_chany_top_out;
  wire [0:0] cby_0__1__8_left_grid_pin_0_;
  wire [0:0] cby_0__1__9_ccff_tail;
  wire [0:19] cby_0__1__9_chany_bottom_out;
  wire [0:19] cby_0__1__9_chany_top_out;
  wire [0:0] cby_0__1__9_left_grid_pin_0_;
  wire [0:0] cby_12__1__0_ccff_tail;
  wire [0:19] cby_12__1__0_chany_bottom_out;
  wire [0:19] cby_12__1__0_chany_top_out;
  wire [0:0] cby_12__1__0_left_grid_pin_16_;
  wire [0:0] cby_12__1__0_left_grid_pin_17_;
  wire [0:0] cby_12__1__0_left_grid_pin_18_;
  wire [0:0] cby_12__1__0_left_grid_pin_19_;
  wire [0:0] cby_12__1__0_left_grid_pin_20_;
  wire [0:0] cby_12__1__0_left_grid_pin_21_;
  wire [0:0] cby_12__1__0_left_grid_pin_22_;
  wire [0:0] cby_12__1__0_left_grid_pin_23_;
  wire [0:0] cby_12__1__0_left_grid_pin_24_;
  wire [0:0] cby_12__1__0_left_grid_pin_25_;
  wire [0:0] cby_12__1__0_left_grid_pin_26_;
  wire [0:0] cby_12__1__0_left_grid_pin_27_;
  wire [0:0] cby_12__1__0_left_grid_pin_28_;
  wire [0:0] cby_12__1__0_left_grid_pin_29_;
  wire [0:0] cby_12__1__0_left_grid_pin_30_;
  wire [0:0] cby_12__1__0_left_grid_pin_31_;
  wire [0:0] cby_12__1__0_right_grid_pin_0_;
  wire [0:0] cby_12__1__10_ccff_tail;
  wire [0:19] cby_12__1__10_chany_bottom_out;
  wire [0:19] cby_12__1__10_chany_top_out;
  wire [0:0] cby_12__1__10_left_grid_pin_16_;
  wire [0:0] cby_12__1__10_left_grid_pin_17_;
  wire [0:0] cby_12__1__10_left_grid_pin_18_;
  wire [0:0] cby_12__1__10_left_grid_pin_19_;
  wire [0:0] cby_12__1__10_left_grid_pin_20_;
  wire [0:0] cby_12__1__10_left_grid_pin_21_;
  wire [0:0] cby_12__1__10_left_grid_pin_22_;
  wire [0:0] cby_12__1__10_left_grid_pin_23_;
  wire [0:0] cby_12__1__10_left_grid_pin_24_;
  wire [0:0] cby_12__1__10_left_grid_pin_25_;
  wire [0:0] cby_12__1__10_left_grid_pin_26_;
  wire [0:0] cby_12__1__10_left_grid_pin_27_;
  wire [0:0] cby_12__1__10_left_grid_pin_28_;
  wire [0:0] cby_12__1__10_left_grid_pin_29_;
  wire [0:0] cby_12__1__10_left_grid_pin_30_;
  wire [0:0] cby_12__1__10_left_grid_pin_31_;
  wire [0:0] cby_12__1__10_right_grid_pin_0_;
  wire [0:0] cby_12__1__11_ccff_tail;
  wire [0:19] cby_12__1__11_chany_bottom_out;
  wire [0:19] cby_12__1__11_chany_top_out;
  wire [0:0] cby_12__1__11_left_grid_pin_16_;
  wire [0:0] cby_12__1__11_left_grid_pin_17_;
  wire [0:0] cby_12__1__11_left_grid_pin_18_;
  wire [0:0] cby_12__1__11_left_grid_pin_19_;
  wire [0:0] cby_12__1__11_left_grid_pin_20_;
  wire [0:0] cby_12__1__11_left_grid_pin_21_;
  wire [0:0] cby_12__1__11_left_grid_pin_22_;
  wire [0:0] cby_12__1__11_left_grid_pin_23_;
  wire [0:0] cby_12__1__11_left_grid_pin_24_;
  wire [0:0] cby_12__1__11_left_grid_pin_25_;
  wire [0:0] cby_12__1__11_left_grid_pin_26_;
  wire [0:0] cby_12__1__11_left_grid_pin_27_;
  wire [0:0] cby_12__1__11_left_grid_pin_28_;
  wire [0:0] cby_12__1__11_left_grid_pin_29_;
  wire [0:0] cby_12__1__11_left_grid_pin_30_;
  wire [0:0] cby_12__1__11_left_grid_pin_31_;
  wire [0:0] cby_12__1__11_right_grid_pin_0_;
  wire [0:0] cby_12__1__1_ccff_tail;
  wire [0:19] cby_12__1__1_chany_bottom_out;
  wire [0:19] cby_12__1__1_chany_top_out;
  wire [0:0] cby_12__1__1_left_grid_pin_16_;
  wire [0:0] cby_12__1__1_left_grid_pin_17_;
  wire [0:0] cby_12__1__1_left_grid_pin_18_;
  wire [0:0] cby_12__1__1_left_grid_pin_19_;
  wire [0:0] cby_12__1__1_left_grid_pin_20_;
  wire [0:0] cby_12__1__1_left_grid_pin_21_;
  wire [0:0] cby_12__1__1_left_grid_pin_22_;
  wire [0:0] cby_12__1__1_left_grid_pin_23_;
  wire [0:0] cby_12__1__1_left_grid_pin_24_;
  wire [0:0] cby_12__1__1_left_grid_pin_25_;
  wire [0:0] cby_12__1__1_left_grid_pin_26_;
  wire [0:0] cby_12__1__1_left_grid_pin_27_;
  wire [0:0] cby_12__1__1_left_grid_pin_28_;
  wire [0:0] cby_12__1__1_left_grid_pin_29_;
  wire [0:0] cby_12__1__1_left_grid_pin_30_;
  wire [0:0] cby_12__1__1_left_grid_pin_31_;
  wire [0:0] cby_12__1__1_right_grid_pin_0_;
  wire [0:0] cby_12__1__2_ccff_tail;
  wire [0:19] cby_12__1__2_chany_bottom_out;
  wire [0:19] cby_12__1__2_chany_top_out;
  wire [0:0] cby_12__1__2_left_grid_pin_16_;
  wire [0:0] cby_12__1__2_left_grid_pin_17_;
  wire [0:0] cby_12__1__2_left_grid_pin_18_;
  wire [0:0] cby_12__1__2_left_grid_pin_19_;
  wire [0:0] cby_12__1__2_left_grid_pin_20_;
  wire [0:0] cby_12__1__2_left_grid_pin_21_;
  wire [0:0] cby_12__1__2_left_grid_pin_22_;
  wire [0:0] cby_12__1__2_left_grid_pin_23_;
  wire [0:0] cby_12__1__2_left_grid_pin_24_;
  wire [0:0] cby_12__1__2_left_grid_pin_25_;
  wire [0:0] cby_12__1__2_left_grid_pin_26_;
  wire [0:0] cby_12__1__2_left_grid_pin_27_;
  wire [0:0] cby_12__1__2_left_grid_pin_28_;
  wire [0:0] cby_12__1__2_left_grid_pin_29_;
  wire [0:0] cby_12__1__2_left_grid_pin_30_;
  wire [0:0] cby_12__1__2_left_grid_pin_31_;
  wire [0:0] cby_12__1__2_right_grid_pin_0_;
  wire [0:0] cby_12__1__3_ccff_tail;
  wire [0:19] cby_12__1__3_chany_bottom_out;
  wire [0:19] cby_12__1__3_chany_top_out;
  wire [0:0] cby_12__1__3_left_grid_pin_16_;
  wire [0:0] cby_12__1__3_left_grid_pin_17_;
  wire [0:0] cby_12__1__3_left_grid_pin_18_;
  wire [0:0] cby_12__1__3_left_grid_pin_19_;
  wire [0:0] cby_12__1__3_left_grid_pin_20_;
  wire [0:0] cby_12__1__3_left_grid_pin_21_;
  wire [0:0] cby_12__1__3_left_grid_pin_22_;
  wire [0:0] cby_12__1__3_left_grid_pin_23_;
  wire [0:0] cby_12__1__3_left_grid_pin_24_;
  wire [0:0] cby_12__1__3_left_grid_pin_25_;
  wire [0:0] cby_12__1__3_left_grid_pin_26_;
  wire [0:0] cby_12__1__3_left_grid_pin_27_;
  wire [0:0] cby_12__1__3_left_grid_pin_28_;
  wire [0:0] cby_12__1__3_left_grid_pin_29_;
  wire [0:0] cby_12__1__3_left_grid_pin_30_;
  wire [0:0] cby_12__1__3_left_grid_pin_31_;
  wire [0:0] cby_12__1__3_right_grid_pin_0_;
  wire [0:0] cby_12__1__4_ccff_tail;
  wire [0:19] cby_12__1__4_chany_bottom_out;
  wire [0:19] cby_12__1__4_chany_top_out;
  wire [0:0] cby_12__1__4_left_grid_pin_16_;
  wire [0:0] cby_12__1__4_left_grid_pin_17_;
  wire [0:0] cby_12__1__4_left_grid_pin_18_;
  wire [0:0] cby_12__1__4_left_grid_pin_19_;
  wire [0:0] cby_12__1__4_left_grid_pin_20_;
  wire [0:0] cby_12__1__4_left_grid_pin_21_;
  wire [0:0] cby_12__1__4_left_grid_pin_22_;
  wire [0:0] cby_12__1__4_left_grid_pin_23_;
  wire [0:0] cby_12__1__4_left_grid_pin_24_;
  wire [0:0] cby_12__1__4_left_grid_pin_25_;
  wire [0:0] cby_12__1__4_left_grid_pin_26_;
  wire [0:0] cby_12__1__4_left_grid_pin_27_;
  wire [0:0] cby_12__1__4_left_grid_pin_28_;
  wire [0:0] cby_12__1__4_left_grid_pin_29_;
  wire [0:0] cby_12__1__4_left_grid_pin_30_;
  wire [0:0] cby_12__1__4_left_grid_pin_31_;
  wire [0:0] cby_12__1__4_right_grid_pin_0_;
  wire [0:0] cby_12__1__5_ccff_tail;
  wire [0:19] cby_12__1__5_chany_bottom_out;
  wire [0:19] cby_12__1__5_chany_top_out;
  wire [0:0] cby_12__1__5_left_grid_pin_16_;
  wire [0:0] cby_12__1__5_left_grid_pin_17_;
  wire [0:0] cby_12__1__5_left_grid_pin_18_;
  wire [0:0] cby_12__1__5_left_grid_pin_19_;
  wire [0:0] cby_12__1__5_left_grid_pin_20_;
  wire [0:0] cby_12__1__5_left_grid_pin_21_;
  wire [0:0] cby_12__1__5_left_grid_pin_22_;
  wire [0:0] cby_12__1__5_left_grid_pin_23_;
  wire [0:0] cby_12__1__5_left_grid_pin_24_;
  wire [0:0] cby_12__1__5_left_grid_pin_25_;
  wire [0:0] cby_12__1__5_left_grid_pin_26_;
  wire [0:0] cby_12__1__5_left_grid_pin_27_;
  wire [0:0] cby_12__1__5_left_grid_pin_28_;
  wire [0:0] cby_12__1__5_left_grid_pin_29_;
  wire [0:0] cby_12__1__5_left_grid_pin_30_;
  wire [0:0] cby_12__1__5_left_grid_pin_31_;
  wire [0:0] cby_12__1__5_right_grid_pin_0_;
  wire [0:0] cby_12__1__6_ccff_tail;
  wire [0:19] cby_12__1__6_chany_bottom_out;
  wire [0:19] cby_12__1__6_chany_top_out;
  wire [0:0] cby_12__1__6_left_grid_pin_16_;
  wire [0:0] cby_12__1__6_left_grid_pin_17_;
  wire [0:0] cby_12__1__6_left_grid_pin_18_;
  wire [0:0] cby_12__1__6_left_grid_pin_19_;
  wire [0:0] cby_12__1__6_left_grid_pin_20_;
  wire [0:0] cby_12__1__6_left_grid_pin_21_;
  wire [0:0] cby_12__1__6_left_grid_pin_22_;
  wire [0:0] cby_12__1__6_left_grid_pin_23_;
  wire [0:0] cby_12__1__6_left_grid_pin_24_;
  wire [0:0] cby_12__1__6_left_grid_pin_25_;
  wire [0:0] cby_12__1__6_left_grid_pin_26_;
  wire [0:0] cby_12__1__6_left_grid_pin_27_;
  wire [0:0] cby_12__1__6_left_grid_pin_28_;
  wire [0:0] cby_12__1__6_left_grid_pin_29_;
  wire [0:0] cby_12__1__6_left_grid_pin_30_;
  wire [0:0] cby_12__1__6_left_grid_pin_31_;
  wire [0:0] cby_12__1__6_right_grid_pin_0_;
  wire [0:0] cby_12__1__7_ccff_tail;
  wire [0:19] cby_12__1__7_chany_bottom_out;
  wire [0:19] cby_12__1__7_chany_top_out;
  wire [0:0] cby_12__1__7_left_grid_pin_16_;
  wire [0:0] cby_12__1__7_left_grid_pin_17_;
  wire [0:0] cby_12__1__7_left_grid_pin_18_;
  wire [0:0] cby_12__1__7_left_grid_pin_19_;
  wire [0:0] cby_12__1__7_left_grid_pin_20_;
  wire [0:0] cby_12__1__7_left_grid_pin_21_;
  wire [0:0] cby_12__1__7_left_grid_pin_22_;
  wire [0:0] cby_12__1__7_left_grid_pin_23_;
  wire [0:0] cby_12__1__7_left_grid_pin_24_;
  wire [0:0] cby_12__1__7_left_grid_pin_25_;
  wire [0:0] cby_12__1__7_left_grid_pin_26_;
  wire [0:0] cby_12__1__7_left_grid_pin_27_;
  wire [0:0] cby_12__1__7_left_grid_pin_28_;
  wire [0:0] cby_12__1__7_left_grid_pin_29_;
  wire [0:0] cby_12__1__7_left_grid_pin_30_;
  wire [0:0] cby_12__1__7_left_grid_pin_31_;
  wire [0:0] cby_12__1__7_right_grid_pin_0_;
  wire [0:0] cby_12__1__8_ccff_tail;
  wire [0:19] cby_12__1__8_chany_bottom_out;
  wire [0:19] cby_12__1__8_chany_top_out;
  wire [0:0] cby_12__1__8_left_grid_pin_16_;
  wire [0:0] cby_12__1__8_left_grid_pin_17_;
  wire [0:0] cby_12__1__8_left_grid_pin_18_;
  wire [0:0] cby_12__1__8_left_grid_pin_19_;
  wire [0:0] cby_12__1__8_left_grid_pin_20_;
  wire [0:0] cby_12__1__8_left_grid_pin_21_;
  wire [0:0] cby_12__1__8_left_grid_pin_22_;
  wire [0:0] cby_12__1__8_left_grid_pin_23_;
  wire [0:0] cby_12__1__8_left_grid_pin_24_;
  wire [0:0] cby_12__1__8_left_grid_pin_25_;
  wire [0:0] cby_12__1__8_left_grid_pin_26_;
  wire [0:0] cby_12__1__8_left_grid_pin_27_;
  wire [0:0] cby_12__1__8_left_grid_pin_28_;
  wire [0:0] cby_12__1__8_left_grid_pin_29_;
  wire [0:0] cby_12__1__8_left_grid_pin_30_;
  wire [0:0] cby_12__1__8_left_grid_pin_31_;
  wire [0:0] cby_12__1__8_right_grid_pin_0_;
  wire [0:0] cby_12__1__9_ccff_tail;
  wire [0:19] cby_12__1__9_chany_bottom_out;
  wire [0:19] cby_12__1__9_chany_top_out;
  wire [0:0] cby_12__1__9_left_grid_pin_16_;
  wire [0:0] cby_12__1__9_left_grid_pin_17_;
  wire [0:0] cby_12__1__9_left_grid_pin_18_;
  wire [0:0] cby_12__1__9_left_grid_pin_19_;
  wire [0:0] cby_12__1__9_left_grid_pin_20_;
  wire [0:0] cby_12__1__9_left_grid_pin_21_;
  wire [0:0] cby_12__1__9_left_grid_pin_22_;
  wire [0:0] cby_12__1__9_left_grid_pin_23_;
  wire [0:0] cby_12__1__9_left_grid_pin_24_;
  wire [0:0] cby_12__1__9_left_grid_pin_25_;
  wire [0:0] cby_12__1__9_left_grid_pin_26_;
  wire [0:0] cby_12__1__9_left_grid_pin_27_;
  wire [0:0] cby_12__1__9_left_grid_pin_28_;
  wire [0:0] cby_12__1__9_left_grid_pin_29_;
  wire [0:0] cby_12__1__9_left_grid_pin_30_;
  wire [0:0] cby_12__1__9_left_grid_pin_31_;
  wire [0:0] cby_12__1__9_right_grid_pin_0_;
  wire [0:0] cby_1__1__0_ccff_tail;
  wire [0:19] cby_1__1__0_chany_bottom_out;
  wire [0:19] cby_1__1__0_chany_top_out;
  wire [0:0] cby_1__1__0_left_grid_pin_16_;
  wire [0:0] cby_1__1__0_left_grid_pin_17_;
  wire [0:0] cby_1__1__0_left_grid_pin_18_;
  wire [0:0] cby_1__1__0_left_grid_pin_19_;
  wire [0:0] cby_1__1__0_left_grid_pin_20_;
  wire [0:0] cby_1__1__0_left_grid_pin_21_;
  wire [0:0] cby_1__1__0_left_grid_pin_22_;
  wire [0:0] cby_1__1__0_left_grid_pin_23_;
  wire [0:0] cby_1__1__0_left_grid_pin_24_;
  wire [0:0] cby_1__1__0_left_grid_pin_25_;
  wire [0:0] cby_1__1__0_left_grid_pin_26_;
  wire [0:0] cby_1__1__0_left_grid_pin_27_;
  wire [0:0] cby_1__1__0_left_grid_pin_28_;
  wire [0:0] cby_1__1__0_left_grid_pin_29_;
  wire [0:0] cby_1__1__0_left_grid_pin_30_;
  wire [0:0] cby_1__1__0_left_grid_pin_31_;
  wire [0:0] cby_1__1__100_ccff_tail;
  wire [0:19] cby_1__1__100_chany_bottom_out;
  wire [0:19] cby_1__1__100_chany_top_out;
  wire [0:0] cby_1__1__100_left_grid_pin_16_;
  wire [0:0] cby_1__1__100_left_grid_pin_17_;
  wire [0:0] cby_1__1__100_left_grid_pin_18_;
  wire [0:0] cby_1__1__100_left_grid_pin_19_;
  wire [0:0] cby_1__1__100_left_grid_pin_20_;
  wire [0:0] cby_1__1__100_left_grid_pin_21_;
  wire [0:0] cby_1__1__100_left_grid_pin_22_;
  wire [0:0] cby_1__1__100_left_grid_pin_23_;
  wire [0:0] cby_1__1__100_left_grid_pin_24_;
  wire [0:0] cby_1__1__100_left_grid_pin_25_;
  wire [0:0] cby_1__1__100_left_grid_pin_26_;
  wire [0:0] cby_1__1__100_left_grid_pin_27_;
  wire [0:0] cby_1__1__100_left_grid_pin_28_;
  wire [0:0] cby_1__1__100_left_grid_pin_29_;
  wire [0:0] cby_1__1__100_left_grid_pin_30_;
  wire [0:0] cby_1__1__100_left_grid_pin_31_;
  wire [0:0] cby_1__1__101_ccff_tail;
  wire [0:19] cby_1__1__101_chany_bottom_out;
  wire [0:19] cby_1__1__101_chany_top_out;
  wire [0:0] cby_1__1__101_left_grid_pin_16_;
  wire [0:0] cby_1__1__101_left_grid_pin_17_;
  wire [0:0] cby_1__1__101_left_grid_pin_18_;
  wire [0:0] cby_1__1__101_left_grid_pin_19_;
  wire [0:0] cby_1__1__101_left_grid_pin_20_;
  wire [0:0] cby_1__1__101_left_grid_pin_21_;
  wire [0:0] cby_1__1__101_left_grid_pin_22_;
  wire [0:0] cby_1__1__101_left_grid_pin_23_;
  wire [0:0] cby_1__1__101_left_grid_pin_24_;
  wire [0:0] cby_1__1__101_left_grid_pin_25_;
  wire [0:0] cby_1__1__101_left_grid_pin_26_;
  wire [0:0] cby_1__1__101_left_grid_pin_27_;
  wire [0:0] cby_1__1__101_left_grid_pin_28_;
  wire [0:0] cby_1__1__101_left_grid_pin_29_;
  wire [0:0] cby_1__1__101_left_grid_pin_30_;
  wire [0:0] cby_1__1__101_left_grid_pin_31_;
  wire [0:0] cby_1__1__102_ccff_tail;
  wire [0:19] cby_1__1__102_chany_bottom_out;
  wire [0:19] cby_1__1__102_chany_top_out;
  wire [0:0] cby_1__1__102_left_grid_pin_16_;
  wire [0:0] cby_1__1__102_left_grid_pin_17_;
  wire [0:0] cby_1__1__102_left_grid_pin_18_;
  wire [0:0] cby_1__1__102_left_grid_pin_19_;
  wire [0:0] cby_1__1__102_left_grid_pin_20_;
  wire [0:0] cby_1__1__102_left_grid_pin_21_;
  wire [0:0] cby_1__1__102_left_grid_pin_22_;
  wire [0:0] cby_1__1__102_left_grid_pin_23_;
  wire [0:0] cby_1__1__102_left_grid_pin_24_;
  wire [0:0] cby_1__1__102_left_grid_pin_25_;
  wire [0:0] cby_1__1__102_left_grid_pin_26_;
  wire [0:0] cby_1__1__102_left_grid_pin_27_;
  wire [0:0] cby_1__1__102_left_grid_pin_28_;
  wire [0:0] cby_1__1__102_left_grid_pin_29_;
  wire [0:0] cby_1__1__102_left_grid_pin_30_;
  wire [0:0] cby_1__1__102_left_grid_pin_31_;
  wire [0:0] cby_1__1__103_ccff_tail;
  wire [0:19] cby_1__1__103_chany_bottom_out;
  wire [0:19] cby_1__1__103_chany_top_out;
  wire [0:0] cby_1__1__103_left_grid_pin_16_;
  wire [0:0] cby_1__1__103_left_grid_pin_17_;
  wire [0:0] cby_1__1__103_left_grid_pin_18_;
  wire [0:0] cby_1__1__103_left_grid_pin_19_;
  wire [0:0] cby_1__1__103_left_grid_pin_20_;
  wire [0:0] cby_1__1__103_left_grid_pin_21_;
  wire [0:0] cby_1__1__103_left_grid_pin_22_;
  wire [0:0] cby_1__1__103_left_grid_pin_23_;
  wire [0:0] cby_1__1__103_left_grid_pin_24_;
  wire [0:0] cby_1__1__103_left_grid_pin_25_;
  wire [0:0] cby_1__1__103_left_grid_pin_26_;
  wire [0:0] cby_1__1__103_left_grid_pin_27_;
  wire [0:0] cby_1__1__103_left_grid_pin_28_;
  wire [0:0] cby_1__1__103_left_grid_pin_29_;
  wire [0:0] cby_1__1__103_left_grid_pin_30_;
  wire [0:0] cby_1__1__103_left_grid_pin_31_;
  wire [0:0] cby_1__1__104_ccff_tail;
  wire [0:19] cby_1__1__104_chany_bottom_out;
  wire [0:19] cby_1__1__104_chany_top_out;
  wire [0:0] cby_1__1__104_left_grid_pin_16_;
  wire [0:0] cby_1__1__104_left_grid_pin_17_;
  wire [0:0] cby_1__1__104_left_grid_pin_18_;
  wire [0:0] cby_1__1__104_left_grid_pin_19_;
  wire [0:0] cby_1__1__104_left_grid_pin_20_;
  wire [0:0] cby_1__1__104_left_grid_pin_21_;
  wire [0:0] cby_1__1__104_left_grid_pin_22_;
  wire [0:0] cby_1__1__104_left_grid_pin_23_;
  wire [0:0] cby_1__1__104_left_grid_pin_24_;
  wire [0:0] cby_1__1__104_left_grid_pin_25_;
  wire [0:0] cby_1__1__104_left_grid_pin_26_;
  wire [0:0] cby_1__1__104_left_grid_pin_27_;
  wire [0:0] cby_1__1__104_left_grid_pin_28_;
  wire [0:0] cby_1__1__104_left_grid_pin_29_;
  wire [0:0] cby_1__1__104_left_grid_pin_30_;
  wire [0:0] cby_1__1__104_left_grid_pin_31_;
  wire [0:0] cby_1__1__105_ccff_tail;
  wire [0:19] cby_1__1__105_chany_bottom_out;
  wire [0:19] cby_1__1__105_chany_top_out;
  wire [0:0] cby_1__1__105_left_grid_pin_16_;
  wire [0:0] cby_1__1__105_left_grid_pin_17_;
  wire [0:0] cby_1__1__105_left_grid_pin_18_;
  wire [0:0] cby_1__1__105_left_grid_pin_19_;
  wire [0:0] cby_1__1__105_left_grid_pin_20_;
  wire [0:0] cby_1__1__105_left_grid_pin_21_;
  wire [0:0] cby_1__1__105_left_grid_pin_22_;
  wire [0:0] cby_1__1__105_left_grid_pin_23_;
  wire [0:0] cby_1__1__105_left_grid_pin_24_;
  wire [0:0] cby_1__1__105_left_grid_pin_25_;
  wire [0:0] cby_1__1__105_left_grid_pin_26_;
  wire [0:0] cby_1__1__105_left_grid_pin_27_;
  wire [0:0] cby_1__1__105_left_grid_pin_28_;
  wire [0:0] cby_1__1__105_left_grid_pin_29_;
  wire [0:0] cby_1__1__105_left_grid_pin_30_;
  wire [0:0] cby_1__1__105_left_grid_pin_31_;
  wire [0:0] cby_1__1__106_ccff_tail;
  wire [0:19] cby_1__1__106_chany_bottom_out;
  wire [0:19] cby_1__1__106_chany_top_out;
  wire [0:0] cby_1__1__106_left_grid_pin_16_;
  wire [0:0] cby_1__1__106_left_grid_pin_17_;
  wire [0:0] cby_1__1__106_left_grid_pin_18_;
  wire [0:0] cby_1__1__106_left_grid_pin_19_;
  wire [0:0] cby_1__1__106_left_grid_pin_20_;
  wire [0:0] cby_1__1__106_left_grid_pin_21_;
  wire [0:0] cby_1__1__106_left_grid_pin_22_;
  wire [0:0] cby_1__1__106_left_grid_pin_23_;
  wire [0:0] cby_1__1__106_left_grid_pin_24_;
  wire [0:0] cby_1__1__106_left_grid_pin_25_;
  wire [0:0] cby_1__1__106_left_grid_pin_26_;
  wire [0:0] cby_1__1__106_left_grid_pin_27_;
  wire [0:0] cby_1__1__106_left_grid_pin_28_;
  wire [0:0] cby_1__1__106_left_grid_pin_29_;
  wire [0:0] cby_1__1__106_left_grid_pin_30_;
  wire [0:0] cby_1__1__106_left_grid_pin_31_;
  wire [0:0] cby_1__1__107_ccff_tail;
  wire [0:19] cby_1__1__107_chany_bottom_out;
  wire [0:19] cby_1__1__107_chany_top_out;
  wire [0:0] cby_1__1__107_left_grid_pin_16_;
  wire [0:0] cby_1__1__107_left_grid_pin_17_;
  wire [0:0] cby_1__1__107_left_grid_pin_18_;
  wire [0:0] cby_1__1__107_left_grid_pin_19_;
  wire [0:0] cby_1__1__107_left_grid_pin_20_;
  wire [0:0] cby_1__1__107_left_grid_pin_21_;
  wire [0:0] cby_1__1__107_left_grid_pin_22_;
  wire [0:0] cby_1__1__107_left_grid_pin_23_;
  wire [0:0] cby_1__1__107_left_grid_pin_24_;
  wire [0:0] cby_1__1__107_left_grid_pin_25_;
  wire [0:0] cby_1__1__107_left_grid_pin_26_;
  wire [0:0] cby_1__1__107_left_grid_pin_27_;
  wire [0:0] cby_1__1__107_left_grid_pin_28_;
  wire [0:0] cby_1__1__107_left_grid_pin_29_;
  wire [0:0] cby_1__1__107_left_grid_pin_30_;
  wire [0:0] cby_1__1__107_left_grid_pin_31_;
  wire [0:0] cby_1__1__108_ccff_tail;
  wire [0:19] cby_1__1__108_chany_bottom_out;
  wire [0:19] cby_1__1__108_chany_top_out;
  wire [0:0] cby_1__1__108_left_grid_pin_16_;
  wire [0:0] cby_1__1__108_left_grid_pin_17_;
  wire [0:0] cby_1__1__108_left_grid_pin_18_;
  wire [0:0] cby_1__1__108_left_grid_pin_19_;
  wire [0:0] cby_1__1__108_left_grid_pin_20_;
  wire [0:0] cby_1__1__108_left_grid_pin_21_;
  wire [0:0] cby_1__1__108_left_grid_pin_22_;
  wire [0:0] cby_1__1__108_left_grid_pin_23_;
  wire [0:0] cby_1__1__108_left_grid_pin_24_;
  wire [0:0] cby_1__1__108_left_grid_pin_25_;
  wire [0:0] cby_1__1__108_left_grid_pin_26_;
  wire [0:0] cby_1__1__108_left_grid_pin_27_;
  wire [0:0] cby_1__1__108_left_grid_pin_28_;
  wire [0:0] cby_1__1__108_left_grid_pin_29_;
  wire [0:0] cby_1__1__108_left_grid_pin_30_;
  wire [0:0] cby_1__1__108_left_grid_pin_31_;
  wire [0:0] cby_1__1__109_ccff_tail;
  wire [0:19] cby_1__1__109_chany_bottom_out;
  wire [0:19] cby_1__1__109_chany_top_out;
  wire [0:0] cby_1__1__109_left_grid_pin_16_;
  wire [0:0] cby_1__1__109_left_grid_pin_17_;
  wire [0:0] cby_1__1__109_left_grid_pin_18_;
  wire [0:0] cby_1__1__109_left_grid_pin_19_;
  wire [0:0] cby_1__1__109_left_grid_pin_20_;
  wire [0:0] cby_1__1__109_left_grid_pin_21_;
  wire [0:0] cby_1__1__109_left_grid_pin_22_;
  wire [0:0] cby_1__1__109_left_grid_pin_23_;
  wire [0:0] cby_1__1__109_left_grid_pin_24_;
  wire [0:0] cby_1__1__109_left_grid_pin_25_;
  wire [0:0] cby_1__1__109_left_grid_pin_26_;
  wire [0:0] cby_1__1__109_left_grid_pin_27_;
  wire [0:0] cby_1__1__109_left_grid_pin_28_;
  wire [0:0] cby_1__1__109_left_grid_pin_29_;
  wire [0:0] cby_1__1__109_left_grid_pin_30_;
  wire [0:0] cby_1__1__109_left_grid_pin_31_;
  wire [0:0] cby_1__1__10_ccff_tail;
  wire [0:19] cby_1__1__10_chany_bottom_out;
  wire [0:19] cby_1__1__10_chany_top_out;
  wire [0:0] cby_1__1__10_left_grid_pin_16_;
  wire [0:0] cby_1__1__10_left_grid_pin_17_;
  wire [0:0] cby_1__1__10_left_grid_pin_18_;
  wire [0:0] cby_1__1__10_left_grid_pin_19_;
  wire [0:0] cby_1__1__10_left_grid_pin_20_;
  wire [0:0] cby_1__1__10_left_grid_pin_21_;
  wire [0:0] cby_1__1__10_left_grid_pin_22_;
  wire [0:0] cby_1__1__10_left_grid_pin_23_;
  wire [0:0] cby_1__1__10_left_grid_pin_24_;
  wire [0:0] cby_1__1__10_left_grid_pin_25_;
  wire [0:0] cby_1__1__10_left_grid_pin_26_;
  wire [0:0] cby_1__1__10_left_grid_pin_27_;
  wire [0:0] cby_1__1__10_left_grid_pin_28_;
  wire [0:0] cby_1__1__10_left_grid_pin_29_;
  wire [0:0] cby_1__1__10_left_grid_pin_30_;
  wire [0:0] cby_1__1__10_left_grid_pin_31_;
  wire [0:0] cby_1__1__110_ccff_tail;
  wire [0:19] cby_1__1__110_chany_bottom_out;
  wire [0:19] cby_1__1__110_chany_top_out;
  wire [0:0] cby_1__1__110_left_grid_pin_16_;
  wire [0:0] cby_1__1__110_left_grid_pin_17_;
  wire [0:0] cby_1__1__110_left_grid_pin_18_;
  wire [0:0] cby_1__1__110_left_grid_pin_19_;
  wire [0:0] cby_1__1__110_left_grid_pin_20_;
  wire [0:0] cby_1__1__110_left_grid_pin_21_;
  wire [0:0] cby_1__1__110_left_grid_pin_22_;
  wire [0:0] cby_1__1__110_left_grid_pin_23_;
  wire [0:0] cby_1__1__110_left_grid_pin_24_;
  wire [0:0] cby_1__1__110_left_grid_pin_25_;
  wire [0:0] cby_1__1__110_left_grid_pin_26_;
  wire [0:0] cby_1__1__110_left_grid_pin_27_;
  wire [0:0] cby_1__1__110_left_grid_pin_28_;
  wire [0:0] cby_1__1__110_left_grid_pin_29_;
  wire [0:0] cby_1__1__110_left_grid_pin_30_;
  wire [0:0] cby_1__1__110_left_grid_pin_31_;
  wire [0:0] cby_1__1__111_ccff_tail;
  wire [0:19] cby_1__1__111_chany_bottom_out;
  wire [0:19] cby_1__1__111_chany_top_out;
  wire [0:0] cby_1__1__111_left_grid_pin_16_;
  wire [0:0] cby_1__1__111_left_grid_pin_17_;
  wire [0:0] cby_1__1__111_left_grid_pin_18_;
  wire [0:0] cby_1__1__111_left_grid_pin_19_;
  wire [0:0] cby_1__1__111_left_grid_pin_20_;
  wire [0:0] cby_1__1__111_left_grid_pin_21_;
  wire [0:0] cby_1__1__111_left_grid_pin_22_;
  wire [0:0] cby_1__1__111_left_grid_pin_23_;
  wire [0:0] cby_1__1__111_left_grid_pin_24_;
  wire [0:0] cby_1__1__111_left_grid_pin_25_;
  wire [0:0] cby_1__1__111_left_grid_pin_26_;
  wire [0:0] cby_1__1__111_left_grid_pin_27_;
  wire [0:0] cby_1__1__111_left_grid_pin_28_;
  wire [0:0] cby_1__1__111_left_grid_pin_29_;
  wire [0:0] cby_1__1__111_left_grid_pin_30_;
  wire [0:0] cby_1__1__111_left_grid_pin_31_;
  wire [0:0] cby_1__1__112_ccff_tail;
  wire [0:19] cby_1__1__112_chany_bottom_out;
  wire [0:19] cby_1__1__112_chany_top_out;
  wire [0:0] cby_1__1__112_left_grid_pin_16_;
  wire [0:0] cby_1__1__112_left_grid_pin_17_;
  wire [0:0] cby_1__1__112_left_grid_pin_18_;
  wire [0:0] cby_1__1__112_left_grid_pin_19_;
  wire [0:0] cby_1__1__112_left_grid_pin_20_;
  wire [0:0] cby_1__1__112_left_grid_pin_21_;
  wire [0:0] cby_1__1__112_left_grid_pin_22_;
  wire [0:0] cby_1__1__112_left_grid_pin_23_;
  wire [0:0] cby_1__1__112_left_grid_pin_24_;
  wire [0:0] cby_1__1__112_left_grid_pin_25_;
  wire [0:0] cby_1__1__112_left_grid_pin_26_;
  wire [0:0] cby_1__1__112_left_grid_pin_27_;
  wire [0:0] cby_1__1__112_left_grid_pin_28_;
  wire [0:0] cby_1__1__112_left_grid_pin_29_;
  wire [0:0] cby_1__1__112_left_grid_pin_30_;
  wire [0:0] cby_1__1__112_left_grid_pin_31_;
  wire [0:0] cby_1__1__113_ccff_tail;
  wire [0:19] cby_1__1__113_chany_bottom_out;
  wire [0:19] cby_1__1__113_chany_top_out;
  wire [0:0] cby_1__1__113_left_grid_pin_16_;
  wire [0:0] cby_1__1__113_left_grid_pin_17_;
  wire [0:0] cby_1__1__113_left_grid_pin_18_;
  wire [0:0] cby_1__1__113_left_grid_pin_19_;
  wire [0:0] cby_1__1__113_left_grid_pin_20_;
  wire [0:0] cby_1__1__113_left_grid_pin_21_;
  wire [0:0] cby_1__1__113_left_grid_pin_22_;
  wire [0:0] cby_1__1__113_left_grid_pin_23_;
  wire [0:0] cby_1__1__113_left_grid_pin_24_;
  wire [0:0] cby_1__1__113_left_grid_pin_25_;
  wire [0:0] cby_1__1__113_left_grid_pin_26_;
  wire [0:0] cby_1__1__113_left_grid_pin_27_;
  wire [0:0] cby_1__1__113_left_grid_pin_28_;
  wire [0:0] cby_1__1__113_left_grid_pin_29_;
  wire [0:0] cby_1__1__113_left_grid_pin_30_;
  wire [0:0] cby_1__1__113_left_grid_pin_31_;
  wire [0:0] cby_1__1__114_ccff_tail;
  wire [0:19] cby_1__1__114_chany_bottom_out;
  wire [0:19] cby_1__1__114_chany_top_out;
  wire [0:0] cby_1__1__114_left_grid_pin_16_;
  wire [0:0] cby_1__1__114_left_grid_pin_17_;
  wire [0:0] cby_1__1__114_left_grid_pin_18_;
  wire [0:0] cby_1__1__114_left_grid_pin_19_;
  wire [0:0] cby_1__1__114_left_grid_pin_20_;
  wire [0:0] cby_1__1__114_left_grid_pin_21_;
  wire [0:0] cby_1__1__114_left_grid_pin_22_;
  wire [0:0] cby_1__1__114_left_grid_pin_23_;
  wire [0:0] cby_1__1__114_left_grid_pin_24_;
  wire [0:0] cby_1__1__114_left_grid_pin_25_;
  wire [0:0] cby_1__1__114_left_grid_pin_26_;
  wire [0:0] cby_1__1__114_left_grid_pin_27_;
  wire [0:0] cby_1__1__114_left_grid_pin_28_;
  wire [0:0] cby_1__1__114_left_grid_pin_29_;
  wire [0:0] cby_1__1__114_left_grid_pin_30_;
  wire [0:0] cby_1__1__114_left_grid_pin_31_;
  wire [0:0] cby_1__1__115_ccff_tail;
  wire [0:19] cby_1__1__115_chany_bottom_out;
  wire [0:19] cby_1__1__115_chany_top_out;
  wire [0:0] cby_1__1__115_left_grid_pin_16_;
  wire [0:0] cby_1__1__115_left_grid_pin_17_;
  wire [0:0] cby_1__1__115_left_grid_pin_18_;
  wire [0:0] cby_1__1__115_left_grid_pin_19_;
  wire [0:0] cby_1__1__115_left_grid_pin_20_;
  wire [0:0] cby_1__1__115_left_grid_pin_21_;
  wire [0:0] cby_1__1__115_left_grid_pin_22_;
  wire [0:0] cby_1__1__115_left_grid_pin_23_;
  wire [0:0] cby_1__1__115_left_grid_pin_24_;
  wire [0:0] cby_1__1__115_left_grid_pin_25_;
  wire [0:0] cby_1__1__115_left_grid_pin_26_;
  wire [0:0] cby_1__1__115_left_grid_pin_27_;
  wire [0:0] cby_1__1__115_left_grid_pin_28_;
  wire [0:0] cby_1__1__115_left_grid_pin_29_;
  wire [0:0] cby_1__1__115_left_grid_pin_30_;
  wire [0:0] cby_1__1__115_left_grid_pin_31_;
  wire [0:0] cby_1__1__116_ccff_tail;
  wire [0:19] cby_1__1__116_chany_bottom_out;
  wire [0:19] cby_1__1__116_chany_top_out;
  wire [0:0] cby_1__1__116_left_grid_pin_16_;
  wire [0:0] cby_1__1__116_left_grid_pin_17_;
  wire [0:0] cby_1__1__116_left_grid_pin_18_;
  wire [0:0] cby_1__1__116_left_grid_pin_19_;
  wire [0:0] cby_1__1__116_left_grid_pin_20_;
  wire [0:0] cby_1__1__116_left_grid_pin_21_;
  wire [0:0] cby_1__1__116_left_grid_pin_22_;
  wire [0:0] cby_1__1__116_left_grid_pin_23_;
  wire [0:0] cby_1__1__116_left_grid_pin_24_;
  wire [0:0] cby_1__1__116_left_grid_pin_25_;
  wire [0:0] cby_1__1__116_left_grid_pin_26_;
  wire [0:0] cby_1__1__116_left_grid_pin_27_;
  wire [0:0] cby_1__1__116_left_grid_pin_28_;
  wire [0:0] cby_1__1__116_left_grid_pin_29_;
  wire [0:0] cby_1__1__116_left_grid_pin_30_;
  wire [0:0] cby_1__1__116_left_grid_pin_31_;
  wire [0:0] cby_1__1__117_ccff_tail;
  wire [0:19] cby_1__1__117_chany_bottom_out;
  wire [0:19] cby_1__1__117_chany_top_out;
  wire [0:0] cby_1__1__117_left_grid_pin_16_;
  wire [0:0] cby_1__1__117_left_grid_pin_17_;
  wire [0:0] cby_1__1__117_left_grid_pin_18_;
  wire [0:0] cby_1__1__117_left_grid_pin_19_;
  wire [0:0] cby_1__1__117_left_grid_pin_20_;
  wire [0:0] cby_1__1__117_left_grid_pin_21_;
  wire [0:0] cby_1__1__117_left_grid_pin_22_;
  wire [0:0] cby_1__1__117_left_grid_pin_23_;
  wire [0:0] cby_1__1__117_left_grid_pin_24_;
  wire [0:0] cby_1__1__117_left_grid_pin_25_;
  wire [0:0] cby_1__1__117_left_grid_pin_26_;
  wire [0:0] cby_1__1__117_left_grid_pin_27_;
  wire [0:0] cby_1__1__117_left_grid_pin_28_;
  wire [0:0] cby_1__1__117_left_grid_pin_29_;
  wire [0:0] cby_1__1__117_left_grid_pin_30_;
  wire [0:0] cby_1__1__117_left_grid_pin_31_;
  wire [0:0] cby_1__1__118_ccff_tail;
  wire [0:19] cby_1__1__118_chany_bottom_out;
  wire [0:19] cby_1__1__118_chany_top_out;
  wire [0:0] cby_1__1__118_left_grid_pin_16_;
  wire [0:0] cby_1__1__118_left_grid_pin_17_;
  wire [0:0] cby_1__1__118_left_grid_pin_18_;
  wire [0:0] cby_1__1__118_left_grid_pin_19_;
  wire [0:0] cby_1__1__118_left_grid_pin_20_;
  wire [0:0] cby_1__1__118_left_grid_pin_21_;
  wire [0:0] cby_1__1__118_left_grid_pin_22_;
  wire [0:0] cby_1__1__118_left_grid_pin_23_;
  wire [0:0] cby_1__1__118_left_grid_pin_24_;
  wire [0:0] cby_1__1__118_left_grid_pin_25_;
  wire [0:0] cby_1__1__118_left_grid_pin_26_;
  wire [0:0] cby_1__1__118_left_grid_pin_27_;
  wire [0:0] cby_1__1__118_left_grid_pin_28_;
  wire [0:0] cby_1__1__118_left_grid_pin_29_;
  wire [0:0] cby_1__1__118_left_grid_pin_30_;
  wire [0:0] cby_1__1__118_left_grid_pin_31_;
  wire [0:0] cby_1__1__119_ccff_tail;
  wire [0:19] cby_1__1__119_chany_bottom_out;
  wire [0:19] cby_1__1__119_chany_top_out;
  wire [0:0] cby_1__1__119_left_grid_pin_16_;
  wire [0:0] cby_1__1__119_left_grid_pin_17_;
  wire [0:0] cby_1__1__119_left_grid_pin_18_;
  wire [0:0] cby_1__1__119_left_grid_pin_19_;
  wire [0:0] cby_1__1__119_left_grid_pin_20_;
  wire [0:0] cby_1__1__119_left_grid_pin_21_;
  wire [0:0] cby_1__1__119_left_grid_pin_22_;
  wire [0:0] cby_1__1__119_left_grid_pin_23_;
  wire [0:0] cby_1__1__119_left_grid_pin_24_;
  wire [0:0] cby_1__1__119_left_grid_pin_25_;
  wire [0:0] cby_1__1__119_left_grid_pin_26_;
  wire [0:0] cby_1__1__119_left_grid_pin_27_;
  wire [0:0] cby_1__1__119_left_grid_pin_28_;
  wire [0:0] cby_1__1__119_left_grid_pin_29_;
  wire [0:0] cby_1__1__119_left_grid_pin_30_;
  wire [0:0] cby_1__1__119_left_grid_pin_31_;
  wire [0:0] cby_1__1__11_ccff_tail;
  wire [0:19] cby_1__1__11_chany_bottom_out;
  wire [0:19] cby_1__1__11_chany_top_out;
  wire [0:0] cby_1__1__11_left_grid_pin_16_;
  wire [0:0] cby_1__1__11_left_grid_pin_17_;
  wire [0:0] cby_1__1__11_left_grid_pin_18_;
  wire [0:0] cby_1__1__11_left_grid_pin_19_;
  wire [0:0] cby_1__1__11_left_grid_pin_20_;
  wire [0:0] cby_1__1__11_left_grid_pin_21_;
  wire [0:0] cby_1__1__11_left_grid_pin_22_;
  wire [0:0] cby_1__1__11_left_grid_pin_23_;
  wire [0:0] cby_1__1__11_left_grid_pin_24_;
  wire [0:0] cby_1__1__11_left_grid_pin_25_;
  wire [0:0] cby_1__1__11_left_grid_pin_26_;
  wire [0:0] cby_1__1__11_left_grid_pin_27_;
  wire [0:0] cby_1__1__11_left_grid_pin_28_;
  wire [0:0] cby_1__1__11_left_grid_pin_29_;
  wire [0:0] cby_1__1__11_left_grid_pin_30_;
  wire [0:0] cby_1__1__11_left_grid_pin_31_;
  wire [0:0] cby_1__1__120_ccff_tail;
  wire [0:19] cby_1__1__120_chany_bottom_out;
  wire [0:19] cby_1__1__120_chany_top_out;
  wire [0:0] cby_1__1__120_left_grid_pin_16_;
  wire [0:0] cby_1__1__120_left_grid_pin_17_;
  wire [0:0] cby_1__1__120_left_grid_pin_18_;
  wire [0:0] cby_1__1__120_left_grid_pin_19_;
  wire [0:0] cby_1__1__120_left_grid_pin_20_;
  wire [0:0] cby_1__1__120_left_grid_pin_21_;
  wire [0:0] cby_1__1__120_left_grid_pin_22_;
  wire [0:0] cby_1__1__120_left_grid_pin_23_;
  wire [0:0] cby_1__1__120_left_grid_pin_24_;
  wire [0:0] cby_1__1__120_left_grid_pin_25_;
  wire [0:0] cby_1__1__120_left_grid_pin_26_;
  wire [0:0] cby_1__1__120_left_grid_pin_27_;
  wire [0:0] cby_1__1__120_left_grid_pin_28_;
  wire [0:0] cby_1__1__120_left_grid_pin_29_;
  wire [0:0] cby_1__1__120_left_grid_pin_30_;
  wire [0:0] cby_1__1__120_left_grid_pin_31_;
  wire [0:0] cby_1__1__121_ccff_tail;
  wire [0:19] cby_1__1__121_chany_bottom_out;
  wire [0:19] cby_1__1__121_chany_top_out;
  wire [0:0] cby_1__1__121_left_grid_pin_16_;
  wire [0:0] cby_1__1__121_left_grid_pin_17_;
  wire [0:0] cby_1__1__121_left_grid_pin_18_;
  wire [0:0] cby_1__1__121_left_grid_pin_19_;
  wire [0:0] cby_1__1__121_left_grid_pin_20_;
  wire [0:0] cby_1__1__121_left_grid_pin_21_;
  wire [0:0] cby_1__1__121_left_grid_pin_22_;
  wire [0:0] cby_1__1__121_left_grid_pin_23_;
  wire [0:0] cby_1__1__121_left_grid_pin_24_;
  wire [0:0] cby_1__1__121_left_grid_pin_25_;
  wire [0:0] cby_1__1__121_left_grid_pin_26_;
  wire [0:0] cby_1__1__121_left_grid_pin_27_;
  wire [0:0] cby_1__1__121_left_grid_pin_28_;
  wire [0:0] cby_1__1__121_left_grid_pin_29_;
  wire [0:0] cby_1__1__121_left_grid_pin_30_;
  wire [0:0] cby_1__1__121_left_grid_pin_31_;
  wire [0:0] cby_1__1__122_ccff_tail;
  wire [0:19] cby_1__1__122_chany_bottom_out;
  wire [0:19] cby_1__1__122_chany_top_out;
  wire [0:0] cby_1__1__122_left_grid_pin_16_;
  wire [0:0] cby_1__1__122_left_grid_pin_17_;
  wire [0:0] cby_1__1__122_left_grid_pin_18_;
  wire [0:0] cby_1__1__122_left_grid_pin_19_;
  wire [0:0] cby_1__1__122_left_grid_pin_20_;
  wire [0:0] cby_1__1__122_left_grid_pin_21_;
  wire [0:0] cby_1__1__122_left_grid_pin_22_;
  wire [0:0] cby_1__1__122_left_grid_pin_23_;
  wire [0:0] cby_1__1__122_left_grid_pin_24_;
  wire [0:0] cby_1__1__122_left_grid_pin_25_;
  wire [0:0] cby_1__1__122_left_grid_pin_26_;
  wire [0:0] cby_1__1__122_left_grid_pin_27_;
  wire [0:0] cby_1__1__122_left_grid_pin_28_;
  wire [0:0] cby_1__1__122_left_grid_pin_29_;
  wire [0:0] cby_1__1__122_left_grid_pin_30_;
  wire [0:0] cby_1__1__122_left_grid_pin_31_;
  wire [0:0] cby_1__1__123_ccff_tail;
  wire [0:19] cby_1__1__123_chany_bottom_out;
  wire [0:19] cby_1__1__123_chany_top_out;
  wire [0:0] cby_1__1__123_left_grid_pin_16_;
  wire [0:0] cby_1__1__123_left_grid_pin_17_;
  wire [0:0] cby_1__1__123_left_grid_pin_18_;
  wire [0:0] cby_1__1__123_left_grid_pin_19_;
  wire [0:0] cby_1__1__123_left_grid_pin_20_;
  wire [0:0] cby_1__1__123_left_grid_pin_21_;
  wire [0:0] cby_1__1__123_left_grid_pin_22_;
  wire [0:0] cby_1__1__123_left_grid_pin_23_;
  wire [0:0] cby_1__1__123_left_grid_pin_24_;
  wire [0:0] cby_1__1__123_left_grid_pin_25_;
  wire [0:0] cby_1__1__123_left_grid_pin_26_;
  wire [0:0] cby_1__1__123_left_grid_pin_27_;
  wire [0:0] cby_1__1__123_left_grid_pin_28_;
  wire [0:0] cby_1__1__123_left_grid_pin_29_;
  wire [0:0] cby_1__1__123_left_grid_pin_30_;
  wire [0:0] cby_1__1__123_left_grid_pin_31_;
  wire [0:0] cby_1__1__124_ccff_tail;
  wire [0:19] cby_1__1__124_chany_bottom_out;
  wire [0:19] cby_1__1__124_chany_top_out;
  wire [0:0] cby_1__1__124_left_grid_pin_16_;
  wire [0:0] cby_1__1__124_left_grid_pin_17_;
  wire [0:0] cby_1__1__124_left_grid_pin_18_;
  wire [0:0] cby_1__1__124_left_grid_pin_19_;
  wire [0:0] cby_1__1__124_left_grid_pin_20_;
  wire [0:0] cby_1__1__124_left_grid_pin_21_;
  wire [0:0] cby_1__1__124_left_grid_pin_22_;
  wire [0:0] cby_1__1__124_left_grid_pin_23_;
  wire [0:0] cby_1__1__124_left_grid_pin_24_;
  wire [0:0] cby_1__1__124_left_grid_pin_25_;
  wire [0:0] cby_1__1__124_left_grid_pin_26_;
  wire [0:0] cby_1__1__124_left_grid_pin_27_;
  wire [0:0] cby_1__1__124_left_grid_pin_28_;
  wire [0:0] cby_1__1__124_left_grid_pin_29_;
  wire [0:0] cby_1__1__124_left_grid_pin_30_;
  wire [0:0] cby_1__1__124_left_grid_pin_31_;
  wire [0:0] cby_1__1__125_ccff_tail;
  wire [0:19] cby_1__1__125_chany_bottom_out;
  wire [0:19] cby_1__1__125_chany_top_out;
  wire [0:0] cby_1__1__125_left_grid_pin_16_;
  wire [0:0] cby_1__1__125_left_grid_pin_17_;
  wire [0:0] cby_1__1__125_left_grid_pin_18_;
  wire [0:0] cby_1__1__125_left_grid_pin_19_;
  wire [0:0] cby_1__1__125_left_grid_pin_20_;
  wire [0:0] cby_1__1__125_left_grid_pin_21_;
  wire [0:0] cby_1__1__125_left_grid_pin_22_;
  wire [0:0] cby_1__1__125_left_grid_pin_23_;
  wire [0:0] cby_1__1__125_left_grid_pin_24_;
  wire [0:0] cby_1__1__125_left_grid_pin_25_;
  wire [0:0] cby_1__1__125_left_grid_pin_26_;
  wire [0:0] cby_1__1__125_left_grid_pin_27_;
  wire [0:0] cby_1__1__125_left_grid_pin_28_;
  wire [0:0] cby_1__1__125_left_grid_pin_29_;
  wire [0:0] cby_1__1__125_left_grid_pin_30_;
  wire [0:0] cby_1__1__125_left_grid_pin_31_;
  wire [0:0] cby_1__1__126_ccff_tail;
  wire [0:19] cby_1__1__126_chany_bottom_out;
  wire [0:19] cby_1__1__126_chany_top_out;
  wire [0:0] cby_1__1__126_left_grid_pin_16_;
  wire [0:0] cby_1__1__126_left_grid_pin_17_;
  wire [0:0] cby_1__1__126_left_grid_pin_18_;
  wire [0:0] cby_1__1__126_left_grid_pin_19_;
  wire [0:0] cby_1__1__126_left_grid_pin_20_;
  wire [0:0] cby_1__1__126_left_grid_pin_21_;
  wire [0:0] cby_1__1__126_left_grid_pin_22_;
  wire [0:0] cby_1__1__126_left_grid_pin_23_;
  wire [0:0] cby_1__1__126_left_grid_pin_24_;
  wire [0:0] cby_1__1__126_left_grid_pin_25_;
  wire [0:0] cby_1__1__126_left_grid_pin_26_;
  wire [0:0] cby_1__1__126_left_grid_pin_27_;
  wire [0:0] cby_1__1__126_left_grid_pin_28_;
  wire [0:0] cby_1__1__126_left_grid_pin_29_;
  wire [0:0] cby_1__1__126_left_grid_pin_30_;
  wire [0:0] cby_1__1__126_left_grid_pin_31_;
  wire [0:0] cby_1__1__127_ccff_tail;
  wire [0:19] cby_1__1__127_chany_bottom_out;
  wire [0:19] cby_1__1__127_chany_top_out;
  wire [0:0] cby_1__1__127_left_grid_pin_16_;
  wire [0:0] cby_1__1__127_left_grid_pin_17_;
  wire [0:0] cby_1__1__127_left_grid_pin_18_;
  wire [0:0] cby_1__1__127_left_grid_pin_19_;
  wire [0:0] cby_1__1__127_left_grid_pin_20_;
  wire [0:0] cby_1__1__127_left_grid_pin_21_;
  wire [0:0] cby_1__1__127_left_grid_pin_22_;
  wire [0:0] cby_1__1__127_left_grid_pin_23_;
  wire [0:0] cby_1__1__127_left_grid_pin_24_;
  wire [0:0] cby_1__1__127_left_grid_pin_25_;
  wire [0:0] cby_1__1__127_left_grid_pin_26_;
  wire [0:0] cby_1__1__127_left_grid_pin_27_;
  wire [0:0] cby_1__1__127_left_grid_pin_28_;
  wire [0:0] cby_1__1__127_left_grid_pin_29_;
  wire [0:0] cby_1__1__127_left_grid_pin_30_;
  wire [0:0] cby_1__1__127_left_grid_pin_31_;
  wire [0:0] cby_1__1__128_ccff_tail;
  wire [0:19] cby_1__1__128_chany_bottom_out;
  wire [0:19] cby_1__1__128_chany_top_out;
  wire [0:0] cby_1__1__128_left_grid_pin_16_;
  wire [0:0] cby_1__1__128_left_grid_pin_17_;
  wire [0:0] cby_1__1__128_left_grid_pin_18_;
  wire [0:0] cby_1__1__128_left_grid_pin_19_;
  wire [0:0] cby_1__1__128_left_grid_pin_20_;
  wire [0:0] cby_1__1__128_left_grid_pin_21_;
  wire [0:0] cby_1__1__128_left_grid_pin_22_;
  wire [0:0] cby_1__1__128_left_grid_pin_23_;
  wire [0:0] cby_1__1__128_left_grid_pin_24_;
  wire [0:0] cby_1__1__128_left_grid_pin_25_;
  wire [0:0] cby_1__1__128_left_grid_pin_26_;
  wire [0:0] cby_1__1__128_left_grid_pin_27_;
  wire [0:0] cby_1__1__128_left_grid_pin_28_;
  wire [0:0] cby_1__1__128_left_grid_pin_29_;
  wire [0:0] cby_1__1__128_left_grid_pin_30_;
  wire [0:0] cby_1__1__128_left_grid_pin_31_;
  wire [0:0] cby_1__1__129_ccff_tail;
  wire [0:19] cby_1__1__129_chany_bottom_out;
  wire [0:19] cby_1__1__129_chany_top_out;
  wire [0:0] cby_1__1__129_left_grid_pin_16_;
  wire [0:0] cby_1__1__129_left_grid_pin_17_;
  wire [0:0] cby_1__1__129_left_grid_pin_18_;
  wire [0:0] cby_1__1__129_left_grid_pin_19_;
  wire [0:0] cby_1__1__129_left_grid_pin_20_;
  wire [0:0] cby_1__1__129_left_grid_pin_21_;
  wire [0:0] cby_1__1__129_left_grid_pin_22_;
  wire [0:0] cby_1__1__129_left_grid_pin_23_;
  wire [0:0] cby_1__1__129_left_grid_pin_24_;
  wire [0:0] cby_1__1__129_left_grid_pin_25_;
  wire [0:0] cby_1__1__129_left_grid_pin_26_;
  wire [0:0] cby_1__1__129_left_grid_pin_27_;
  wire [0:0] cby_1__1__129_left_grid_pin_28_;
  wire [0:0] cby_1__1__129_left_grid_pin_29_;
  wire [0:0] cby_1__1__129_left_grid_pin_30_;
  wire [0:0] cby_1__1__129_left_grid_pin_31_;
  wire [0:0] cby_1__1__12_ccff_tail;
  wire [0:19] cby_1__1__12_chany_bottom_out;
  wire [0:19] cby_1__1__12_chany_top_out;
  wire [0:0] cby_1__1__12_left_grid_pin_16_;
  wire [0:0] cby_1__1__12_left_grid_pin_17_;
  wire [0:0] cby_1__1__12_left_grid_pin_18_;
  wire [0:0] cby_1__1__12_left_grid_pin_19_;
  wire [0:0] cby_1__1__12_left_grid_pin_20_;
  wire [0:0] cby_1__1__12_left_grid_pin_21_;
  wire [0:0] cby_1__1__12_left_grid_pin_22_;
  wire [0:0] cby_1__1__12_left_grid_pin_23_;
  wire [0:0] cby_1__1__12_left_grid_pin_24_;
  wire [0:0] cby_1__1__12_left_grid_pin_25_;
  wire [0:0] cby_1__1__12_left_grid_pin_26_;
  wire [0:0] cby_1__1__12_left_grid_pin_27_;
  wire [0:0] cby_1__1__12_left_grid_pin_28_;
  wire [0:0] cby_1__1__12_left_grid_pin_29_;
  wire [0:0] cby_1__1__12_left_grid_pin_30_;
  wire [0:0] cby_1__1__12_left_grid_pin_31_;
  wire [0:0] cby_1__1__130_ccff_tail;
  wire [0:19] cby_1__1__130_chany_bottom_out;
  wire [0:19] cby_1__1__130_chany_top_out;
  wire [0:0] cby_1__1__130_left_grid_pin_16_;
  wire [0:0] cby_1__1__130_left_grid_pin_17_;
  wire [0:0] cby_1__1__130_left_grid_pin_18_;
  wire [0:0] cby_1__1__130_left_grid_pin_19_;
  wire [0:0] cby_1__1__130_left_grid_pin_20_;
  wire [0:0] cby_1__1__130_left_grid_pin_21_;
  wire [0:0] cby_1__1__130_left_grid_pin_22_;
  wire [0:0] cby_1__1__130_left_grid_pin_23_;
  wire [0:0] cby_1__1__130_left_grid_pin_24_;
  wire [0:0] cby_1__1__130_left_grid_pin_25_;
  wire [0:0] cby_1__1__130_left_grid_pin_26_;
  wire [0:0] cby_1__1__130_left_grid_pin_27_;
  wire [0:0] cby_1__1__130_left_grid_pin_28_;
  wire [0:0] cby_1__1__130_left_grid_pin_29_;
  wire [0:0] cby_1__1__130_left_grid_pin_30_;
  wire [0:0] cby_1__1__130_left_grid_pin_31_;
  wire [0:0] cby_1__1__131_ccff_tail;
  wire [0:19] cby_1__1__131_chany_bottom_out;
  wire [0:19] cby_1__1__131_chany_top_out;
  wire [0:0] cby_1__1__131_left_grid_pin_16_;
  wire [0:0] cby_1__1__131_left_grid_pin_17_;
  wire [0:0] cby_1__1__131_left_grid_pin_18_;
  wire [0:0] cby_1__1__131_left_grid_pin_19_;
  wire [0:0] cby_1__1__131_left_grid_pin_20_;
  wire [0:0] cby_1__1__131_left_grid_pin_21_;
  wire [0:0] cby_1__1__131_left_grid_pin_22_;
  wire [0:0] cby_1__1__131_left_grid_pin_23_;
  wire [0:0] cby_1__1__131_left_grid_pin_24_;
  wire [0:0] cby_1__1__131_left_grid_pin_25_;
  wire [0:0] cby_1__1__131_left_grid_pin_26_;
  wire [0:0] cby_1__1__131_left_grid_pin_27_;
  wire [0:0] cby_1__1__131_left_grid_pin_28_;
  wire [0:0] cby_1__1__131_left_grid_pin_29_;
  wire [0:0] cby_1__1__131_left_grid_pin_30_;
  wire [0:0] cby_1__1__131_left_grid_pin_31_;
  wire [0:0] cby_1__1__13_ccff_tail;
  wire [0:19] cby_1__1__13_chany_bottom_out;
  wire [0:19] cby_1__1__13_chany_top_out;
  wire [0:0] cby_1__1__13_left_grid_pin_16_;
  wire [0:0] cby_1__1__13_left_grid_pin_17_;
  wire [0:0] cby_1__1__13_left_grid_pin_18_;
  wire [0:0] cby_1__1__13_left_grid_pin_19_;
  wire [0:0] cby_1__1__13_left_grid_pin_20_;
  wire [0:0] cby_1__1__13_left_grid_pin_21_;
  wire [0:0] cby_1__1__13_left_grid_pin_22_;
  wire [0:0] cby_1__1__13_left_grid_pin_23_;
  wire [0:0] cby_1__1__13_left_grid_pin_24_;
  wire [0:0] cby_1__1__13_left_grid_pin_25_;
  wire [0:0] cby_1__1__13_left_grid_pin_26_;
  wire [0:0] cby_1__1__13_left_grid_pin_27_;
  wire [0:0] cby_1__1__13_left_grid_pin_28_;
  wire [0:0] cby_1__1__13_left_grid_pin_29_;
  wire [0:0] cby_1__1__13_left_grid_pin_30_;
  wire [0:0] cby_1__1__13_left_grid_pin_31_;
  wire [0:0] cby_1__1__14_ccff_tail;
  wire [0:19] cby_1__1__14_chany_bottom_out;
  wire [0:19] cby_1__1__14_chany_top_out;
  wire [0:0] cby_1__1__14_left_grid_pin_16_;
  wire [0:0] cby_1__1__14_left_grid_pin_17_;
  wire [0:0] cby_1__1__14_left_grid_pin_18_;
  wire [0:0] cby_1__1__14_left_grid_pin_19_;
  wire [0:0] cby_1__1__14_left_grid_pin_20_;
  wire [0:0] cby_1__1__14_left_grid_pin_21_;
  wire [0:0] cby_1__1__14_left_grid_pin_22_;
  wire [0:0] cby_1__1__14_left_grid_pin_23_;
  wire [0:0] cby_1__1__14_left_grid_pin_24_;
  wire [0:0] cby_1__1__14_left_grid_pin_25_;
  wire [0:0] cby_1__1__14_left_grid_pin_26_;
  wire [0:0] cby_1__1__14_left_grid_pin_27_;
  wire [0:0] cby_1__1__14_left_grid_pin_28_;
  wire [0:0] cby_1__1__14_left_grid_pin_29_;
  wire [0:0] cby_1__1__14_left_grid_pin_30_;
  wire [0:0] cby_1__1__14_left_grid_pin_31_;
  wire [0:0] cby_1__1__15_ccff_tail;
  wire [0:19] cby_1__1__15_chany_bottom_out;
  wire [0:19] cby_1__1__15_chany_top_out;
  wire [0:0] cby_1__1__15_left_grid_pin_16_;
  wire [0:0] cby_1__1__15_left_grid_pin_17_;
  wire [0:0] cby_1__1__15_left_grid_pin_18_;
  wire [0:0] cby_1__1__15_left_grid_pin_19_;
  wire [0:0] cby_1__1__15_left_grid_pin_20_;
  wire [0:0] cby_1__1__15_left_grid_pin_21_;
  wire [0:0] cby_1__1__15_left_grid_pin_22_;
  wire [0:0] cby_1__1__15_left_grid_pin_23_;
  wire [0:0] cby_1__1__15_left_grid_pin_24_;
  wire [0:0] cby_1__1__15_left_grid_pin_25_;
  wire [0:0] cby_1__1__15_left_grid_pin_26_;
  wire [0:0] cby_1__1__15_left_grid_pin_27_;
  wire [0:0] cby_1__1__15_left_grid_pin_28_;
  wire [0:0] cby_1__1__15_left_grid_pin_29_;
  wire [0:0] cby_1__1__15_left_grid_pin_30_;
  wire [0:0] cby_1__1__15_left_grid_pin_31_;
  wire [0:0] cby_1__1__16_ccff_tail;
  wire [0:19] cby_1__1__16_chany_bottom_out;
  wire [0:19] cby_1__1__16_chany_top_out;
  wire [0:0] cby_1__1__16_left_grid_pin_16_;
  wire [0:0] cby_1__1__16_left_grid_pin_17_;
  wire [0:0] cby_1__1__16_left_grid_pin_18_;
  wire [0:0] cby_1__1__16_left_grid_pin_19_;
  wire [0:0] cby_1__1__16_left_grid_pin_20_;
  wire [0:0] cby_1__1__16_left_grid_pin_21_;
  wire [0:0] cby_1__1__16_left_grid_pin_22_;
  wire [0:0] cby_1__1__16_left_grid_pin_23_;
  wire [0:0] cby_1__1__16_left_grid_pin_24_;
  wire [0:0] cby_1__1__16_left_grid_pin_25_;
  wire [0:0] cby_1__1__16_left_grid_pin_26_;
  wire [0:0] cby_1__1__16_left_grid_pin_27_;
  wire [0:0] cby_1__1__16_left_grid_pin_28_;
  wire [0:0] cby_1__1__16_left_grid_pin_29_;
  wire [0:0] cby_1__1__16_left_grid_pin_30_;
  wire [0:0] cby_1__1__16_left_grid_pin_31_;
  wire [0:0] cby_1__1__17_ccff_tail;
  wire [0:19] cby_1__1__17_chany_bottom_out;
  wire [0:19] cby_1__1__17_chany_top_out;
  wire [0:0] cby_1__1__17_left_grid_pin_16_;
  wire [0:0] cby_1__1__17_left_grid_pin_17_;
  wire [0:0] cby_1__1__17_left_grid_pin_18_;
  wire [0:0] cby_1__1__17_left_grid_pin_19_;
  wire [0:0] cby_1__1__17_left_grid_pin_20_;
  wire [0:0] cby_1__1__17_left_grid_pin_21_;
  wire [0:0] cby_1__1__17_left_grid_pin_22_;
  wire [0:0] cby_1__1__17_left_grid_pin_23_;
  wire [0:0] cby_1__1__17_left_grid_pin_24_;
  wire [0:0] cby_1__1__17_left_grid_pin_25_;
  wire [0:0] cby_1__1__17_left_grid_pin_26_;
  wire [0:0] cby_1__1__17_left_grid_pin_27_;
  wire [0:0] cby_1__1__17_left_grid_pin_28_;
  wire [0:0] cby_1__1__17_left_grid_pin_29_;
  wire [0:0] cby_1__1__17_left_grid_pin_30_;
  wire [0:0] cby_1__1__17_left_grid_pin_31_;
  wire [0:0] cby_1__1__18_ccff_tail;
  wire [0:19] cby_1__1__18_chany_bottom_out;
  wire [0:19] cby_1__1__18_chany_top_out;
  wire [0:0] cby_1__1__18_left_grid_pin_16_;
  wire [0:0] cby_1__1__18_left_grid_pin_17_;
  wire [0:0] cby_1__1__18_left_grid_pin_18_;
  wire [0:0] cby_1__1__18_left_grid_pin_19_;
  wire [0:0] cby_1__1__18_left_grid_pin_20_;
  wire [0:0] cby_1__1__18_left_grid_pin_21_;
  wire [0:0] cby_1__1__18_left_grid_pin_22_;
  wire [0:0] cby_1__1__18_left_grid_pin_23_;
  wire [0:0] cby_1__1__18_left_grid_pin_24_;
  wire [0:0] cby_1__1__18_left_grid_pin_25_;
  wire [0:0] cby_1__1__18_left_grid_pin_26_;
  wire [0:0] cby_1__1__18_left_grid_pin_27_;
  wire [0:0] cby_1__1__18_left_grid_pin_28_;
  wire [0:0] cby_1__1__18_left_grid_pin_29_;
  wire [0:0] cby_1__1__18_left_grid_pin_30_;
  wire [0:0] cby_1__1__18_left_grid_pin_31_;
  wire [0:0] cby_1__1__19_ccff_tail;
  wire [0:19] cby_1__1__19_chany_bottom_out;
  wire [0:19] cby_1__1__19_chany_top_out;
  wire [0:0] cby_1__1__19_left_grid_pin_16_;
  wire [0:0] cby_1__1__19_left_grid_pin_17_;
  wire [0:0] cby_1__1__19_left_grid_pin_18_;
  wire [0:0] cby_1__1__19_left_grid_pin_19_;
  wire [0:0] cby_1__1__19_left_grid_pin_20_;
  wire [0:0] cby_1__1__19_left_grid_pin_21_;
  wire [0:0] cby_1__1__19_left_grid_pin_22_;
  wire [0:0] cby_1__1__19_left_grid_pin_23_;
  wire [0:0] cby_1__1__19_left_grid_pin_24_;
  wire [0:0] cby_1__1__19_left_grid_pin_25_;
  wire [0:0] cby_1__1__19_left_grid_pin_26_;
  wire [0:0] cby_1__1__19_left_grid_pin_27_;
  wire [0:0] cby_1__1__19_left_grid_pin_28_;
  wire [0:0] cby_1__1__19_left_grid_pin_29_;
  wire [0:0] cby_1__1__19_left_grid_pin_30_;
  wire [0:0] cby_1__1__19_left_grid_pin_31_;
  wire [0:0] cby_1__1__1_ccff_tail;
  wire [0:19] cby_1__1__1_chany_bottom_out;
  wire [0:19] cby_1__1__1_chany_top_out;
  wire [0:0] cby_1__1__1_left_grid_pin_16_;
  wire [0:0] cby_1__1__1_left_grid_pin_17_;
  wire [0:0] cby_1__1__1_left_grid_pin_18_;
  wire [0:0] cby_1__1__1_left_grid_pin_19_;
  wire [0:0] cby_1__1__1_left_grid_pin_20_;
  wire [0:0] cby_1__1__1_left_grid_pin_21_;
  wire [0:0] cby_1__1__1_left_grid_pin_22_;
  wire [0:0] cby_1__1__1_left_grid_pin_23_;
  wire [0:0] cby_1__1__1_left_grid_pin_24_;
  wire [0:0] cby_1__1__1_left_grid_pin_25_;
  wire [0:0] cby_1__1__1_left_grid_pin_26_;
  wire [0:0] cby_1__1__1_left_grid_pin_27_;
  wire [0:0] cby_1__1__1_left_grid_pin_28_;
  wire [0:0] cby_1__1__1_left_grid_pin_29_;
  wire [0:0] cby_1__1__1_left_grid_pin_30_;
  wire [0:0] cby_1__1__1_left_grid_pin_31_;
  wire [0:0] cby_1__1__20_ccff_tail;
  wire [0:19] cby_1__1__20_chany_bottom_out;
  wire [0:19] cby_1__1__20_chany_top_out;
  wire [0:0] cby_1__1__20_left_grid_pin_16_;
  wire [0:0] cby_1__1__20_left_grid_pin_17_;
  wire [0:0] cby_1__1__20_left_grid_pin_18_;
  wire [0:0] cby_1__1__20_left_grid_pin_19_;
  wire [0:0] cby_1__1__20_left_grid_pin_20_;
  wire [0:0] cby_1__1__20_left_grid_pin_21_;
  wire [0:0] cby_1__1__20_left_grid_pin_22_;
  wire [0:0] cby_1__1__20_left_grid_pin_23_;
  wire [0:0] cby_1__1__20_left_grid_pin_24_;
  wire [0:0] cby_1__1__20_left_grid_pin_25_;
  wire [0:0] cby_1__1__20_left_grid_pin_26_;
  wire [0:0] cby_1__1__20_left_grid_pin_27_;
  wire [0:0] cby_1__1__20_left_grid_pin_28_;
  wire [0:0] cby_1__1__20_left_grid_pin_29_;
  wire [0:0] cby_1__1__20_left_grid_pin_30_;
  wire [0:0] cby_1__1__20_left_grid_pin_31_;
  wire [0:0] cby_1__1__21_ccff_tail;
  wire [0:19] cby_1__1__21_chany_bottom_out;
  wire [0:19] cby_1__1__21_chany_top_out;
  wire [0:0] cby_1__1__21_left_grid_pin_16_;
  wire [0:0] cby_1__1__21_left_grid_pin_17_;
  wire [0:0] cby_1__1__21_left_grid_pin_18_;
  wire [0:0] cby_1__1__21_left_grid_pin_19_;
  wire [0:0] cby_1__1__21_left_grid_pin_20_;
  wire [0:0] cby_1__1__21_left_grid_pin_21_;
  wire [0:0] cby_1__1__21_left_grid_pin_22_;
  wire [0:0] cby_1__1__21_left_grid_pin_23_;
  wire [0:0] cby_1__1__21_left_grid_pin_24_;
  wire [0:0] cby_1__1__21_left_grid_pin_25_;
  wire [0:0] cby_1__1__21_left_grid_pin_26_;
  wire [0:0] cby_1__1__21_left_grid_pin_27_;
  wire [0:0] cby_1__1__21_left_grid_pin_28_;
  wire [0:0] cby_1__1__21_left_grid_pin_29_;
  wire [0:0] cby_1__1__21_left_grid_pin_30_;
  wire [0:0] cby_1__1__21_left_grid_pin_31_;
  wire [0:0] cby_1__1__22_ccff_tail;
  wire [0:19] cby_1__1__22_chany_bottom_out;
  wire [0:19] cby_1__1__22_chany_top_out;
  wire [0:0] cby_1__1__22_left_grid_pin_16_;
  wire [0:0] cby_1__1__22_left_grid_pin_17_;
  wire [0:0] cby_1__1__22_left_grid_pin_18_;
  wire [0:0] cby_1__1__22_left_grid_pin_19_;
  wire [0:0] cby_1__1__22_left_grid_pin_20_;
  wire [0:0] cby_1__1__22_left_grid_pin_21_;
  wire [0:0] cby_1__1__22_left_grid_pin_22_;
  wire [0:0] cby_1__1__22_left_grid_pin_23_;
  wire [0:0] cby_1__1__22_left_grid_pin_24_;
  wire [0:0] cby_1__1__22_left_grid_pin_25_;
  wire [0:0] cby_1__1__22_left_grid_pin_26_;
  wire [0:0] cby_1__1__22_left_grid_pin_27_;
  wire [0:0] cby_1__1__22_left_grid_pin_28_;
  wire [0:0] cby_1__1__22_left_grid_pin_29_;
  wire [0:0] cby_1__1__22_left_grid_pin_30_;
  wire [0:0] cby_1__1__22_left_grid_pin_31_;
  wire [0:0] cby_1__1__23_ccff_tail;
  wire [0:19] cby_1__1__23_chany_bottom_out;
  wire [0:19] cby_1__1__23_chany_top_out;
  wire [0:0] cby_1__1__23_left_grid_pin_16_;
  wire [0:0] cby_1__1__23_left_grid_pin_17_;
  wire [0:0] cby_1__1__23_left_grid_pin_18_;
  wire [0:0] cby_1__1__23_left_grid_pin_19_;
  wire [0:0] cby_1__1__23_left_grid_pin_20_;
  wire [0:0] cby_1__1__23_left_grid_pin_21_;
  wire [0:0] cby_1__1__23_left_grid_pin_22_;
  wire [0:0] cby_1__1__23_left_grid_pin_23_;
  wire [0:0] cby_1__1__23_left_grid_pin_24_;
  wire [0:0] cby_1__1__23_left_grid_pin_25_;
  wire [0:0] cby_1__1__23_left_grid_pin_26_;
  wire [0:0] cby_1__1__23_left_grid_pin_27_;
  wire [0:0] cby_1__1__23_left_grid_pin_28_;
  wire [0:0] cby_1__1__23_left_grid_pin_29_;
  wire [0:0] cby_1__1__23_left_grid_pin_30_;
  wire [0:0] cby_1__1__23_left_grid_pin_31_;
  wire [0:0] cby_1__1__24_ccff_tail;
  wire [0:19] cby_1__1__24_chany_bottom_out;
  wire [0:19] cby_1__1__24_chany_top_out;
  wire [0:0] cby_1__1__24_left_grid_pin_16_;
  wire [0:0] cby_1__1__24_left_grid_pin_17_;
  wire [0:0] cby_1__1__24_left_grid_pin_18_;
  wire [0:0] cby_1__1__24_left_grid_pin_19_;
  wire [0:0] cby_1__1__24_left_grid_pin_20_;
  wire [0:0] cby_1__1__24_left_grid_pin_21_;
  wire [0:0] cby_1__1__24_left_grid_pin_22_;
  wire [0:0] cby_1__1__24_left_grid_pin_23_;
  wire [0:0] cby_1__1__24_left_grid_pin_24_;
  wire [0:0] cby_1__1__24_left_grid_pin_25_;
  wire [0:0] cby_1__1__24_left_grid_pin_26_;
  wire [0:0] cby_1__1__24_left_grid_pin_27_;
  wire [0:0] cby_1__1__24_left_grid_pin_28_;
  wire [0:0] cby_1__1__24_left_grid_pin_29_;
  wire [0:0] cby_1__1__24_left_grid_pin_30_;
  wire [0:0] cby_1__1__24_left_grid_pin_31_;
  wire [0:0] cby_1__1__25_ccff_tail;
  wire [0:19] cby_1__1__25_chany_bottom_out;
  wire [0:19] cby_1__1__25_chany_top_out;
  wire [0:0] cby_1__1__25_left_grid_pin_16_;
  wire [0:0] cby_1__1__25_left_grid_pin_17_;
  wire [0:0] cby_1__1__25_left_grid_pin_18_;
  wire [0:0] cby_1__1__25_left_grid_pin_19_;
  wire [0:0] cby_1__1__25_left_grid_pin_20_;
  wire [0:0] cby_1__1__25_left_grid_pin_21_;
  wire [0:0] cby_1__1__25_left_grid_pin_22_;
  wire [0:0] cby_1__1__25_left_grid_pin_23_;
  wire [0:0] cby_1__1__25_left_grid_pin_24_;
  wire [0:0] cby_1__1__25_left_grid_pin_25_;
  wire [0:0] cby_1__1__25_left_grid_pin_26_;
  wire [0:0] cby_1__1__25_left_grid_pin_27_;
  wire [0:0] cby_1__1__25_left_grid_pin_28_;
  wire [0:0] cby_1__1__25_left_grid_pin_29_;
  wire [0:0] cby_1__1__25_left_grid_pin_30_;
  wire [0:0] cby_1__1__25_left_grid_pin_31_;
  wire [0:0] cby_1__1__26_ccff_tail;
  wire [0:19] cby_1__1__26_chany_bottom_out;
  wire [0:19] cby_1__1__26_chany_top_out;
  wire [0:0] cby_1__1__26_left_grid_pin_16_;
  wire [0:0] cby_1__1__26_left_grid_pin_17_;
  wire [0:0] cby_1__1__26_left_grid_pin_18_;
  wire [0:0] cby_1__1__26_left_grid_pin_19_;
  wire [0:0] cby_1__1__26_left_grid_pin_20_;
  wire [0:0] cby_1__1__26_left_grid_pin_21_;
  wire [0:0] cby_1__1__26_left_grid_pin_22_;
  wire [0:0] cby_1__1__26_left_grid_pin_23_;
  wire [0:0] cby_1__1__26_left_grid_pin_24_;
  wire [0:0] cby_1__1__26_left_grid_pin_25_;
  wire [0:0] cby_1__1__26_left_grid_pin_26_;
  wire [0:0] cby_1__1__26_left_grid_pin_27_;
  wire [0:0] cby_1__1__26_left_grid_pin_28_;
  wire [0:0] cby_1__1__26_left_grid_pin_29_;
  wire [0:0] cby_1__1__26_left_grid_pin_30_;
  wire [0:0] cby_1__1__26_left_grid_pin_31_;
  wire [0:0] cby_1__1__27_ccff_tail;
  wire [0:19] cby_1__1__27_chany_bottom_out;
  wire [0:19] cby_1__1__27_chany_top_out;
  wire [0:0] cby_1__1__27_left_grid_pin_16_;
  wire [0:0] cby_1__1__27_left_grid_pin_17_;
  wire [0:0] cby_1__1__27_left_grid_pin_18_;
  wire [0:0] cby_1__1__27_left_grid_pin_19_;
  wire [0:0] cby_1__1__27_left_grid_pin_20_;
  wire [0:0] cby_1__1__27_left_grid_pin_21_;
  wire [0:0] cby_1__1__27_left_grid_pin_22_;
  wire [0:0] cby_1__1__27_left_grid_pin_23_;
  wire [0:0] cby_1__1__27_left_grid_pin_24_;
  wire [0:0] cby_1__1__27_left_grid_pin_25_;
  wire [0:0] cby_1__1__27_left_grid_pin_26_;
  wire [0:0] cby_1__1__27_left_grid_pin_27_;
  wire [0:0] cby_1__1__27_left_grid_pin_28_;
  wire [0:0] cby_1__1__27_left_grid_pin_29_;
  wire [0:0] cby_1__1__27_left_grid_pin_30_;
  wire [0:0] cby_1__1__27_left_grid_pin_31_;
  wire [0:0] cby_1__1__28_ccff_tail;
  wire [0:19] cby_1__1__28_chany_bottom_out;
  wire [0:19] cby_1__1__28_chany_top_out;
  wire [0:0] cby_1__1__28_left_grid_pin_16_;
  wire [0:0] cby_1__1__28_left_grid_pin_17_;
  wire [0:0] cby_1__1__28_left_grid_pin_18_;
  wire [0:0] cby_1__1__28_left_grid_pin_19_;
  wire [0:0] cby_1__1__28_left_grid_pin_20_;
  wire [0:0] cby_1__1__28_left_grid_pin_21_;
  wire [0:0] cby_1__1__28_left_grid_pin_22_;
  wire [0:0] cby_1__1__28_left_grid_pin_23_;
  wire [0:0] cby_1__1__28_left_grid_pin_24_;
  wire [0:0] cby_1__1__28_left_grid_pin_25_;
  wire [0:0] cby_1__1__28_left_grid_pin_26_;
  wire [0:0] cby_1__1__28_left_grid_pin_27_;
  wire [0:0] cby_1__1__28_left_grid_pin_28_;
  wire [0:0] cby_1__1__28_left_grid_pin_29_;
  wire [0:0] cby_1__1__28_left_grid_pin_30_;
  wire [0:0] cby_1__1__28_left_grid_pin_31_;
  wire [0:0] cby_1__1__29_ccff_tail;
  wire [0:19] cby_1__1__29_chany_bottom_out;
  wire [0:19] cby_1__1__29_chany_top_out;
  wire [0:0] cby_1__1__29_left_grid_pin_16_;
  wire [0:0] cby_1__1__29_left_grid_pin_17_;
  wire [0:0] cby_1__1__29_left_grid_pin_18_;
  wire [0:0] cby_1__1__29_left_grid_pin_19_;
  wire [0:0] cby_1__1__29_left_grid_pin_20_;
  wire [0:0] cby_1__1__29_left_grid_pin_21_;
  wire [0:0] cby_1__1__29_left_grid_pin_22_;
  wire [0:0] cby_1__1__29_left_grid_pin_23_;
  wire [0:0] cby_1__1__29_left_grid_pin_24_;
  wire [0:0] cby_1__1__29_left_grid_pin_25_;
  wire [0:0] cby_1__1__29_left_grid_pin_26_;
  wire [0:0] cby_1__1__29_left_grid_pin_27_;
  wire [0:0] cby_1__1__29_left_grid_pin_28_;
  wire [0:0] cby_1__1__29_left_grid_pin_29_;
  wire [0:0] cby_1__1__29_left_grid_pin_30_;
  wire [0:0] cby_1__1__29_left_grid_pin_31_;
  wire [0:0] cby_1__1__2_ccff_tail;
  wire [0:19] cby_1__1__2_chany_bottom_out;
  wire [0:19] cby_1__1__2_chany_top_out;
  wire [0:0] cby_1__1__2_left_grid_pin_16_;
  wire [0:0] cby_1__1__2_left_grid_pin_17_;
  wire [0:0] cby_1__1__2_left_grid_pin_18_;
  wire [0:0] cby_1__1__2_left_grid_pin_19_;
  wire [0:0] cby_1__1__2_left_grid_pin_20_;
  wire [0:0] cby_1__1__2_left_grid_pin_21_;
  wire [0:0] cby_1__1__2_left_grid_pin_22_;
  wire [0:0] cby_1__1__2_left_grid_pin_23_;
  wire [0:0] cby_1__1__2_left_grid_pin_24_;
  wire [0:0] cby_1__1__2_left_grid_pin_25_;
  wire [0:0] cby_1__1__2_left_grid_pin_26_;
  wire [0:0] cby_1__1__2_left_grid_pin_27_;
  wire [0:0] cby_1__1__2_left_grid_pin_28_;
  wire [0:0] cby_1__1__2_left_grid_pin_29_;
  wire [0:0] cby_1__1__2_left_grid_pin_30_;
  wire [0:0] cby_1__1__2_left_grid_pin_31_;
  wire [0:0] cby_1__1__30_ccff_tail;
  wire [0:19] cby_1__1__30_chany_bottom_out;
  wire [0:19] cby_1__1__30_chany_top_out;
  wire [0:0] cby_1__1__30_left_grid_pin_16_;
  wire [0:0] cby_1__1__30_left_grid_pin_17_;
  wire [0:0] cby_1__1__30_left_grid_pin_18_;
  wire [0:0] cby_1__1__30_left_grid_pin_19_;
  wire [0:0] cby_1__1__30_left_grid_pin_20_;
  wire [0:0] cby_1__1__30_left_grid_pin_21_;
  wire [0:0] cby_1__1__30_left_grid_pin_22_;
  wire [0:0] cby_1__1__30_left_grid_pin_23_;
  wire [0:0] cby_1__1__30_left_grid_pin_24_;
  wire [0:0] cby_1__1__30_left_grid_pin_25_;
  wire [0:0] cby_1__1__30_left_grid_pin_26_;
  wire [0:0] cby_1__1__30_left_grid_pin_27_;
  wire [0:0] cby_1__1__30_left_grid_pin_28_;
  wire [0:0] cby_1__1__30_left_grid_pin_29_;
  wire [0:0] cby_1__1__30_left_grid_pin_30_;
  wire [0:0] cby_1__1__30_left_grid_pin_31_;
  wire [0:0] cby_1__1__31_ccff_tail;
  wire [0:19] cby_1__1__31_chany_bottom_out;
  wire [0:19] cby_1__1__31_chany_top_out;
  wire [0:0] cby_1__1__31_left_grid_pin_16_;
  wire [0:0] cby_1__1__31_left_grid_pin_17_;
  wire [0:0] cby_1__1__31_left_grid_pin_18_;
  wire [0:0] cby_1__1__31_left_grid_pin_19_;
  wire [0:0] cby_1__1__31_left_grid_pin_20_;
  wire [0:0] cby_1__1__31_left_grid_pin_21_;
  wire [0:0] cby_1__1__31_left_grid_pin_22_;
  wire [0:0] cby_1__1__31_left_grid_pin_23_;
  wire [0:0] cby_1__1__31_left_grid_pin_24_;
  wire [0:0] cby_1__1__31_left_grid_pin_25_;
  wire [0:0] cby_1__1__31_left_grid_pin_26_;
  wire [0:0] cby_1__1__31_left_grid_pin_27_;
  wire [0:0] cby_1__1__31_left_grid_pin_28_;
  wire [0:0] cby_1__1__31_left_grid_pin_29_;
  wire [0:0] cby_1__1__31_left_grid_pin_30_;
  wire [0:0] cby_1__1__31_left_grid_pin_31_;
  wire [0:0] cby_1__1__32_ccff_tail;
  wire [0:19] cby_1__1__32_chany_bottom_out;
  wire [0:19] cby_1__1__32_chany_top_out;
  wire [0:0] cby_1__1__32_left_grid_pin_16_;
  wire [0:0] cby_1__1__32_left_grid_pin_17_;
  wire [0:0] cby_1__1__32_left_grid_pin_18_;
  wire [0:0] cby_1__1__32_left_grid_pin_19_;
  wire [0:0] cby_1__1__32_left_grid_pin_20_;
  wire [0:0] cby_1__1__32_left_grid_pin_21_;
  wire [0:0] cby_1__1__32_left_grid_pin_22_;
  wire [0:0] cby_1__1__32_left_grid_pin_23_;
  wire [0:0] cby_1__1__32_left_grid_pin_24_;
  wire [0:0] cby_1__1__32_left_grid_pin_25_;
  wire [0:0] cby_1__1__32_left_grid_pin_26_;
  wire [0:0] cby_1__1__32_left_grid_pin_27_;
  wire [0:0] cby_1__1__32_left_grid_pin_28_;
  wire [0:0] cby_1__1__32_left_grid_pin_29_;
  wire [0:0] cby_1__1__32_left_grid_pin_30_;
  wire [0:0] cby_1__1__32_left_grid_pin_31_;
  wire [0:0] cby_1__1__33_ccff_tail;
  wire [0:19] cby_1__1__33_chany_bottom_out;
  wire [0:19] cby_1__1__33_chany_top_out;
  wire [0:0] cby_1__1__33_left_grid_pin_16_;
  wire [0:0] cby_1__1__33_left_grid_pin_17_;
  wire [0:0] cby_1__1__33_left_grid_pin_18_;
  wire [0:0] cby_1__1__33_left_grid_pin_19_;
  wire [0:0] cby_1__1__33_left_grid_pin_20_;
  wire [0:0] cby_1__1__33_left_grid_pin_21_;
  wire [0:0] cby_1__1__33_left_grid_pin_22_;
  wire [0:0] cby_1__1__33_left_grid_pin_23_;
  wire [0:0] cby_1__1__33_left_grid_pin_24_;
  wire [0:0] cby_1__1__33_left_grid_pin_25_;
  wire [0:0] cby_1__1__33_left_grid_pin_26_;
  wire [0:0] cby_1__1__33_left_grid_pin_27_;
  wire [0:0] cby_1__1__33_left_grid_pin_28_;
  wire [0:0] cby_1__1__33_left_grid_pin_29_;
  wire [0:0] cby_1__1__33_left_grid_pin_30_;
  wire [0:0] cby_1__1__33_left_grid_pin_31_;
  wire [0:0] cby_1__1__34_ccff_tail;
  wire [0:19] cby_1__1__34_chany_bottom_out;
  wire [0:19] cby_1__1__34_chany_top_out;
  wire [0:0] cby_1__1__34_left_grid_pin_16_;
  wire [0:0] cby_1__1__34_left_grid_pin_17_;
  wire [0:0] cby_1__1__34_left_grid_pin_18_;
  wire [0:0] cby_1__1__34_left_grid_pin_19_;
  wire [0:0] cby_1__1__34_left_grid_pin_20_;
  wire [0:0] cby_1__1__34_left_grid_pin_21_;
  wire [0:0] cby_1__1__34_left_grid_pin_22_;
  wire [0:0] cby_1__1__34_left_grid_pin_23_;
  wire [0:0] cby_1__1__34_left_grid_pin_24_;
  wire [0:0] cby_1__1__34_left_grid_pin_25_;
  wire [0:0] cby_1__1__34_left_grid_pin_26_;
  wire [0:0] cby_1__1__34_left_grid_pin_27_;
  wire [0:0] cby_1__1__34_left_grid_pin_28_;
  wire [0:0] cby_1__1__34_left_grid_pin_29_;
  wire [0:0] cby_1__1__34_left_grid_pin_30_;
  wire [0:0] cby_1__1__34_left_grid_pin_31_;
  wire [0:0] cby_1__1__35_ccff_tail;
  wire [0:19] cby_1__1__35_chany_bottom_out;
  wire [0:19] cby_1__1__35_chany_top_out;
  wire [0:0] cby_1__1__35_left_grid_pin_16_;
  wire [0:0] cby_1__1__35_left_grid_pin_17_;
  wire [0:0] cby_1__1__35_left_grid_pin_18_;
  wire [0:0] cby_1__1__35_left_grid_pin_19_;
  wire [0:0] cby_1__1__35_left_grid_pin_20_;
  wire [0:0] cby_1__1__35_left_grid_pin_21_;
  wire [0:0] cby_1__1__35_left_grid_pin_22_;
  wire [0:0] cby_1__1__35_left_grid_pin_23_;
  wire [0:0] cby_1__1__35_left_grid_pin_24_;
  wire [0:0] cby_1__1__35_left_grid_pin_25_;
  wire [0:0] cby_1__1__35_left_grid_pin_26_;
  wire [0:0] cby_1__1__35_left_grid_pin_27_;
  wire [0:0] cby_1__1__35_left_grid_pin_28_;
  wire [0:0] cby_1__1__35_left_grid_pin_29_;
  wire [0:0] cby_1__1__35_left_grid_pin_30_;
  wire [0:0] cby_1__1__35_left_grid_pin_31_;
  wire [0:0] cby_1__1__36_ccff_tail;
  wire [0:19] cby_1__1__36_chany_bottom_out;
  wire [0:19] cby_1__1__36_chany_top_out;
  wire [0:0] cby_1__1__36_left_grid_pin_16_;
  wire [0:0] cby_1__1__36_left_grid_pin_17_;
  wire [0:0] cby_1__1__36_left_grid_pin_18_;
  wire [0:0] cby_1__1__36_left_grid_pin_19_;
  wire [0:0] cby_1__1__36_left_grid_pin_20_;
  wire [0:0] cby_1__1__36_left_grid_pin_21_;
  wire [0:0] cby_1__1__36_left_grid_pin_22_;
  wire [0:0] cby_1__1__36_left_grid_pin_23_;
  wire [0:0] cby_1__1__36_left_grid_pin_24_;
  wire [0:0] cby_1__1__36_left_grid_pin_25_;
  wire [0:0] cby_1__1__36_left_grid_pin_26_;
  wire [0:0] cby_1__1__36_left_grid_pin_27_;
  wire [0:0] cby_1__1__36_left_grid_pin_28_;
  wire [0:0] cby_1__1__36_left_grid_pin_29_;
  wire [0:0] cby_1__1__36_left_grid_pin_30_;
  wire [0:0] cby_1__1__36_left_grid_pin_31_;
  wire [0:0] cby_1__1__37_ccff_tail;
  wire [0:19] cby_1__1__37_chany_bottom_out;
  wire [0:19] cby_1__1__37_chany_top_out;
  wire [0:0] cby_1__1__37_left_grid_pin_16_;
  wire [0:0] cby_1__1__37_left_grid_pin_17_;
  wire [0:0] cby_1__1__37_left_grid_pin_18_;
  wire [0:0] cby_1__1__37_left_grid_pin_19_;
  wire [0:0] cby_1__1__37_left_grid_pin_20_;
  wire [0:0] cby_1__1__37_left_grid_pin_21_;
  wire [0:0] cby_1__1__37_left_grid_pin_22_;
  wire [0:0] cby_1__1__37_left_grid_pin_23_;
  wire [0:0] cby_1__1__37_left_grid_pin_24_;
  wire [0:0] cby_1__1__37_left_grid_pin_25_;
  wire [0:0] cby_1__1__37_left_grid_pin_26_;
  wire [0:0] cby_1__1__37_left_grid_pin_27_;
  wire [0:0] cby_1__1__37_left_grid_pin_28_;
  wire [0:0] cby_1__1__37_left_grid_pin_29_;
  wire [0:0] cby_1__1__37_left_grid_pin_30_;
  wire [0:0] cby_1__1__37_left_grid_pin_31_;
  wire [0:0] cby_1__1__38_ccff_tail;
  wire [0:19] cby_1__1__38_chany_bottom_out;
  wire [0:19] cby_1__1__38_chany_top_out;
  wire [0:0] cby_1__1__38_left_grid_pin_16_;
  wire [0:0] cby_1__1__38_left_grid_pin_17_;
  wire [0:0] cby_1__1__38_left_grid_pin_18_;
  wire [0:0] cby_1__1__38_left_grid_pin_19_;
  wire [0:0] cby_1__1__38_left_grid_pin_20_;
  wire [0:0] cby_1__1__38_left_grid_pin_21_;
  wire [0:0] cby_1__1__38_left_grid_pin_22_;
  wire [0:0] cby_1__1__38_left_grid_pin_23_;
  wire [0:0] cby_1__1__38_left_grid_pin_24_;
  wire [0:0] cby_1__1__38_left_grid_pin_25_;
  wire [0:0] cby_1__1__38_left_grid_pin_26_;
  wire [0:0] cby_1__1__38_left_grid_pin_27_;
  wire [0:0] cby_1__1__38_left_grid_pin_28_;
  wire [0:0] cby_1__1__38_left_grid_pin_29_;
  wire [0:0] cby_1__1__38_left_grid_pin_30_;
  wire [0:0] cby_1__1__38_left_grid_pin_31_;
  wire [0:0] cby_1__1__39_ccff_tail;
  wire [0:19] cby_1__1__39_chany_bottom_out;
  wire [0:19] cby_1__1__39_chany_top_out;
  wire [0:0] cby_1__1__39_left_grid_pin_16_;
  wire [0:0] cby_1__1__39_left_grid_pin_17_;
  wire [0:0] cby_1__1__39_left_grid_pin_18_;
  wire [0:0] cby_1__1__39_left_grid_pin_19_;
  wire [0:0] cby_1__1__39_left_grid_pin_20_;
  wire [0:0] cby_1__1__39_left_grid_pin_21_;
  wire [0:0] cby_1__1__39_left_grid_pin_22_;
  wire [0:0] cby_1__1__39_left_grid_pin_23_;
  wire [0:0] cby_1__1__39_left_grid_pin_24_;
  wire [0:0] cby_1__1__39_left_grid_pin_25_;
  wire [0:0] cby_1__1__39_left_grid_pin_26_;
  wire [0:0] cby_1__1__39_left_grid_pin_27_;
  wire [0:0] cby_1__1__39_left_grid_pin_28_;
  wire [0:0] cby_1__1__39_left_grid_pin_29_;
  wire [0:0] cby_1__1__39_left_grid_pin_30_;
  wire [0:0] cby_1__1__39_left_grid_pin_31_;
  wire [0:0] cby_1__1__3_ccff_tail;
  wire [0:19] cby_1__1__3_chany_bottom_out;
  wire [0:19] cby_1__1__3_chany_top_out;
  wire [0:0] cby_1__1__3_left_grid_pin_16_;
  wire [0:0] cby_1__1__3_left_grid_pin_17_;
  wire [0:0] cby_1__1__3_left_grid_pin_18_;
  wire [0:0] cby_1__1__3_left_grid_pin_19_;
  wire [0:0] cby_1__1__3_left_grid_pin_20_;
  wire [0:0] cby_1__1__3_left_grid_pin_21_;
  wire [0:0] cby_1__1__3_left_grid_pin_22_;
  wire [0:0] cby_1__1__3_left_grid_pin_23_;
  wire [0:0] cby_1__1__3_left_grid_pin_24_;
  wire [0:0] cby_1__1__3_left_grid_pin_25_;
  wire [0:0] cby_1__1__3_left_grid_pin_26_;
  wire [0:0] cby_1__1__3_left_grid_pin_27_;
  wire [0:0] cby_1__1__3_left_grid_pin_28_;
  wire [0:0] cby_1__1__3_left_grid_pin_29_;
  wire [0:0] cby_1__1__3_left_grid_pin_30_;
  wire [0:0] cby_1__1__3_left_grid_pin_31_;
  wire [0:0] cby_1__1__40_ccff_tail;
  wire [0:19] cby_1__1__40_chany_bottom_out;
  wire [0:19] cby_1__1__40_chany_top_out;
  wire [0:0] cby_1__1__40_left_grid_pin_16_;
  wire [0:0] cby_1__1__40_left_grid_pin_17_;
  wire [0:0] cby_1__1__40_left_grid_pin_18_;
  wire [0:0] cby_1__1__40_left_grid_pin_19_;
  wire [0:0] cby_1__1__40_left_grid_pin_20_;
  wire [0:0] cby_1__1__40_left_grid_pin_21_;
  wire [0:0] cby_1__1__40_left_grid_pin_22_;
  wire [0:0] cby_1__1__40_left_grid_pin_23_;
  wire [0:0] cby_1__1__40_left_grid_pin_24_;
  wire [0:0] cby_1__1__40_left_grid_pin_25_;
  wire [0:0] cby_1__1__40_left_grid_pin_26_;
  wire [0:0] cby_1__1__40_left_grid_pin_27_;
  wire [0:0] cby_1__1__40_left_grid_pin_28_;
  wire [0:0] cby_1__1__40_left_grid_pin_29_;
  wire [0:0] cby_1__1__40_left_grid_pin_30_;
  wire [0:0] cby_1__1__40_left_grid_pin_31_;
  wire [0:0] cby_1__1__41_ccff_tail;
  wire [0:19] cby_1__1__41_chany_bottom_out;
  wire [0:19] cby_1__1__41_chany_top_out;
  wire [0:0] cby_1__1__41_left_grid_pin_16_;
  wire [0:0] cby_1__1__41_left_grid_pin_17_;
  wire [0:0] cby_1__1__41_left_grid_pin_18_;
  wire [0:0] cby_1__1__41_left_grid_pin_19_;
  wire [0:0] cby_1__1__41_left_grid_pin_20_;
  wire [0:0] cby_1__1__41_left_grid_pin_21_;
  wire [0:0] cby_1__1__41_left_grid_pin_22_;
  wire [0:0] cby_1__1__41_left_grid_pin_23_;
  wire [0:0] cby_1__1__41_left_grid_pin_24_;
  wire [0:0] cby_1__1__41_left_grid_pin_25_;
  wire [0:0] cby_1__1__41_left_grid_pin_26_;
  wire [0:0] cby_1__1__41_left_grid_pin_27_;
  wire [0:0] cby_1__1__41_left_grid_pin_28_;
  wire [0:0] cby_1__1__41_left_grid_pin_29_;
  wire [0:0] cby_1__1__41_left_grid_pin_30_;
  wire [0:0] cby_1__1__41_left_grid_pin_31_;
  wire [0:0] cby_1__1__42_ccff_tail;
  wire [0:19] cby_1__1__42_chany_bottom_out;
  wire [0:19] cby_1__1__42_chany_top_out;
  wire [0:0] cby_1__1__42_left_grid_pin_16_;
  wire [0:0] cby_1__1__42_left_grid_pin_17_;
  wire [0:0] cby_1__1__42_left_grid_pin_18_;
  wire [0:0] cby_1__1__42_left_grid_pin_19_;
  wire [0:0] cby_1__1__42_left_grid_pin_20_;
  wire [0:0] cby_1__1__42_left_grid_pin_21_;
  wire [0:0] cby_1__1__42_left_grid_pin_22_;
  wire [0:0] cby_1__1__42_left_grid_pin_23_;
  wire [0:0] cby_1__1__42_left_grid_pin_24_;
  wire [0:0] cby_1__1__42_left_grid_pin_25_;
  wire [0:0] cby_1__1__42_left_grid_pin_26_;
  wire [0:0] cby_1__1__42_left_grid_pin_27_;
  wire [0:0] cby_1__1__42_left_grid_pin_28_;
  wire [0:0] cby_1__1__42_left_grid_pin_29_;
  wire [0:0] cby_1__1__42_left_grid_pin_30_;
  wire [0:0] cby_1__1__42_left_grid_pin_31_;
  wire [0:0] cby_1__1__43_ccff_tail;
  wire [0:19] cby_1__1__43_chany_bottom_out;
  wire [0:19] cby_1__1__43_chany_top_out;
  wire [0:0] cby_1__1__43_left_grid_pin_16_;
  wire [0:0] cby_1__1__43_left_grid_pin_17_;
  wire [0:0] cby_1__1__43_left_grid_pin_18_;
  wire [0:0] cby_1__1__43_left_grid_pin_19_;
  wire [0:0] cby_1__1__43_left_grid_pin_20_;
  wire [0:0] cby_1__1__43_left_grid_pin_21_;
  wire [0:0] cby_1__1__43_left_grid_pin_22_;
  wire [0:0] cby_1__1__43_left_grid_pin_23_;
  wire [0:0] cby_1__1__43_left_grid_pin_24_;
  wire [0:0] cby_1__1__43_left_grid_pin_25_;
  wire [0:0] cby_1__1__43_left_grid_pin_26_;
  wire [0:0] cby_1__1__43_left_grid_pin_27_;
  wire [0:0] cby_1__1__43_left_grid_pin_28_;
  wire [0:0] cby_1__1__43_left_grid_pin_29_;
  wire [0:0] cby_1__1__43_left_grid_pin_30_;
  wire [0:0] cby_1__1__43_left_grid_pin_31_;
  wire [0:0] cby_1__1__44_ccff_tail;
  wire [0:19] cby_1__1__44_chany_bottom_out;
  wire [0:19] cby_1__1__44_chany_top_out;
  wire [0:0] cby_1__1__44_left_grid_pin_16_;
  wire [0:0] cby_1__1__44_left_grid_pin_17_;
  wire [0:0] cby_1__1__44_left_grid_pin_18_;
  wire [0:0] cby_1__1__44_left_grid_pin_19_;
  wire [0:0] cby_1__1__44_left_grid_pin_20_;
  wire [0:0] cby_1__1__44_left_grid_pin_21_;
  wire [0:0] cby_1__1__44_left_grid_pin_22_;
  wire [0:0] cby_1__1__44_left_grid_pin_23_;
  wire [0:0] cby_1__1__44_left_grid_pin_24_;
  wire [0:0] cby_1__1__44_left_grid_pin_25_;
  wire [0:0] cby_1__1__44_left_grid_pin_26_;
  wire [0:0] cby_1__1__44_left_grid_pin_27_;
  wire [0:0] cby_1__1__44_left_grid_pin_28_;
  wire [0:0] cby_1__1__44_left_grid_pin_29_;
  wire [0:0] cby_1__1__44_left_grid_pin_30_;
  wire [0:0] cby_1__1__44_left_grid_pin_31_;
  wire [0:0] cby_1__1__45_ccff_tail;
  wire [0:19] cby_1__1__45_chany_bottom_out;
  wire [0:19] cby_1__1__45_chany_top_out;
  wire [0:0] cby_1__1__45_left_grid_pin_16_;
  wire [0:0] cby_1__1__45_left_grid_pin_17_;
  wire [0:0] cby_1__1__45_left_grid_pin_18_;
  wire [0:0] cby_1__1__45_left_grid_pin_19_;
  wire [0:0] cby_1__1__45_left_grid_pin_20_;
  wire [0:0] cby_1__1__45_left_grid_pin_21_;
  wire [0:0] cby_1__1__45_left_grid_pin_22_;
  wire [0:0] cby_1__1__45_left_grid_pin_23_;
  wire [0:0] cby_1__1__45_left_grid_pin_24_;
  wire [0:0] cby_1__1__45_left_grid_pin_25_;
  wire [0:0] cby_1__1__45_left_grid_pin_26_;
  wire [0:0] cby_1__1__45_left_grid_pin_27_;
  wire [0:0] cby_1__1__45_left_grid_pin_28_;
  wire [0:0] cby_1__1__45_left_grid_pin_29_;
  wire [0:0] cby_1__1__45_left_grid_pin_30_;
  wire [0:0] cby_1__1__45_left_grid_pin_31_;
  wire [0:0] cby_1__1__46_ccff_tail;
  wire [0:19] cby_1__1__46_chany_bottom_out;
  wire [0:19] cby_1__1__46_chany_top_out;
  wire [0:0] cby_1__1__46_left_grid_pin_16_;
  wire [0:0] cby_1__1__46_left_grid_pin_17_;
  wire [0:0] cby_1__1__46_left_grid_pin_18_;
  wire [0:0] cby_1__1__46_left_grid_pin_19_;
  wire [0:0] cby_1__1__46_left_grid_pin_20_;
  wire [0:0] cby_1__1__46_left_grid_pin_21_;
  wire [0:0] cby_1__1__46_left_grid_pin_22_;
  wire [0:0] cby_1__1__46_left_grid_pin_23_;
  wire [0:0] cby_1__1__46_left_grid_pin_24_;
  wire [0:0] cby_1__1__46_left_grid_pin_25_;
  wire [0:0] cby_1__1__46_left_grid_pin_26_;
  wire [0:0] cby_1__1__46_left_grid_pin_27_;
  wire [0:0] cby_1__1__46_left_grid_pin_28_;
  wire [0:0] cby_1__1__46_left_grid_pin_29_;
  wire [0:0] cby_1__1__46_left_grid_pin_30_;
  wire [0:0] cby_1__1__46_left_grid_pin_31_;
  wire [0:0] cby_1__1__47_ccff_tail;
  wire [0:19] cby_1__1__47_chany_bottom_out;
  wire [0:19] cby_1__1__47_chany_top_out;
  wire [0:0] cby_1__1__47_left_grid_pin_16_;
  wire [0:0] cby_1__1__47_left_grid_pin_17_;
  wire [0:0] cby_1__1__47_left_grid_pin_18_;
  wire [0:0] cby_1__1__47_left_grid_pin_19_;
  wire [0:0] cby_1__1__47_left_grid_pin_20_;
  wire [0:0] cby_1__1__47_left_grid_pin_21_;
  wire [0:0] cby_1__1__47_left_grid_pin_22_;
  wire [0:0] cby_1__1__47_left_grid_pin_23_;
  wire [0:0] cby_1__1__47_left_grid_pin_24_;
  wire [0:0] cby_1__1__47_left_grid_pin_25_;
  wire [0:0] cby_1__1__47_left_grid_pin_26_;
  wire [0:0] cby_1__1__47_left_grid_pin_27_;
  wire [0:0] cby_1__1__47_left_grid_pin_28_;
  wire [0:0] cby_1__1__47_left_grid_pin_29_;
  wire [0:0] cby_1__1__47_left_grid_pin_30_;
  wire [0:0] cby_1__1__47_left_grid_pin_31_;
  wire [0:0] cby_1__1__48_ccff_tail;
  wire [0:19] cby_1__1__48_chany_bottom_out;
  wire [0:19] cby_1__1__48_chany_top_out;
  wire [0:0] cby_1__1__48_left_grid_pin_16_;
  wire [0:0] cby_1__1__48_left_grid_pin_17_;
  wire [0:0] cby_1__1__48_left_grid_pin_18_;
  wire [0:0] cby_1__1__48_left_grid_pin_19_;
  wire [0:0] cby_1__1__48_left_grid_pin_20_;
  wire [0:0] cby_1__1__48_left_grid_pin_21_;
  wire [0:0] cby_1__1__48_left_grid_pin_22_;
  wire [0:0] cby_1__1__48_left_grid_pin_23_;
  wire [0:0] cby_1__1__48_left_grid_pin_24_;
  wire [0:0] cby_1__1__48_left_grid_pin_25_;
  wire [0:0] cby_1__1__48_left_grid_pin_26_;
  wire [0:0] cby_1__1__48_left_grid_pin_27_;
  wire [0:0] cby_1__1__48_left_grid_pin_28_;
  wire [0:0] cby_1__1__48_left_grid_pin_29_;
  wire [0:0] cby_1__1__48_left_grid_pin_30_;
  wire [0:0] cby_1__1__48_left_grid_pin_31_;
  wire [0:0] cby_1__1__49_ccff_tail;
  wire [0:19] cby_1__1__49_chany_bottom_out;
  wire [0:19] cby_1__1__49_chany_top_out;
  wire [0:0] cby_1__1__49_left_grid_pin_16_;
  wire [0:0] cby_1__1__49_left_grid_pin_17_;
  wire [0:0] cby_1__1__49_left_grid_pin_18_;
  wire [0:0] cby_1__1__49_left_grid_pin_19_;
  wire [0:0] cby_1__1__49_left_grid_pin_20_;
  wire [0:0] cby_1__1__49_left_grid_pin_21_;
  wire [0:0] cby_1__1__49_left_grid_pin_22_;
  wire [0:0] cby_1__1__49_left_grid_pin_23_;
  wire [0:0] cby_1__1__49_left_grid_pin_24_;
  wire [0:0] cby_1__1__49_left_grid_pin_25_;
  wire [0:0] cby_1__1__49_left_grid_pin_26_;
  wire [0:0] cby_1__1__49_left_grid_pin_27_;
  wire [0:0] cby_1__1__49_left_grid_pin_28_;
  wire [0:0] cby_1__1__49_left_grid_pin_29_;
  wire [0:0] cby_1__1__49_left_grid_pin_30_;
  wire [0:0] cby_1__1__49_left_grid_pin_31_;
  wire [0:0] cby_1__1__4_ccff_tail;
  wire [0:19] cby_1__1__4_chany_bottom_out;
  wire [0:19] cby_1__1__4_chany_top_out;
  wire [0:0] cby_1__1__4_left_grid_pin_16_;
  wire [0:0] cby_1__1__4_left_grid_pin_17_;
  wire [0:0] cby_1__1__4_left_grid_pin_18_;
  wire [0:0] cby_1__1__4_left_grid_pin_19_;
  wire [0:0] cby_1__1__4_left_grid_pin_20_;
  wire [0:0] cby_1__1__4_left_grid_pin_21_;
  wire [0:0] cby_1__1__4_left_grid_pin_22_;
  wire [0:0] cby_1__1__4_left_grid_pin_23_;
  wire [0:0] cby_1__1__4_left_grid_pin_24_;
  wire [0:0] cby_1__1__4_left_grid_pin_25_;
  wire [0:0] cby_1__1__4_left_grid_pin_26_;
  wire [0:0] cby_1__1__4_left_grid_pin_27_;
  wire [0:0] cby_1__1__4_left_grid_pin_28_;
  wire [0:0] cby_1__1__4_left_grid_pin_29_;
  wire [0:0] cby_1__1__4_left_grid_pin_30_;
  wire [0:0] cby_1__1__4_left_grid_pin_31_;
  wire [0:0] cby_1__1__50_ccff_tail;
  wire [0:19] cby_1__1__50_chany_bottom_out;
  wire [0:19] cby_1__1__50_chany_top_out;
  wire [0:0] cby_1__1__50_left_grid_pin_16_;
  wire [0:0] cby_1__1__50_left_grid_pin_17_;
  wire [0:0] cby_1__1__50_left_grid_pin_18_;
  wire [0:0] cby_1__1__50_left_grid_pin_19_;
  wire [0:0] cby_1__1__50_left_grid_pin_20_;
  wire [0:0] cby_1__1__50_left_grid_pin_21_;
  wire [0:0] cby_1__1__50_left_grid_pin_22_;
  wire [0:0] cby_1__1__50_left_grid_pin_23_;
  wire [0:0] cby_1__1__50_left_grid_pin_24_;
  wire [0:0] cby_1__1__50_left_grid_pin_25_;
  wire [0:0] cby_1__1__50_left_grid_pin_26_;
  wire [0:0] cby_1__1__50_left_grid_pin_27_;
  wire [0:0] cby_1__1__50_left_grid_pin_28_;
  wire [0:0] cby_1__1__50_left_grid_pin_29_;
  wire [0:0] cby_1__1__50_left_grid_pin_30_;
  wire [0:0] cby_1__1__50_left_grid_pin_31_;
  wire [0:0] cby_1__1__51_ccff_tail;
  wire [0:19] cby_1__1__51_chany_bottom_out;
  wire [0:19] cby_1__1__51_chany_top_out;
  wire [0:0] cby_1__1__51_left_grid_pin_16_;
  wire [0:0] cby_1__1__51_left_grid_pin_17_;
  wire [0:0] cby_1__1__51_left_grid_pin_18_;
  wire [0:0] cby_1__1__51_left_grid_pin_19_;
  wire [0:0] cby_1__1__51_left_grid_pin_20_;
  wire [0:0] cby_1__1__51_left_grid_pin_21_;
  wire [0:0] cby_1__1__51_left_grid_pin_22_;
  wire [0:0] cby_1__1__51_left_grid_pin_23_;
  wire [0:0] cby_1__1__51_left_grid_pin_24_;
  wire [0:0] cby_1__1__51_left_grid_pin_25_;
  wire [0:0] cby_1__1__51_left_grid_pin_26_;
  wire [0:0] cby_1__1__51_left_grid_pin_27_;
  wire [0:0] cby_1__1__51_left_grid_pin_28_;
  wire [0:0] cby_1__1__51_left_grid_pin_29_;
  wire [0:0] cby_1__1__51_left_grid_pin_30_;
  wire [0:0] cby_1__1__51_left_grid_pin_31_;
  wire [0:0] cby_1__1__52_ccff_tail;
  wire [0:19] cby_1__1__52_chany_bottom_out;
  wire [0:19] cby_1__1__52_chany_top_out;
  wire [0:0] cby_1__1__52_left_grid_pin_16_;
  wire [0:0] cby_1__1__52_left_grid_pin_17_;
  wire [0:0] cby_1__1__52_left_grid_pin_18_;
  wire [0:0] cby_1__1__52_left_grid_pin_19_;
  wire [0:0] cby_1__1__52_left_grid_pin_20_;
  wire [0:0] cby_1__1__52_left_grid_pin_21_;
  wire [0:0] cby_1__1__52_left_grid_pin_22_;
  wire [0:0] cby_1__1__52_left_grid_pin_23_;
  wire [0:0] cby_1__1__52_left_grid_pin_24_;
  wire [0:0] cby_1__1__52_left_grid_pin_25_;
  wire [0:0] cby_1__1__52_left_grid_pin_26_;
  wire [0:0] cby_1__1__52_left_grid_pin_27_;
  wire [0:0] cby_1__1__52_left_grid_pin_28_;
  wire [0:0] cby_1__1__52_left_grid_pin_29_;
  wire [0:0] cby_1__1__52_left_grid_pin_30_;
  wire [0:0] cby_1__1__52_left_grid_pin_31_;
  wire [0:0] cby_1__1__53_ccff_tail;
  wire [0:19] cby_1__1__53_chany_bottom_out;
  wire [0:19] cby_1__1__53_chany_top_out;
  wire [0:0] cby_1__1__53_left_grid_pin_16_;
  wire [0:0] cby_1__1__53_left_grid_pin_17_;
  wire [0:0] cby_1__1__53_left_grid_pin_18_;
  wire [0:0] cby_1__1__53_left_grid_pin_19_;
  wire [0:0] cby_1__1__53_left_grid_pin_20_;
  wire [0:0] cby_1__1__53_left_grid_pin_21_;
  wire [0:0] cby_1__1__53_left_grid_pin_22_;
  wire [0:0] cby_1__1__53_left_grid_pin_23_;
  wire [0:0] cby_1__1__53_left_grid_pin_24_;
  wire [0:0] cby_1__1__53_left_grid_pin_25_;
  wire [0:0] cby_1__1__53_left_grid_pin_26_;
  wire [0:0] cby_1__1__53_left_grid_pin_27_;
  wire [0:0] cby_1__1__53_left_grid_pin_28_;
  wire [0:0] cby_1__1__53_left_grid_pin_29_;
  wire [0:0] cby_1__1__53_left_grid_pin_30_;
  wire [0:0] cby_1__1__53_left_grid_pin_31_;
  wire [0:0] cby_1__1__54_ccff_tail;
  wire [0:19] cby_1__1__54_chany_bottom_out;
  wire [0:19] cby_1__1__54_chany_top_out;
  wire [0:0] cby_1__1__54_left_grid_pin_16_;
  wire [0:0] cby_1__1__54_left_grid_pin_17_;
  wire [0:0] cby_1__1__54_left_grid_pin_18_;
  wire [0:0] cby_1__1__54_left_grid_pin_19_;
  wire [0:0] cby_1__1__54_left_grid_pin_20_;
  wire [0:0] cby_1__1__54_left_grid_pin_21_;
  wire [0:0] cby_1__1__54_left_grid_pin_22_;
  wire [0:0] cby_1__1__54_left_grid_pin_23_;
  wire [0:0] cby_1__1__54_left_grid_pin_24_;
  wire [0:0] cby_1__1__54_left_grid_pin_25_;
  wire [0:0] cby_1__1__54_left_grid_pin_26_;
  wire [0:0] cby_1__1__54_left_grid_pin_27_;
  wire [0:0] cby_1__1__54_left_grid_pin_28_;
  wire [0:0] cby_1__1__54_left_grid_pin_29_;
  wire [0:0] cby_1__1__54_left_grid_pin_30_;
  wire [0:0] cby_1__1__54_left_grid_pin_31_;
  wire [0:0] cby_1__1__55_ccff_tail;
  wire [0:19] cby_1__1__55_chany_bottom_out;
  wire [0:19] cby_1__1__55_chany_top_out;
  wire [0:0] cby_1__1__55_left_grid_pin_16_;
  wire [0:0] cby_1__1__55_left_grid_pin_17_;
  wire [0:0] cby_1__1__55_left_grid_pin_18_;
  wire [0:0] cby_1__1__55_left_grid_pin_19_;
  wire [0:0] cby_1__1__55_left_grid_pin_20_;
  wire [0:0] cby_1__1__55_left_grid_pin_21_;
  wire [0:0] cby_1__1__55_left_grid_pin_22_;
  wire [0:0] cby_1__1__55_left_grid_pin_23_;
  wire [0:0] cby_1__1__55_left_grid_pin_24_;
  wire [0:0] cby_1__1__55_left_grid_pin_25_;
  wire [0:0] cby_1__1__55_left_grid_pin_26_;
  wire [0:0] cby_1__1__55_left_grid_pin_27_;
  wire [0:0] cby_1__1__55_left_grid_pin_28_;
  wire [0:0] cby_1__1__55_left_grid_pin_29_;
  wire [0:0] cby_1__1__55_left_grid_pin_30_;
  wire [0:0] cby_1__1__55_left_grid_pin_31_;
  wire [0:0] cby_1__1__56_ccff_tail;
  wire [0:19] cby_1__1__56_chany_bottom_out;
  wire [0:19] cby_1__1__56_chany_top_out;
  wire [0:0] cby_1__1__56_left_grid_pin_16_;
  wire [0:0] cby_1__1__56_left_grid_pin_17_;
  wire [0:0] cby_1__1__56_left_grid_pin_18_;
  wire [0:0] cby_1__1__56_left_grid_pin_19_;
  wire [0:0] cby_1__1__56_left_grid_pin_20_;
  wire [0:0] cby_1__1__56_left_grid_pin_21_;
  wire [0:0] cby_1__1__56_left_grid_pin_22_;
  wire [0:0] cby_1__1__56_left_grid_pin_23_;
  wire [0:0] cby_1__1__56_left_grid_pin_24_;
  wire [0:0] cby_1__1__56_left_grid_pin_25_;
  wire [0:0] cby_1__1__56_left_grid_pin_26_;
  wire [0:0] cby_1__1__56_left_grid_pin_27_;
  wire [0:0] cby_1__1__56_left_grid_pin_28_;
  wire [0:0] cby_1__1__56_left_grid_pin_29_;
  wire [0:0] cby_1__1__56_left_grid_pin_30_;
  wire [0:0] cby_1__1__56_left_grid_pin_31_;
  wire [0:0] cby_1__1__57_ccff_tail;
  wire [0:19] cby_1__1__57_chany_bottom_out;
  wire [0:19] cby_1__1__57_chany_top_out;
  wire [0:0] cby_1__1__57_left_grid_pin_16_;
  wire [0:0] cby_1__1__57_left_grid_pin_17_;
  wire [0:0] cby_1__1__57_left_grid_pin_18_;
  wire [0:0] cby_1__1__57_left_grid_pin_19_;
  wire [0:0] cby_1__1__57_left_grid_pin_20_;
  wire [0:0] cby_1__1__57_left_grid_pin_21_;
  wire [0:0] cby_1__1__57_left_grid_pin_22_;
  wire [0:0] cby_1__1__57_left_grid_pin_23_;
  wire [0:0] cby_1__1__57_left_grid_pin_24_;
  wire [0:0] cby_1__1__57_left_grid_pin_25_;
  wire [0:0] cby_1__1__57_left_grid_pin_26_;
  wire [0:0] cby_1__1__57_left_grid_pin_27_;
  wire [0:0] cby_1__1__57_left_grid_pin_28_;
  wire [0:0] cby_1__1__57_left_grid_pin_29_;
  wire [0:0] cby_1__1__57_left_grid_pin_30_;
  wire [0:0] cby_1__1__57_left_grid_pin_31_;
  wire [0:0] cby_1__1__58_ccff_tail;
  wire [0:19] cby_1__1__58_chany_bottom_out;
  wire [0:19] cby_1__1__58_chany_top_out;
  wire [0:0] cby_1__1__58_left_grid_pin_16_;
  wire [0:0] cby_1__1__58_left_grid_pin_17_;
  wire [0:0] cby_1__1__58_left_grid_pin_18_;
  wire [0:0] cby_1__1__58_left_grid_pin_19_;
  wire [0:0] cby_1__1__58_left_grid_pin_20_;
  wire [0:0] cby_1__1__58_left_grid_pin_21_;
  wire [0:0] cby_1__1__58_left_grid_pin_22_;
  wire [0:0] cby_1__1__58_left_grid_pin_23_;
  wire [0:0] cby_1__1__58_left_grid_pin_24_;
  wire [0:0] cby_1__1__58_left_grid_pin_25_;
  wire [0:0] cby_1__1__58_left_grid_pin_26_;
  wire [0:0] cby_1__1__58_left_grid_pin_27_;
  wire [0:0] cby_1__1__58_left_grid_pin_28_;
  wire [0:0] cby_1__1__58_left_grid_pin_29_;
  wire [0:0] cby_1__1__58_left_grid_pin_30_;
  wire [0:0] cby_1__1__58_left_grid_pin_31_;
  wire [0:0] cby_1__1__59_ccff_tail;
  wire [0:19] cby_1__1__59_chany_bottom_out;
  wire [0:19] cby_1__1__59_chany_top_out;
  wire [0:0] cby_1__1__59_left_grid_pin_16_;
  wire [0:0] cby_1__1__59_left_grid_pin_17_;
  wire [0:0] cby_1__1__59_left_grid_pin_18_;
  wire [0:0] cby_1__1__59_left_grid_pin_19_;
  wire [0:0] cby_1__1__59_left_grid_pin_20_;
  wire [0:0] cby_1__1__59_left_grid_pin_21_;
  wire [0:0] cby_1__1__59_left_grid_pin_22_;
  wire [0:0] cby_1__1__59_left_grid_pin_23_;
  wire [0:0] cby_1__1__59_left_grid_pin_24_;
  wire [0:0] cby_1__1__59_left_grid_pin_25_;
  wire [0:0] cby_1__1__59_left_grid_pin_26_;
  wire [0:0] cby_1__1__59_left_grid_pin_27_;
  wire [0:0] cby_1__1__59_left_grid_pin_28_;
  wire [0:0] cby_1__1__59_left_grid_pin_29_;
  wire [0:0] cby_1__1__59_left_grid_pin_30_;
  wire [0:0] cby_1__1__59_left_grid_pin_31_;
  wire [0:0] cby_1__1__5_ccff_tail;
  wire [0:19] cby_1__1__5_chany_bottom_out;
  wire [0:19] cby_1__1__5_chany_top_out;
  wire [0:0] cby_1__1__5_left_grid_pin_16_;
  wire [0:0] cby_1__1__5_left_grid_pin_17_;
  wire [0:0] cby_1__1__5_left_grid_pin_18_;
  wire [0:0] cby_1__1__5_left_grid_pin_19_;
  wire [0:0] cby_1__1__5_left_grid_pin_20_;
  wire [0:0] cby_1__1__5_left_grid_pin_21_;
  wire [0:0] cby_1__1__5_left_grid_pin_22_;
  wire [0:0] cby_1__1__5_left_grid_pin_23_;
  wire [0:0] cby_1__1__5_left_grid_pin_24_;
  wire [0:0] cby_1__1__5_left_grid_pin_25_;
  wire [0:0] cby_1__1__5_left_grid_pin_26_;
  wire [0:0] cby_1__1__5_left_grid_pin_27_;
  wire [0:0] cby_1__1__5_left_grid_pin_28_;
  wire [0:0] cby_1__1__5_left_grid_pin_29_;
  wire [0:0] cby_1__1__5_left_grid_pin_30_;
  wire [0:0] cby_1__1__5_left_grid_pin_31_;
  wire [0:0] cby_1__1__60_ccff_tail;
  wire [0:19] cby_1__1__60_chany_bottom_out;
  wire [0:19] cby_1__1__60_chany_top_out;
  wire [0:0] cby_1__1__60_left_grid_pin_16_;
  wire [0:0] cby_1__1__60_left_grid_pin_17_;
  wire [0:0] cby_1__1__60_left_grid_pin_18_;
  wire [0:0] cby_1__1__60_left_grid_pin_19_;
  wire [0:0] cby_1__1__60_left_grid_pin_20_;
  wire [0:0] cby_1__1__60_left_grid_pin_21_;
  wire [0:0] cby_1__1__60_left_grid_pin_22_;
  wire [0:0] cby_1__1__60_left_grid_pin_23_;
  wire [0:0] cby_1__1__60_left_grid_pin_24_;
  wire [0:0] cby_1__1__60_left_grid_pin_25_;
  wire [0:0] cby_1__1__60_left_grid_pin_26_;
  wire [0:0] cby_1__1__60_left_grid_pin_27_;
  wire [0:0] cby_1__1__60_left_grid_pin_28_;
  wire [0:0] cby_1__1__60_left_grid_pin_29_;
  wire [0:0] cby_1__1__60_left_grid_pin_30_;
  wire [0:0] cby_1__1__60_left_grid_pin_31_;
  wire [0:0] cby_1__1__61_ccff_tail;
  wire [0:19] cby_1__1__61_chany_bottom_out;
  wire [0:19] cby_1__1__61_chany_top_out;
  wire [0:0] cby_1__1__61_left_grid_pin_16_;
  wire [0:0] cby_1__1__61_left_grid_pin_17_;
  wire [0:0] cby_1__1__61_left_grid_pin_18_;
  wire [0:0] cby_1__1__61_left_grid_pin_19_;
  wire [0:0] cby_1__1__61_left_grid_pin_20_;
  wire [0:0] cby_1__1__61_left_grid_pin_21_;
  wire [0:0] cby_1__1__61_left_grid_pin_22_;
  wire [0:0] cby_1__1__61_left_grid_pin_23_;
  wire [0:0] cby_1__1__61_left_grid_pin_24_;
  wire [0:0] cby_1__1__61_left_grid_pin_25_;
  wire [0:0] cby_1__1__61_left_grid_pin_26_;
  wire [0:0] cby_1__1__61_left_grid_pin_27_;
  wire [0:0] cby_1__1__61_left_grid_pin_28_;
  wire [0:0] cby_1__1__61_left_grid_pin_29_;
  wire [0:0] cby_1__1__61_left_grid_pin_30_;
  wire [0:0] cby_1__1__61_left_grid_pin_31_;
  wire [0:0] cby_1__1__62_ccff_tail;
  wire [0:19] cby_1__1__62_chany_bottom_out;
  wire [0:19] cby_1__1__62_chany_top_out;
  wire [0:0] cby_1__1__62_left_grid_pin_16_;
  wire [0:0] cby_1__1__62_left_grid_pin_17_;
  wire [0:0] cby_1__1__62_left_grid_pin_18_;
  wire [0:0] cby_1__1__62_left_grid_pin_19_;
  wire [0:0] cby_1__1__62_left_grid_pin_20_;
  wire [0:0] cby_1__1__62_left_grid_pin_21_;
  wire [0:0] cby_1__1__62_left_grid_pin_22_;
  wire [0:0] cby_1__1__62_left_grid_pin_23_;
  wire [0:0] cby_1__1__62_left_grid_pin_24_;
  wire [0:0] cby_1__1__62_left_grid_pin_25_;
  wire [0:0] cby_1__1__62_left_grid_pin_26_;
  wire [0:0] cby_1__1__62_left_grid_pin_27_;
  wire [0:0] cby_1__1__62_left_grid_pin_28_;
  wire [0:0] cby_1__1__62_left_grid_pin_29_;
  wire [0:0] cby_1__1__62_left_grid_pin_30_;
  wire [0:0] cby_1__1__62_left_grid_pin_31_;
  wire [0:0] cby_1__1__63_ccff_tail;
  wire [0:19] cby_1__1__63_chany_bottom_out;
  wire [0:19] cby_1__1__63_chany_top_out;
  wire [0:0] cby_1__1__63_left_grid_pin_16_;
  wire [0:0] cby_1__1__63_left_grid_pin_17_;
  wire [0:0] cby_1__1__63_left_grid_pin_18_;
  wire [0:0] cby_1__1__63_left_grid_pin_19_;
  wire [0:0] cby_1__1__63_left_grid_pin_20_;
  wire [0:0] cby_1__1__63_left_grid_pin_21_;
  wire [0:0] cby_1__1__63_left_grid_pin_22_;
  wire [0:0] cby_1__1__63_left_grid_pin_23_;
  wire [0:0] cby_1__1__63_left_grid_pin_24_;
  wire [0:0] cby_1__1__63_left_grid_pin_25_;
  wire [0:0] cby_1__1__63_left_grid_pin_26_;
  wire [0:0] cby_1__1__63_left_grid_pin_27_;
  wire [0:0] cby_1__1__63_left_grid_pin_28_;
  wire [0:0] cby_1__1__63_left_grid_pin_29_;
  wire [0:0] cby_1__1__63_left_grid_pin_30_;
  wire [0:0] cby_1__1__63_left_grid_pin_31_;
  wire [0:0] cby_1__1__64_ccff_tail;
  wire [0:19] cby_1__1__64_chany_bottom_out;
  wire [0:19] cby_1__1__64_chany_top_out;
  wire [0:0] cby_1__1__64_left_grid_pin_16_;
  wire [0:0] cby_1__1__64_left_grid_pin_17_;
  wire [0:0] cby_1__1__64_left_grid_pin_18_;
  wire [0:0] cby_1__1__64_left_grid_pin_19_;
  wire [0:0] cby_1__1__64_left_grid_pin_20_;
  wire [0:0] cby_1__1__64_left_grid_pin_21_;
  wire [0:0] cby_1__1__64_left_grid_pin_22_;
  wire [0:0] cby_1__1__64_left_grid_pin_23_;
  wire [0:0] cby_1__1__64_left_grid_pin_24_;
  wire [0:0] cby_1__1__64_left_grid_pin_25_;
  wire [0:0] cby_1__1__64_left_grid_pin_26_;
  wire [0:0] cby_1__1__64_left_grid_pin_27_;
  wire [0:0] cby_1__1__64_left_grid_pin_28_;
  wire [0:0] cby_1__1__64_left_grid_pin_29_;
  wire [0:0] cby_1__1__64_left_grid_pin_30_;
  wire [0:0] cby_1__1__64_left_grid_pin_31_;
  wire [0:0] cby_1__1__65_ccff_tail;
  wire [0:19] cby_1__1__65_chany_bottom_out;
  wire [0:19] cby_1__1__65_chany_top_out;
  wire [0:0] cby_1__1__65_left_grid_pin_16_;
  wire [0:0] cby_1__1__65_left_grid_pin_17_;
  wire [0:0] cby_1__1__65_left_grid_pin_18_;
  wire [0:0] cby_1__1__65_left_grid_pin_19_;
  wire [0:0] cby_1__1__65_left_grid_pin_20_;
  wire [0:0] cby_1__1__65_left_grid_pin_21_;
  wire [0:0] cby_1__1__65_left_grid_pin_22_;
  wire [0:0] cby_1__1__65_left_grid_pin_23_;
  wire [0:0] cby_1__1__65_left_grid_pin_24_;
  wire [0:0] cby_1__1__65_left_grid_pin_25_;
  wire [0:0] cby_1__1__65_left_grid_pin_26_;
  wire [0:0] cby_1__1__65_left_grid_pin_27_;
  wire [0:0] cby_1__1__65_left_grid_pin_28_;
  wire [0:0] cby_1__1__65_left_grid_pin_29_;
  wire [0:0] cby_1__1__65_left_grid_pin_30_;
  wire [0:0] cby_1__1__65_left_grid_pin_31_;
  wire [0:0] cby_1__1__66_ccff_tail;
  wire [0:19] cby_1__1__66_chany_bottom_out;
  wire [0:19] cby_1__1__66_chany_top_out;
  wire [0:0] cby_1__1__66_left_grid_pin_16_;
  wire [0:0] cby_1__1__66_left_grid_pin_17_;
  wire [0:0] cby_1__1__66_left_grid_pin_18_;
  wire [0:0] cby_1__1__66_left_grid_pin_19_;
  wire [0:0] cby_1__1__66_left_grid_pin_20_;
  wire [0:0] cby_1__1__66_left_grid_pin_21_;
  wire [0:0] cby_1__1__66_left_grid_pin_22_;
  wire [0:0] cby_1__1__66_left_grid_pin_23_;
  wire [0:0] cby_1__1__66_left_grid_pin_24_;
  wire [0:0] cby_1__1__66_left_grid_pin_25_;
  wire [0:0] cby_1__1__66_left_grid_pin_26_;
  wire [0:0] cby_1__1__66_left_grid_pin_27_;
  wire [0:0] cby_1__1__66_left_grid_pin_28_;
  wire [0:0] cby_1__1__66_left_grid_pin_29_;
  wire [0:0] cby_1__1__66_left_grid_pin_30_;
  wire [0:0] cby_1__1__66_left_grid_pin_31_;
  wire [0:0] cby_1__1__67_ccff_tail;
  wire [0:19] cby_1__1__67_chany_bottom_out;
  wire [0:19] cby_1__1__67_chany_top_out;
  wire [0:0] cby_1__1__67_left_grid_pin_16_;
  wire [0:0] cby_1__1__67_left_grid_pin_17_;
  wire [0:0] cby_1__1__67_left_grid_pin_18_;
  wire [0:0] cby_1__1__67_left_grid_pin_19_;
  wire [0:0] cby_1__1__67_left_grid_pin_20_;
  wire [0:0] cby_1__1__67_left_grid_pin_21_;
  wire [0:0] cby_1__1__67_left_grid_pin_22_;
  wire [0:0] cby_1__1__67_left_grid_pin_23_;
  wire [0:0] cby_1__1__67_left_grid_pin_24_;
  wire [0:0] cby_1__1__67_left_grid_pin_25_;
  wire [0:0] cby_1__1__67_left_grid_pin_26_;
  wire [0:0] cby_1__1__67_left_grid_pin_27_;
  wire [0:0] cby_1__1__67_left_grid_pin_28_;
  wire [0:0] cby_1__1__67_left_grid_pin_29_;
  wire [0:0] cby_1__1__67_left_grid_pin_30_;
  wire [0:0] cby_1__1__67_left_grid_pin_31_;
  wire [0:0] cby_1__1__68_ccff_tail;
  wire [0:19] cby_1__1__68_chany_bottom_out;
  wire [0:19] cby_1__1__68_chany_top_out;
  wire [0:0] cby_1__1__68_left_grid_pin_16_;
  wire [0:0] cby_1__1__68_left_grid_pin_17_;
  wire [0:0] cby_1__1__68_left_grid_pin_18_;
  wire [0:0] cby_1__1__68_left_grid_pin_19_;
  wire [0:0] cby_1__1__68_left_grid_pin_20_;
  wire [0:0] cby_1__1__68_left_grid_pin_21_;
  wire [0:0] cby_1__1__68_left_grid_pin_22_;
  wire [0:0] cby_1__1__68_left_grid_pin_23_;
  wire [0:0] cby_1__1__68_left_grid_pin_24_;
  wire [0:0] cby_1__1__68_left_grid_pin_25_;
  wire [0:0] cby_1__1__68_left_grid_pin_26_;
  wire [0:0] cby_1__1__68_left_grid_pin_27_;
  wire [0:0] cby_1__1__68_left_grid_pin_28_;
  wire [0:0] cby_1__1__68_left_grid_pin_29_;
  wire [0:0] cby_1__1__68_left_grid_pin_30_;
  wire [0:0] cby_1__1__68_left_grid_pin_31_;
  wire [0:0] cby_1__1__69_ccff_tail;
  wire [0:19] cby_1__1__69_chany_bottom_out;
  wire [0:19] cby_1__1__69_chany_top_out;
  wire [0:0] cby_1__1__69_left_grid_pin_16_;
  wire [0:0] cby_1__1__69_left_grid_pin_17_;
  wire [0:0] cby_1__1__69_left_grid_pin_18_;
  wire [0:0] cby_1__1__69_left_grid_pin_19_;
  wire [0:0] cby_1__1__69_left_grid_pin_20_;
  wire [0:0] cby_1__1__69_left_grid_pin_21_;
  wire [0:0] cby_1__1__69_left_grid_pin_22_;
  wire [0:0] cby_1__1__69_left_grid_pin_23_;
  wire [0:0] cby_1__1__69_left_grid_pin_24_;
  wire [0:0] cby_1__1__69_left_grid_pin_25_;
  wire [0:0] cby_1__1__69_left_grid_pin_26_;
  wire [0:0] cby_1__1__69_left_grid_pin_27_;
  wire [0:0] cby_1__1__69_left_grid_pin_28_;
  wire [0:0] cby_1__1__69_left_grid_pin_29_;
  wire [0:0] cby_1__1__69_left_grid_pin_30_;
  wire [0:0] cby_1__1__69_left_grid_pin_31_;
  wire [0:0] cby_1__1__6_ccff_tail;
  wire [0:19] cby_1__1__6_chany_bottom_out;
  wire [0:19] cby_1__1__6_chany_top_out;
  wire [0:0] cby_1__1__6_left_grid_pin_16_;
  wire [0:0] cby_1__1__6_left_grid_pin_17_;
  wire [0:0] cby_1__1__6_left_grid_pin_18_;
  wire [0:0] cby_1__1__6_left_grid_pin_19_;
  wire [0:0] cby_1__1__6_left_grid_pin_20_;
  wire [0:0] cby_1__1__6_left_grid_pin_21_;
  wire [0:0] cby_1__1__6_left_grid_pin_22_;
  wire [0:0] cby_1__1__6_left_grid_pin_23_;
  wire [0:0] cby_1__1__6_left_grid_pin_24_;
  wire [0:0] cby_1__1__6_left_grid_pin_25_;
  wire [0:0] cby_1__1__6_left_grid_pin_26_;
  wire [0:0] cby_1__1__6_left_grid_pin_27_;
  wire [0:0] cby_1__1__6_left_grid_pin_28_;
  wire [0:0] cby_1__1__6_left_grid_pin_29_;
  wire [0:0] cby_1__1__6_left_grid_pin_30_;
  wire [0:0] cby_1__1__6_left_grid_pin_31_;
  wire [0:0] cby_1__1__70_ccff_tail;
  wire [0:19] cby_1__1__70_chany_bottom_out;
  wire [0:19] cby_1__1__70_chany_top_out;
  wire [0:0] cby_1__1__70_left_grid_pin_16_;
  wire [0:0] cby_1__1__70_left_grid_pin_17_;
  wire [0:0] cby_1__1__70_left_grid_pin_18_;
  wire [0:0] cby_1__1__70_left_grid_pin_19_;
  wire [0:0] cby_1__1__70_left_grid_pin_20_;
  wire [0:0] cby_1__1__70_left_grid_pin_21_;
  wire [0:0] cby_1__1__70_left_grid_pin_22_;
  wire [0:0] cby_1__1__70_left_grid_pin_23_;
  wire [0:0] cby_1__1__70_left_grid_pin_24_;
  wire [0:0] cby_1__1__70_left_grid_pin_25_;
  wire [0:0] cby_1__1__70_left_grid_pin_26_;
  wire [0:0] cby_1__1__70_left_grid_pin_27_;
  wire [0:0] cby_1__1__70_left_grid_pin_28_;
  wire [0:0] cby_1__1__70_left_grid_pin_29_;
  wire [0:0] cby_1__1__70_left_grid_pin_30_;
  wire [0:0] cby_1__1__70_left_grid_pin_31_;
  wire [0:0] cby_1__1__71_ccff_tail;
  wire [0:19] cby_1__1__71_chany_bottom_out;
  wire [0:19] cby_1__1__71_chany_top_out;
  wire [0:0] cby_1__1__71_left_grid_pin_16_;
  wire [0:0] cby_1__1__71_left_grid_pin_17_;
  wire [0:0] cby_1__1__71_left_grid_pin_18_;
  wire [0:0] cby_1__1__71_left_grid_pin_19_;
  wire [0:0] cby_1__1__71_left_grid_pin_20_;
  wire [0:0] cby_1__1__71_left_grid_pin_21_;
  wire [0:0] cby_1__1__71_left_grid_pin_22_;
  wire [0:0] cby_1__1__71_left_grid_pin_23_;
  wire [0:0] cby_1__1__71_left_grid_pin_24_;
  wire [0:0] cby_1__1__71_left_grid_pin_25_;
  wire [0:0] cby_1__1__71_left_grid_pin_26_;
  wire [0:0] cby_1__1__71_left_grid_pin_27_;
  wire [0:0] cby_1__1__71_left_grid_pin_28_;
  wire [0:0] cby_1__1__71_left_grid_pin_29_;
  wire [0:0] cby_1__1__71_left_grid_pin_30_;
  wire [0:0] cby_1__1__71_left_grid_pin_31_;
  wire [0:0] cby_1__1__72_ccff_tail;
  wire [0:19] cby_1__1__72_chany_bottom_out;
  wire [0:19] cby_1__1__72_chany_top_out;
  wire [0:0] cby_1__1__72_left_grid_pin_16_;
  wire [0:0] cby_1__1__72_left_grid_pin_17_;
  wire [0:0] cby_1__1__72_left_grid_pin_18_;
  wire [0:0] cby_1__1__72_left_grid_pin_19_;
  wire [0:0] cby_1__1__72_left_grid_pin_20_;
  wire [0:0] cby_1__1__72_left_grid_pin_21_;
  wire [0:0] cby_1__1__72_left_grid_pin_22_;
  wire [0:0] cby_1__1__72_left_grid_pin_23_;
  wire [0:0] cby_1__1__72_left_grid_pin_24_;
  wire [0:0] cby_1__1__72_left_grid_pin_25_;
  wire [0:0] cby_1__1__72_left_grid_pin_26_;
  wire [0:0] cby_1__1__72_left_grid_pin_27_;
  wire [0:0] cby_1__1__72_left_grid_pin_28_;
  wire [0:0] cby_1__1__72_left_grid_pin_29_;
  wire [0:0] cby_1__1__72_left_grid_pin_30_;
  wire [0:0] cby_1__1__72_left_grid_pin_31_;
  wire [0:0] cby_1__1__73_ccff_tail;
  wire [0:19] cby_1__1__73_chany_bottom_out;
  wire [0:19] cby_1__1__73_chany_top_out;
  wire [0:0] cby_1__1__73_left_grid_pin_16_;
  wire [0:0] cby_1__1__73_left_grid_pin_17_;
  wire [0:0] cby_1__1__73_left_grid_pin_18_;
  wire [0:0] cby_1__1__73_left_grid_pin_19_;
  wire [0:0] cby_1__1__73_left_grid_pin_20_;
  wire [0:0] cby_1__1__73_left_grid_pin_21_;
  wire [0:0] cby_1__1__73_left_grid_pin_22_;
  wire [0:0] cby_1__1__73_left_grid_pin_23_;
  wire [0:0] cby_1__1__73_left_grid_pin_24_;
  wire [0:0] cby_1__1__73_left_grid_pin_25_;
  wire [0:0] cby_1__1__73_left_grid_pin_26_;
  wire [0:0] cby_1__1__73_left_grid_pin_27_;
  wire [0:0] cby_1__1__73_left_grid_pin_28_;
  wire [0:0] cby_1__1__73_left_grid_pin_29_;
  wire [0:0] cby_1__1__73_left_grid_pin_30_;
  wire [0:0] cby_1__1__73_left_grid_pin_31_;
  wire [0:0] cby_1__1__74_ccff_tail;
  wire [0:19] cby_1__1__74_chany_bottom_out;
  wire [0:19] cby_1__1__74_chany_top_out;
  wire [0:0] cby_1__1__74_left_grid_pin_16_;
  wire [0:0] cby_1__1__74_left_grid_pin_17_;
  wire [0:0] cby_1__1__74_left_grid_pin_18_;
  wire [0:0] cby_1__1__74_left_grid_pin_19_;
  wire [0:0] cby_1__1__74_left_grid_pin_20_;
  wire [0:0] cby_1__1__74_left_grid_pin_21_;
  wire [0:0] cby_1__1__74_left_grid_pin_22_;
  wire [0:0] cby_1__1__74_left_grid_pin_23_;
  wire [0:0] cby_1__1__74_left_grid_pin_24_;
  wire [0:0] cby_1__1__74_left_grid_pin_25_;
  wire [0:0] cby_1__1__74_left_grid_pin_26_;
  wire [0:0] cby_1__1__74_left_grid_pin_27_;
  wire [0:0] cby_1__1__74_left_grid_pin_28_;
  wire [0:0] cby_1__1__74_left_grid_pin_29_;
  wire [0:0] cby_1__1__74_left_grid_pin_30_;
  wire [0:0] cby_1__1__74_left_grid_pin_31_;
  wire [0:0] cby_1__1__75_ccff_tail;
  wire [0:19] cby_1__1__75_chany_bottom_out;
  wire [0:19] cby_1__1__75_chany_top_out;
  wire [0:0] cby_1__1__75_left_grid_pin_16_;
  wire [0:0] cby_1__1__75_left_grid_pin_17_;
  wire [0:0] cby_1__1__75_left_grid_pin_18_;
  wire [0:0] cby_1__1__75_left_grid_pin_19_;
  wire [0:0] cby_1__1__75_left_grid_pin_20_;
  wire [0:0] cby_1__1__75_left_grid_pin_21_;
  wire [0:0] cby_1__1__75_left_grid_pin_22_;
  wire [0:0] cby_1__1__75_left_grid_pin_23_;
  wire [0:0] cby_1__1__75_left_grid_pin_24_;
  wire [0:0] cby_1__1__75_left_grid_pin_25_;
  wire [0:0] cby_1__1__75_left_grid_pin_26_;
  wire [0:0] cby_1__1__75_left_grid_pin_27_;
  wire [0:0] cby_1__1__75_left_grid_pin_28_;
  wire [0:0] cby_1__1__75_left_grid_pin_29_;
  wire [0:0] cby_1__1__75_left_grid_pin_30_;
  wire [0:0] cby_1__1__75_left_grid_pin_31_;
  wire [0:0] cby_1__1__76_ccff_tail;
  wire [0:19] cby_1__1__76_chany_bottom_out;
  wire [0:19] cby_1__1__76_chany_top_out;
  wire [0:0] cby_1__1__76_left_grid_pin_16_;
  wire [0:0] cby_1__1__76_left_grid_pin_17_;
  wire [0:0] cby_1__1__76_left_grid_pin_18_;
  wire [0:0] cby_1__1__76_left_grid_pin_19_;
  wire [0:0] cby_1__1__76_left_grid_pin_20_;
  wire [0:0] cby_1__1__76_left_grid_pin_21_;
  wire [0:0] cby_1__1__76_left_grid_pin_22_;
  wire [0:0] cby_1__1__76_left_grid_pin_23_;
  wire [0:0] cby_1__1__76_left_grid_pin_24_;
  wire [0:0] cby_1__1__76_left_grid_pin_25_;
  wire [0:0] cby_1__1__76_left_grid_pin_26_;
  wire [0:0] cby_1__1__76_left_grid_pin_27_;
  wire [0:0] cby_1__1__76_left_grid_pin_28_;
  wire [0:0] cby_1__1__76_left_grid_pin_29_;
  wire [0:0] cby_1__1__76_left_grid_pin_30_;
  wire [0:0] cby_1__1__76_left_grid_pin_31_;
  wire [0:0] cby_1__1__77_ccff_tail;
  wire [0:19] cby_1__1__77_chany_bottom_out;
  wire [0:19] cby_1__1__77_chany_top_out;
  wire [0:0] cby_1__1__77_left_grid_pin_16_;
  wire [0:0] cby_1__1__77_left_grid_pin_17_;
  wire [0:0] cby_1__1__77_left_grid_pin_18_;
  wire [0:0] cby_1__1__77_left_grid_pin_19_;
  wire [0:0] cby_1__1__77_left_grid_pin_20_;
  wire [0:0] cby_1__1__77_left_grid_pin_21_;
  wire [0:0] cby_1__1__77_left_grid_pin_22_;
  wire [0:0] cby_1__1__77_left_grid_pin_23_;
  wire [0:0] cby_1__1__77_left_grid_pin_24_;
  wire [0:0] cby_1__1__77_left_grid_pin_25_;
  wire [0:0] cby_1__1__77_left_grid_pin_26_;
  wire [0:0] cby_1__1__77_left_grid_pin_27_;
  wire [0:0] cby_1__1__77_left_grid_pin_28_;
  wire [0:0] cby_1__1__77_left_grid_pin_29_;
  wire [0:0] cby_1__1__77_left_grid_pin_30_;
  wire [0:0] cby_1__1__77_left_grid_pin_31_;
  wire [0:0] cby_1__1__78_ccff_tail;
  wire [0:19] cby_1__1__78_chany_bottom_out;
  wire [0:19] cby_1__1__78_chany_top_out;
  wire [0:0] cby_1__1__78_left_grid_pin_16_;
  wire [0:0] cby_1__1__78_left_grid_pin_17_;
  wire [0:0] cby_1__1__78_left_grid_pin_18_;
  wire [0:0] cby_1__1__78_left_grid_pin_19_;
  wire [0:0] cby_1__1__78_left_grid_pin_20_;
  wire [0:0] cby_1__1__78_left_grid_pin_21_;
  wire [0:0] cby_1__1__78_left_grid_pin_22_;
  wire [0:0] cby_1__1__78_left_grid_pin_23_;
  wire [0:0] cby_1__1__78_left_grid_pin_24_;
  wire [0:0] cby_1__1__78_left_grid_pin_25_;
  wire [0:0] cby_1__1__78_left_grid_pin_26_;
  wire [0:0] cby_1__1__78_left_grid_pin_27_;
  wire [0:0] cby_1__1__78_left_grid_pin_28_;
  wire [0:0] cby_1__1__78_left_grid_pin_29_;
  wire [0:0] cby_1__1__78_left_grid_pin_30_;
  wire [0:0] cby_1__1__78_left_grid_pin_31_;
  wire [0:0] cby_1__1__79_ccff_tail;
  wire [0:19] cby_1__1__79_chany_bottom_out;
  wire [0:19] cby_1__1__79_chany_top_out;
  wire [0:0] cby_1__1__79_left_grid_pin_16_;
  wire [0:0] cby_1__1__79_left_grid_pin_17_;
  wire [0:0] cby_1__1__79_left_grid_pin_18_;
  wire [0:0] cby_1__1__79_left_grid_pin_19_;
  wire [0:0] cby_1__1__79_left_grid_pin_20_;
  wire [0:0] cby_1__1__79_left_grid_pin_21_;
  wire [0:0] cby_1__1__79_left_grid_pin_22_;
  wire [0:0] cby_1__1__79_left_grid_pin_23_;
  wire [0:0] cby_1__1__79_left_grid_pin_24_;
  wire [0:0] cby_1__1__79_left_grid_pin_25_;
  wire [0:0] cby_1__1__79_left_grid_pin_26_;
  wire [0:0] cby_1__1__79_left_grid_pin_27_;
  wire [0:0] cby_1__1__79_left_grid_pin_28_;
  wire [0:0] cby_1__1__79_left_grid_pin_29_;
  wire [0:0] cby_1__1__79_left_grid_pin_30_;
  wire [0:0] cby_1__1__79_left_grid_pin_31_;
  wire [0:0] cby_1__1__7_ccff_tail;
  wire [0:19] cby_1__1__7_chany_bottom_out;
  wire [0:19] cby_1__1__7_chany_top_out;
  wire [0:0] cby_1__1__7_left_grid_pin_16_;
  wire [0:0] cby_1__1__7_left_grid_pin_17_;
  wire [0:0] cby_1__1__7_left_grid_pin_18_;
  wire [0:0] cby_1__1__7_left_grid_pin_19_;
  wire [0:0] cby_1__1__7_left_grid_pin_20_;
  wire [0:0] cby_1__1__7_left_grid_pin_21_;
  wire [0:0] cby_1__1__7_left_grid_pin_22_;
  wire [0:0] cby_1__1__7_left_grid_pin_23_;
  wire [0:0] cby_1__1__7_left_grid_pin_24_;
  wire [0:0] cby_1__1__7_left_grid_pin_25_;
  wire [0:0] cby_1__1__7_left_grid_pin_26_;
  wire [0:0] cby_1__1__7_left_grid_pin_27_;
  wire [0:0] cby_1__1__7_left_grid_pin_28_;
  wire [0:0] cby_1__1__7_left_grid_pin_29_;
  wire [0:0] cby_1__1__7_left_grid_pin_30_;
  wire [0:0] cby_1__1__7_left_grid_pin_31_;
  wire [0:0] cby_1__1__80_ccff_tail;
  wire [0:19] cby_1__1__80_chany_bottom_out;
  wire [0:19] cby_1__1__80_chany_top_out;
  wire [0:0] cby_1__1__80_left_grid_pin_16_;
  wire [0:0] cby_1__1__80_left_grid_pin_17_;
  wire [0:0] cby_1__1__80_left_grid_pin_18_;
  wire [0:0] cby_1__1__80_left_grid_pin_19_;
  wire [0:0] cby_1__1__80_left_grid_pin_20_;
  wire [0:0] cby_1__1__80_left_grid_pin_21_;
  wire [0:0] cby_1__1__80_left_grid_pin_22_;
  wire [0:0] cby_1__1__80_left_grid_pin_23_;
  wire [0:0] cby_1__1__80_left_grid_pin_24_;
  wire [0:0] cby_1__1__80_left_grid_pin_25_;
  wire [0:0] cby_1__1__80_left_grid_pin_26_;
  wire [0:0] cby_1__1__80_left_grid_pin_27_;
  wire [0:0] cby_1__1__80_left_grid_pin_28_;
  wire [0:0] cby_1__1__80_left_grid_pin_29_;
  wire [0:0] cby_1__1__80_left_grid_pin_30_;
  wire [0:0] cby_1__1__80_left_grid_pin_31_;
  wire [0:0] cby_1__1__81_ccff_tail;
  wire [0:19] cby_1__1__81_chany_bottom_out;
  wire [0:19] cby_1__1__81_chany_top_out;
  wire [0:0] cby_1__1__81_left_grid_pin_16_;
  wire [0:0] cby_1__1__81_left_grid_pin_17_;
  wire [0:0] cby_1__1__81_left_grid_pin_18_;
  wire [0:0] cby_1__1__81_left_grid_pin_19_;
  wire [0:0] cby_1__1__81_left_grid_pin_20_;
  wire [0:0] cby_1__1__81_left_grid_pin_21_;
  wire [0:0] cby_1__1__81_left_grid_pin_22_;
  wire [0:0] cby_1__1__81_left_grid_pin_23_;
  wire [0:0] cby_1__1__81_left_grid_pin_24_;
  wire [0:0] cby_1__1__81_left_grid_pin_25_;
  wire [0:0] cby_1__1__81_left_grid_pin_26_;
  wire [0:0] cby_1__1__81_left_grid_pin_27_;
  wire [0:0] cby_1__1__81_left_grid_pin_28_;
  wire [0:0] cby_1__1__81_left_grid_pin_29_;
  wire [0:0] cby_1__1__81_left_grid_pin_30_;
  wire [0:0] cby_1__1__81_left_grid_pin_31_;
  wire [0:0] cby_1__1__82_ccff_tail;
  wire [0:19] cby_1__1__82_chany_bottom_out;
  wire [0:19] cby_1__1__82_chany_top_out;
  wire [0:0] cby_1__1__82_left_grid_pin_16_;
  wire [0:0] cby_1__1__82_left_grid_pin_17_;
  wire [0:0] cby_1__1__82_left_grid_pin_18_;
  wire [0:0] cby_1__1__82_left_grid_pin_19_;
  wire [0:0] cby_1__1__82_left_grid_pin_20_;
  wire [0:0] cby_1__1__82_left_grid_pin_21_;
  wire [0:0] cby_1__1__82_left_grid_pin_22_;
  wire [0:0] cby_1__1__82_left_grid_pin_23_;
  wire [0:0] cby_1__1__82_left_grid_pin_24_;
  wire [0:0] cby_1__1__82_left_grid_pin_25_;
  wire [0:0] cby_1__1__82_left_grid_pin_26_;
  wire [0:0] cby_1__1__82_left_grid_pin_27_;
  wire [0:0] cby_1__1__82_left_grid_pin_28_;
  wire [0:0] cby_1__1__82_left_grid_pin_29_;
  wire [0:0] cby_1__1__82_left_grid_pin_30_;
  wire [0:0] cby_1__1__82_left_grid_pin_31_;
  wire [0:0] cby_1__1__83_ccff_tail;
  wire [0:19] cby_1__1__83_chany_bottom_out;
  wire [0:19] cby_1__1__83_chany_top_out;
  wire [0:0] cby_1__1__83_left_grid_pin_16_;
  wire [0:0] cby_1__1__83_left_grid_pin_17_;
  wire [0:0] cby_1__1__83_left_grid_pin_18_;
  wire [0:0] cby_1__1__83_left_grid_pin_19_;
  wire [0:0] cby_1__1__83_left_grid_pin_20_;
  wire [0:0] cby_1__1__83_left_grid_pin_21_;
  wire [0:0] cby_1__1__83_left_grid_pin_22_;
  wire [0:0] cby_1__1__83_left_grid_pin_23_;
  wire [0:0] cby_1__1__83_left_grid_pin_24_;
  wire [0:0] cby_1__1__83_left_grid_pin_25_;
  wire [0:0] cby_1__1__83_left_grid_pin_26_;
  wire [0:0] cby_1__1__83_left_grid_pin_27_;
  wire [0:0] cby_1__1__83_left_grid_pin_28_;
  wire [0:0] cby_1__1__83_left_grid_pin_29_;
  wire [0:0] cby_1__1__83_left_grid_pin_30_;
  wire [0:0] cby_1__1__83_left_grid_pin_31_;
  wire [0:0] cby_1__1__84_ccff_tail;
  wire [0:19] cby_1__1__84_chany_bottom_out;
  wire [0:19] cby_1__1__84_chany_top_out;
  wire [0:0] cby_1__1__84_left_grid_pin_16_;
  wire [0:0] cby_1__1__84_left_grid_pin_17_;
  wire [0:0] cby_1__1__84_left_grid_pin_18_;
  wire [0:0] cby_1__1__84_left_grid_pin_19_;
  wire [0:0] cby_1__1__84_left_grid_pin_20_;
  wire [0:0] cby_1__1__84_left_grid_pin_21_;
  wire [0:0] cby_1__1__84_left_grid_pin_22_;
  wire [0:0] cby_1__1__84_left_grid_pin_23_;
  wire [0:0] cby_1__1__84_left_grid_pin_24_;
  wire [0:0] cby_1__1__84_left_grid_pin_25_;
  wire [0:0] cby_1__1__84_left_grid_pin_26_;
  wire [0:0] cby_1__1__84_left_grid_pin_27_;
  wire [0:0] cby_1__1__84_left_grid_pin_28_;
  wire [0:0] cby_1__1__84_left_grid_pin_29_;
  wire [0:0] cby_1__1__84_left_grid_pin_30_;
  wire [0:0] cby_1__1__84_left_grid_pin_31_;
  wire [0:0] cby_1__1__85_ccff_tail;
  wire [0:19] cby_1__1__85_chany_bottom_out;
  wire [0:19] cby_1__1__85_chany_top_out;
  wire [0:0] cby_1__1__85_left_grid_pin_16_;
  wire [0:0] cby_1__1__85_left_grid_pin_17_;
  wire [0:0] cby_1__1__85_left_grid_pin_18_;
  wire [0:0] cby_1__1__85_left_grid_pin_19_;
  wire [0:0] cby_1__1__85_left_grid_pin_20_;
  wire [0:0] cby_1__1__85_left_grid_pin_21_;
  wire [0:0] cby_1__1__85_left_grid_pin_22_;
  wire [0:0] cby_1__1__85_left_grid_pin_23_;
  wire [0:0] cby_1__1__85_left_grid_pin_24_;
  wire [0:0] cby_1__1__85_left_grid_pin_25_;
  wire [0:0] cby_1__1__85_left_grid_pin_26_;
  wire [0:0] cby_1__1__85_left_grid_pin_27_;
  wire [0:0] cby_1__1__85_left_grid_pin_28_;
  wire [0:0] cby_1__1__85_left_grid_pin_29_;
  wire [0:0] cby_1__1__85_left_grid_pin_30_;
  wire [0:0] cby_1__1__85_left_grid_pin_31_;
  wire [0:0] cby_1__1__86_ccff_tail;
  wire [0:19] cby_1__1__86_chany_bottom_out;
  wire [0:19] cby_1__1__86_chany_top_out;
  wire [0:0] cby_1__1__86_left_grid_pin_16_;
  wire [0:0] cby_1__1__86_left_grid_pin_17_;
  wire [0:0] cby_1__1__86_left_grid_pin_18_;
  wire [0:0] cby_1__1__86_left_grid_pin_19_;
  wire [0:0] cby_1__1__86_left_grid_pin_20_;
  wire [0:0] cby_1__1__86_left_grid_pin_21_;
  wire [0:0] cby_1__1__86_left_grid_pin_22_;
  wire [0:0] cby_1__1__86_left_grid_pin_23_;
  wire [0:0] cby_1__1__86_left_grid_pin_24_;
  wire [0:0] cby_1__1__86_left_grid_pin_25_;
  wire [0:0] cby_1__1__86_left_grid_pin_26_;
  wire [0:0] cby_1__1__86_left_grid_pin_27_;
  wire [0:0] cby_1__1__86_left_grid_pin_28_;
  wire [0:0] cby_1__1__86_left_grid_pin_29_;
  wire [0:0] cby_1__1__86_left_grid_pin_30_;
  wire [0:0] cby_1__1__86_left_grid_pin_31_;
  wire [0:0] cby_1__1__87_ccff_tail;
  wire [0:19] cby_1__1__87_chany_bottom_out;
  wire [0:19] cby_1__1__87_chany_top_out;
  wire [0:0] cby_1__1__87_left_grid_pin_16_;
  wire [0:0] cby_1__1__87_left_grid_pin_17_;
  wire [0:0] cby_1__1__87_left_grid_pin_18_;
  wire [0:0] cby_1__1__87_left_grid_pin_19_;
  wire [0:0] cby_1__1__87_left_grid_pin_20_;
  wire [0:0] cby_1__1__87_left_grid_pin_21_;
  wire [0:0] cby_1__1__87_left_grid_pin_22_;
  wire [0:0] cby_1__1__87_left_grid_pin_23_;
  wire [0:0] cby_1__1__87_left_grid_pin_24_;
  wire [0:0] cby_1__1__87_left_grid_pin_25_;
  wire [0:0] cby_1__1__87_left_grid_pin_26_;
  wire [0:0] cby_1__1__87_left_grid_pin_27_;
  wire [0:0] cby_1__1__87_left_grid_pin_28_;
  wire [0:0] cby_1__1__87_left_grid_pin_29_;
  wire [0:0] cby_1__1__87_left_grid_pin_30_;
  wire [0:0] cby_1__1__87_left_grid_pin_31_;
  wire [0:0] cby_1__1__88_ccff_tail;
  wire [0:19] cby_1__1__88_chany_bottom_out;
  wire [0:19] cby_1__1__88_chany_top_out;
  wire [0:0] cby_1__1__88_left_grid_pin_16_;
  wire [0:0] cby_1__1__88_left_grid_pin_17_;
  wire [0:0] cby_1__1__88_left_grid_pin_18_;
  wire [0:0] cby_1__1__88_left_grid_pin_19_;
  wire [0:0] cby_1__1__88_left_grid_pin_20_;
  wire [0:0] cby_1__1__88_left_grid_pin_21_;
  wire [0:0] cby_1__1__88_left_grid_pin_22_;
  wire [0:0] cby_1__1__88_left_grid_pin_23_;
  wire [0:0] cby_1__1__88_left_grid_pin_24_;
  wire [0:0] cby_1__1__88_left_grid_pin_25_;
  wire [0:0] cby_1__1__88_left_grid_pin_26_;
  wire [0:0] cby_1__1__88_left_grid_pin_27_;
  wire [0:0] cby_1__1__88_left_grid_pin_28_;
  wire [0:0] cby_1__1__88_left_grid_pin_29_;
  wire [0:0] cby_1__1__88_left_grid_pin_30_;
  wire [0:0] cby_1__1__88_left_grid_pin_31_;
  wire [0:0] cby_1__1__89_ccff_tail;
  wire [0:19] cby_1__1__89_chany_bottom_out;
  wire [0:19] cby_1__1__89_chany_top_out;
  wire [0:0] cby_1__1__89_left_grid_pin_16_;
  wire [0:0] cby_1__1__89_left_grid_pin_17_;
  wire [0:0] cby_1__1__89_left_grid_pin_18_;
  wire [0:0] cby_1__1__89_left_grid_pin_19_;
  wire [0:0] cby_1__1__89_left_grid_pin_20_;
  wire [0:0] cby_1__1__89_left_grid_pin_21_;
  wire [0:0] cby_1__1__89_left_grid_pin_22_;
  wire [0:0] cby_1__1__89_left_grid_pin_23_;
  wire [0:0] cby_1__1__89_left_grid_pin_24_;
  wire [0:0] cby_1__1__89_left_grid_pin_25_;
  wire [0:0] cby_1__1__89_left_grid_pin_26_;
  wire [0:0] cby_1__1__89_left_grid_pin_27_;
  wire [0:0] cby_1__1__89_left_grid_pin_28_;
  wire [0:0] cby_1__1__89_left_grid_pin_29_;
  wire [0:0] cby_1__1__89_left_grid_pin_30_;
  wire [0:0] cby_1__1__89_left_grid_pin_31_;
  wire [0:0] cby_1__1__8_ccff_tail;
  wire [0:19] cby_1__1__8_chany_bottom_out;
  wire [0:19] cby_1__1__8_chany_top_out;
  wire [0:0] cby_1__1__8_left_grid_pin_16_;
  wire [0:0] cby_1__1__8_left_grid_pin_17_;
  wire [0:0] cby_1__1__8_left_grid_pin_18_;
  wire [0:0] cby_1__1__8_left_grid_pin_19_;
  wire [0:0] cby_1__1__8_left_grid_pin_20_;
  wire [0:0] cby_1__1__8_left_grid_pin_21_;
  wire [0:0] cby_1__1__8_left_grid_pin_22_;
  wire [0:0] cby_1__1__8_left_grid_pin_23_;
  wire [0:0] cby_1__1__8_left_grid_pin_24_;
  wire [0:0] cby_1__1__8_left_grid_pin_25_;
  wire [0:0] cby_1__1__8_left_grid_pin_26_;
  wire [0:0] cby_1__1__8_left_grid_pin_27_;
  wire [0:0] cby_1__1__8_left_grid_pin_28_;
  wire [0:0] cby_1__1__8_left_grid_pin_29_;
  wire [0:0] cby_1__1__8_left_grid_pin_30_;
  wire [0:0] cby_1__1__8_left_grid_pin_31_;
  wire [0:0] cby_1__1__90_ccff_tail;
  wire [0:19] cby_1__1__90_chany_bottom_out;
  wire [0:19] cby_1__1__90_chany_top_out;
  wire [0:0] cby_1__1__90_left_grid_pin_16_;
  wire [0:0] cby_1__1__90_left_grid_pin_17_;
  wire [0:0] cby_1__1__90_left_grid_pin_18_;
  wire [0:0] cby_1__1__90_left_grid_pin_19_;
  wire [0:0] cby_1__1__90_left_grid_pin_20_;
  wire [0:0] cby_1__1__90_left_grid_pin_21_;
  wire [0:0] cby_1__1__90_left_grid_pin_22_;
  wire [0:0] cby_1__1__90_left_grid_pin_23_;
  wire [0:0] cby_1__1__90_left_grid_pin_24_;
  wire [0:0] cby_1__1__90_left_grid_pin_25_;
  wire [0:0] cby_1__1__90_left_grid_pin_26_;
  wire [0:0] cby_1__1__90_left_grid_pin_27_;
  wire [0:0] cby_1__1__90_left_grid_pin_28_;
  wire [0:0] cby_1__1__90_left_grid_pin_29_;
  wire [0:0] cby_1__1__90_left_grid_pin_30_;
  wire [0:0] cby_1__1__90_left_grid_pin_31_;
  wire [0:0] cby_1__1__91_ccff_tail;
  wire [0:19] cby_1__1__91_chany_bottom_out;
  wire [0:19] cby_1__1__91_chany_top_out;
  wire [0:0] cby_1__1__91_left_grid_pin_16_;
  wire [0:0] cby_1__1__91_left_grid_pin_17_;
  wire [0:0] cby_1__1__91_left_grid_pin_18_;
  wire [0:0] cby_1__1__91_left_grid_pin_19_;
  wire [0:0] cby_1__1__91_left_grid_pin_20_;
  wire [0:0] cby_1__1__91_left_grid_pin_21_;
  wire [0:0] cby_1__1__91_left_grid_pin_22_;
  wire [0:0] cby_1__1__91_left_grid_pin_23_;
  wire [0:0] cby_1__1__91_left_grid_pin_24_;
  wire [0:0] cby_1__1__91_left_grid_pin_25_;
  wire [0:0] cby_1__1__91_left_grid_pin_26_;
  wire [0:0] cby_1__1__91_left_grid_pin_27_;
  wire [0:0] cby_1__1__91_left_grid_pin_28_;
  wire [0:0] cby_1__1__91_left_grid_pin_29_;
  wire [0:0] cby_1__1__91_left_grid_pin_30_;
  wire [0:0] cby_1__1__91_left_grid_pin_31_;
  wire [0:0] cby_1__1__92_ccff_tail;
  wire [0:19] cby_1__1__92_chany_bottom_out;
  wire [0:19] cby_1__1__92_chany_top_out;
  wire [0:0] cby_1__1__92_left_grid_pin_16_;
  wire [0:0] cby_1__1__92_left_grid_pin_17_;
  wire [0:0] cby_1__1__92_left_grid_pin_18_;
  wire [0:0] cby_1__1__92_left_grid_pin_19_;
  wire [0:0] cby_1__1__92_left_grid_pin_20_;
  wire [0:0] cby_1__1__92_left_grid_pin_21_;
  wire [0:0] cby_1__1__92_left_grid_pin_22_;
  wire [0:0] cby_1__1__92_left_grid_pin_23_;
  wire [0:0] cby_1__1__92_left_grid_pin_24_;
  wire [0:0] cby_1__1__92_left_grid_pin_25_;
  wire [0:0] cby_1__1__92_left_grid_pin_26_;
  wire [0:0] cby_1__1__92_left_grid_pin_27_;
  wire [0:0] cby_1__1__92_left_grid_pin_28_;
  wire [0:0] cby_1__1__92_left_grid_pin_29_;
  wire [0:0] cby_1__1__92_left_grid_pin_30_;
  wire [0:0] cby_1__1__92_left_grid_pin_31_;
  wire [0:0] cby_1__1__93_ccff_tail;
  wire [0:19] cby_1__1__93_chany_bottom_out;
  wire [0:19] cby_1__1__93_chany_top_out;
  wire [0:0] cby_1__1__93_left_grid_pin_16_;
  wire [0:0] cby_1__1__93_left_grid_pin_17_;
  wire [0:0] cby_1__1__93_left_grid_pin_18_;
  wire [0:0] cby_1__1__93_left_grid_pin_19_;
  wire [0:0] cby_1__1__93_left_grid_pin_20_;
  wire [0:0] cby_1__1__93_left_grid_pin_21_;
  wire [0:0] cby_1__1__93_left_grid_pin_22_;
  wire [0:0] cby_1__1__93_left_grid_pin_23_;
  wire [0:0] cby_1__1__93_left_grid_pin_24_;
  wire [0:0] cby_1__1__93_left_grid_pin_25_;
  wire [0:0] cby_1__1__93_left_grid_pin_26_;
  wire [0:0] cby_1__1__93_left_grid_pin_27_;
  wire [0:0] cby_1__1__93_left_grid_pin_28_;
  wire [0:0] cby_1__1__93_left_grid_pin_29_;
  wire [0:0] cby_1__1__93_left_grid_pin_30_;
  wire [0:0] cby_1__1__93_left_grid_pin_31_;
  wire [0:0] cby_1__1__94_ccff_tail;
  wire [0:19] cby_1__1__94_chany_bottom_out;
  wire [0:19] cby_1__1__94_chany_top_out;
  wire [0:0] cby_1__1__94_left_grid_pin_16_;
  wire [0:0] cby_1__1__94_left_grid_pin_17_;
  wire [0:0] cby_1__1__94_left_grid_pin_18_;
  wire [0:0] cby_1__1__94_left_grid_pin_19_;
  wire [0:0] cby_1__1__94_left_grid_pin_20_;
  wire [0:0] cby_1__1__94_left_grid_pin_21_;
  wire [0:0] cby_1__1__94_left_grid_pin_22_;
  wire [0:0] cby_1__1__94_left_grid_pin_23_;
  wire [0:0] cby_1__1__94_left_grid_pin_24_;
  wire [0:0] cby_1__1__94_left_grid_pin_25_;
  wire [0:0] cby_1__1__94_left_grid_pin_26_;
  wire [0:0] cby_1__1__94_left_grid_pin_27_;
  wire [0:0] cby_1__1__94_left_grid_pin_28_;
  wire [0:0] cby_1__1__94_left_grid_pin_29_;
  wire [0:0] cby_1__1__94_left_grid_pin_30_;
  wire [0:0] cby_1__1__94_left_grid_pin_31_;
  wire [0:0] cby_1__1__95_ccff_tail;
  wire [0:19] cby_1__1__95_chany_bottom_out;
  wire [0:19] cby_1__1__95_chany_top_out;
  wire [0:0] cby_1__1__95_left_grid_pin_16_;
  wire [0:0] cby_1__1__95_left_grid_pin_17_;
  wire [0:0] cby_1__1__95_left_grid_pin_18_;
  wire [0:0] cby_1__1__95_left_grid_pin_19_;
  wire [0:0] cby_1__1__95_left_grid_pin_20_;
  wire [0:0] cby_1__1__95_left_grid_pin_21_;
  wire [0:0] cby_1__1__95_left_grid_pin_22_;
  wire [0:0] cby_1__1__95_left_grid_pin_23_;
  wire [0:0] cby_1__1__95_left_grid_pin_24_;
  wire [0:0] cby_1__1__95_left_grid_pin_25_;
  wire [0:0] cby_1__1__95_left_grid_pin_26_;
  wire [0:0] cby_1__1__95_left_grid_pin_27_;
  wire [0:0] cby_1__1__95_left_grid_pin_28_;
  wire [0:0] cby_1__1__95_left_grid_pin_29_;
  wire [0:0] cby_1__1__95_left_grid_pin_30_;
  wire [0:0] cby_1__1__95_left_grid_pin_31_;
  wire [0:0] cby_1__1__96_ccff_tail;
  wire [0:19] cby_1__1__96_chany_bottom_out;
  wire [0:19] cby_1__1__96_chany_top_out;
  wire [0:0] cby_1__1__96_left_grid_pin_16_;
  wire [0:0] cby_1__1__96_left_grid_pin_17_;
  wire [0:0] cby_1__1__96_left_grid_pin_18_;
  wire [0:0] cby_1__1__96_left_grid_pin_19_;
  wire [0:0] cby_1__1__96_left_grid_pin_20_;
  wire [0:0] cby_1__1__96_left_grid_pin_21_;
  wire [0:0] cby_1__1__96_left_grid_pin_22_;
  wire [0:0] cby_1__1__96_left_grid_pin_23_;
  wire [0:0] cby_1__1__96_left_grid_pin_24_;
  wire [0:0] cby_1__1__96_left_grid_pin_25_;
  wire [0:0] cby_1__1__96_left_grid_pin_26_;
  wire [0:0] cby_1__1__96_left_grid_pin_27_;
  wire [0:0] cby_1__1__96_left_grid_pin_28_;
  wire [0:0] cby_1__1__96_left_grid_pin_29_;
  wire [0:0] cby_1__1__96_left_grid_pin_30_;
  wire [0:0] cby_1__1__96_left_grid_pin_31_;
  wire [0:0] cby_1__1__97_ccff_tail;
  wire [0:19] cby_1__1__97_chany_bottom_out;
  wire [0:19] cby_1__1__97_chany_top_out;
  wire [0:0] cby_1__1__97_left_grid_pin_16_;
  wire [0:0] cby_1__1__97_left_grid_pin_17_;
  wire [0:0] cby_1__1__97_left_grid_pin_18_;
  wire [0:0] cby_1__1__97_left_grid_pin_19_;
  wire [0:0] cby_1__1__97_left_grid_pin_20_;
  wire [0:0] cby_1__1__97_left_grid_pin_21_;
  wire [0:0] cby_1__1__97_left_grid_pin_22_;
  wire [0:0] cby_1__1__97_left_grid_pin_23_;
  wire [0:0] cby_1__1__97_left_grid_pin_24_;
  wire [0:0] cby_1__1__97_left_grid_pin_25_;
  wire [0:0] cby_1__1__97_left_grid_pin_26_;
  wire [0:0] cby_1__1__97_left_grid_pin_27_;
  wire [0:0] cby_1__1__97_left_grid_pin_28_;
  wire [0:0] cby_1__1__97_left_grid_pin_29_;
  wire [0:0] cby_1__1__97_left_grid_pin_30_;
  wire [0:0] cby_1__1__97_left_grid_pin_31_;
  wire [0:0] cby_1__1__98_ccff_tail;
  wire [0:19] cby_1__1__98_chany_bottom_out;
  wire [0:19] cby_1__1__98_chany_top_out;
  wire [0:0] cby_1__1__98_left_grid_pin_16_;
  wire [0:0] cby_1__1__98_left_grid_pin_17_;
  wire [0:0] cby_1__1__98_left_grid_pin_18_;
  wire [0:0] cby_1__1__98_left_grid_pin_19_;
  wire [0:0] cby_1__1__98_left_grid_pin_20_;
  wire [0:0] cby_1__1__98_left_grid_pin_21_;
  wire [0:0] cby_1__1__98_left_grid_pin_22_;
  wire [0:0] cby_1__1__98_left_grid_pin_23_;
  wire [0:0] cby_1__1__98_left_grid_pin_24_;
  wire [0:0] cby_1__1__98_left_grid_pin_25_;
  wire [0:0] cby_1__1__98_left_grid_pin_26_;
  wire [0:0] cby_1__1__98_left_grid_pin_27_;
  wire [0:0] cby_1__1__98_left_grid_pin_28_;
  wire [0:0] cby_1__1__98_left_grid_pin_29_;
  wire [0:0] cby_1__1__98_left_grid_pin_30_;
  wire [0:0] cby_1__1__98_left_grid_pin_31_;
  wire [0:0] cby_1__1__99_ccff_tail;
  wire [0:19] cby_1__1__99_chany_bottom_out;
  wire [0:19] cby_1__1__99_chany_top_out;
  wire [0:0] cby_1__1__99_left_grid_pin_16_;
  wire [0:0] cby_1__1__99_left_grid_pin_17_;
  wire [0:0] cby_1__1__99_left_grid_pin_18_;
  wire [0:0] cby_1__1__99_left_grid_pin_19_;
  wire [0:0] cby_1__1__99_left_grid_pin_20_;
  wire [0:0] cby_1__1__99_left_grid_pin_21_;
  wire [0:0] cby_1__1__99_left_grid_pin_22_;
  wire [0:0] cby_1__1__99_left_grid_pin_23_;
  wire [0:0] cby_1__1__99_left_grid_pin_24_;
  wire [0:0] cby_1__1__99_left_grid_pin_25_;
  wire [0:0] cby_1__1__99_left_grid_pin_26_;
  wire [0:0] cby_1__1__99_left_grid_pin_27_;
  wire [0:0] cby_1__1__99_left_grid_pin_28_;
  wire [0:0] cby_1__1__99_left_grid_pin_29_;
  wire [0:0] cby_1__1__99_left_grid_pin_30_;
  wire [0:0] cby_1__1__99_left_grid_pin_31_;
  wire [0:0] cby_1__1__9_ccff_tail;
  wire [0:19] cby_1__1__9_chany_bottom_out;
  wire [0:19] cby_1__1__9_chany_top_out;
  wire [0:0] cby_1__1__9_left_grid_pin_16_;
  wire [0:0] cby_1__1__9_left_grid_pin_17_;
  wire [0:0] cby_1__1__9_left_grid_pin_18_;
  wire [0:0] cby_1__1__9_left_grid_pin_19_;
  wire [0:0] cby_1__1__9_left_grid_pin_20_;
  wire [0:0] cby_1__1__9_left_grid_pin_21_;
  wire [0:0] cby_1__1__9_left_grid_pin_22_;
  wire [0:0] cby_1__1__9_left_grid_pin_23_;
  wire [0:0] cby_1__1__9_left_grid_pin_24_;
  wire [0:0] cby_1__1__9_left_grid_pin_25_;
  wire [0:0] cby_1__1__9_left_grid_pin_26_;
  wire [0:0] cby_1__1__9_left_grid_pin_27_;
  wire [0:0] cby_1__1__9_left_grid_pin_28_;
  wire [0:0] cby_1__1__9_left_grid_pin_29_;
  wire [0:0] cby_1__1__9_left_grid_pin_30_;
  wire [0:0] cby_1__1__9_left_grid_pin_31_;
  wire [0:0] direct_interc_0_out;
  wire [0:0] direct_interc_100_out;
  wire [0:0] direct_interc_101_out;
  wire [0:0] direct_interc_102_out;
  wire [0:0] direct_interc_103_out;
  wire [0:0] direct_interc_104_out;
  wire [0:0] direct_interc_105_out;
  wire [0:0] direct_interc_106_out;
  wire [0:0] direct_interc_107_out;
  wire [0:0] direct_interc_108_out;
  wire [0:0] direct_interc_109_out;
  wire [0:0] direct_interc_10_out;
  wire [0:0] direct_interc_110_out;
  wire [0:0] direct_interc_111_out;
  wire [0:0] direct_interc_112_out;
  wire [0:0] direct_interc_113_out;
  wire [0:0] direct_interc_114_out;
  wire [0:0] direct_interc_115_out;
  wire [0:0] direct_interc_116_out;
  wire [0:0] direct_interc_117_out;
  wire [0:0] direct_interc_118_out;
  wire [0:0] direct_interc_119_out;
  wire [0:0] direct_interc_11_out;
  wire [0:0] direct_interc_120_out;
  wire [0:0] direct_interc_121_out;
  wire [0:0] direct_interc_122_out;
  wire [0:0] direct_interc_123_out;
  wire [0:0] direct_interc_124_out;
  wire [0:0] direct_interc_125_out;
  wire [0:0] direct_interc_126_out;
  wire [0:0] direct_interc_127_out;
  wire [0:0] direct_interc_128_out;
  wire [0:0] direct_interc_129_out;
  wire [0:0] direct_interc_12_out;
  wire [0:0] direct_interc_130_out;
  wire [0:0] direct_interc_131_out;
  wire [0:0] direct_interc_132_out;
  wire [0:0] direct_interc_133_out;
  wire [0:0] direct_interc_134_out;
  wire [0:0] direct_interc_135_out;
  wire [0:0] direct_interc_136_out;
  wire [0:0] direct_interc_137_out;
  wire [0:0] direct_interc_138_out;
  wire [0:0] direct_interc_139_out;
  wire [0:0] direct_interc_13_out;
  wire [0:0] direct_interc_140_out;
  wire [0:0] direct_interc_141_out;
  wire [0:0] direct_interc_142_out;
  wire [0:0] direct_interc_143_out;
  wire [0:0] direct_interc_144_out;
  wire [0:0] direct_interc_145_out;
  wire [0:0] direct_interc_146_out;
  wire [0:0] direct_interc_147_out;
  wire [0:0] direct_interc_148_out;
  wire [0:0] direct_interc_149_out;
  wire [0:0] direct_interc_14_out;
  wire [0:0] direct_interc_150_out;
  wire [0:0] direct_interc_151_out;
  wire [0:0] direct_interc_152_out;
  wire [0:0] direct_interc_153_out;
  wire [0:0] direct_interc_154_out;
  wire [0:0] direct_interc_155_out;
  wire [0:0] direct_interc_156_out;
  wire [0:0] direct_interc_157_out;
  wire [0:0] direct_interc_158_out;
  wire [0:0] direct_interc_159_out;
  wire [0:0] direct_interc_15_out;
  wire [0:0] direct_interc_160_out;
  wire [0:0] direct_interc_161_out;
  wire [0:0] direct_interc_162_out;
  wire [0:0] direct_interc_163_out;
  wire [0:0] direct_interc_164_out;
  wire [0:0] direct_interc_165_out;
  wire [0:0] direct_interc_166_out;
  wire [0:0] direct_interc_167_out;
  wire [0:0] direct_interc_168_out;
  wire [0:0] direct_interc_169_out;
  wire [0:0] direct_interc_16_out;
  wire [0:0] direct_interc_170_out;
  wire [0:0] direct_interc_171_out;
  wire [0:0] direct_interc_172_out;
  wire [0:0] direct_interc_173_out;
  wire [0:0] direct_interc_174_out;
  wire [0:0] direct_interc_175_out;
  wire [0:0] direct_interc_176_out;
  wire [0:0] direct_interc_177_out;
  wire [0:0] direct_interc_178_out;
  wire [0:0] direct_interc_179_out;
  wire [0:0] direct_interc_17_out;
  wire [0:0] direct_interc_180_out;
  wire [0:0] direct_interc_181_out;
  wire [0:0] direct_interc_182_out;
  wire [0:0] direct_interc_183_out;
  wire [0:0] direct_interc_184_out;
  wire [0:0] direct_interc_185_out;
  wire [0:0] direct_interc_186_out;
  wire [0:0] direct_interc_187_out;
  wire [0:0] direct_interc_188_out;
  wire [0:0] direct_interc_189_out;
  wire [0:0] direct_interc_18_out;
  wire [0:0] direct_interc_190_out;
  wire [0:0] direct_interc_191_out;
  wire [0:0] direct_interc_192_out;
  wire [0:0] direct_interc_193_out;
  wire [0:0] direct_interc_194_out;
  wire [0:0] direct_interc_195_out;
  wire [0:0] direct_interc_196_out;
  wire [0:0] direct_interc_197_out;
  wire [0:0] direct_interc_198_out;
  wire [0:0] direct_interc_199_out;
  wire [0:0] direct_interc_19_out;
  wire [0:0] direct_interc_1_out;
  wire [0:0] direct_interc_200_out;
  wire [0:0] direct_interc_201_out;
  wire [0:0] direct_interc_202_out;
  wire [0:0] direct_interc_203_out;
  wire [0:0] direct_interc_204_out;
  wire [0:0] direct_interc_205_out;
  wire [0:0] direct_interc_206_out;
  wire [0:0] direct_interc_207_out;
  wire [0:0] direct_interc_208_out;
  wire [0:0] direct_interc_209_out;
  wire [0:0] direct_interc_20_out;
  wire [0:0] direct_interc_210_out;
  wire [0:0] direct_interc_211_out;
  wire [0:0] direct_interc_212_out;
  wire [0:0] direct_interc_213_out;
  wire [0:0] direct_interc_214_out;
  wire [0:0] direct_interc_215_out;
  wire [0:0] direct_interc_216_out;
  wire [0:0] direct_interc_217_out;
  wire [0:0] direct_interc_218_out;
  wire [0:0] direct_interc_219_out;
  wire [0:0] direct_interc_21_out;
  wire [0:0] direct_interc_220_out;
  wire [0:0] direct_interc_221_out;
  wire [0:0] direct_interc_222_out;
  wire [0:0] direct_interc_223_out;
  wire [0:0] direct_interc_224_out;
  wire [0:0] direct_interc_225_out;
  wire [0:0] direct_interc_226_out;
  wire [0:0] direct_interc_227_out;
  wire [0:0] direct_interc_228_out;
  wire [0:0] direct_interc_229_out;
  wire [0:0] direct_interc_22_out;
  wire [0:0] direct_interc_230_out;
  wire [0:0] direct_interc_231_out;
  wire [0:0] direct_interc_232_out;
  wire [0:0] direct_interc_233_out;
  wire [0:0] direct_interc_234_out;
  wire [0:0] direct_interc_235_out;
  wire [0:0] direct_interc_236_out;
  wire [0:0] direct_interc_237_out;
  wire [0:0] direct_interc_238_out;
  wire [0:0] direct_interc_239_out;
  wire [0:0] direct_interc_23_out;
  wire [0:0] direct_interc_240_out;
  wire [0:0] direct_interc_241_out;
  wire [0:0] direct_interc_242_out;
  wire [0:0] direct_interc_243_out;
  wire [0:0] direct_interc_244_out;
  wire [0:0] direct_interc_245_out;
  wire [0:0] direct_interc_246_out;
  wire [0:0] direct_interc_247_out;
  wire [0:0] direct_interc_248_out;
  wire [0:0] direct_interc_249_out;
  wire [0:0] direct_interc_24_out;
  wire [0:0] direct_interc_250_out;
  wire [0:0] direct_interc_251_out;
  wire [0:0] direct_interc_252_out;
  wire [0:0] direct_interc_253_out;
  wire [0:0] direct_interc_254_out;
  wire [0:0] direct_interc_255_out;
  wire [0:0] direct_interc_256_out;
  wire [0:0] direct_interc_257_out;
  wire [0:0] direct_interc_258_out;
  wire [0:0] direct_interc_259_out;
  wire [0:0] direct_interc_25_out;
  wire [0:0] direct_interc_260_out;
  wire [0:0] direct_interc_261_out;
  wire [0:0] direct_interc_262_out;
  wire [0:0] direct_interc_263_out;
  wire [0:0] direct_interc_264_out;
  wire [0:0] direct_interc_265_out;
  wire [0:0] direct_interc_266_out;
  wire [0:0] direct_interc_267_out;
  wire [0:0] direct_interc_268_out;
  wire [0:0] direct_interc_269_out;
  wire [0:0] direct_interc_26_out;
  wire [0:0] direct_interc_270_out;
  wire [0:0] direct_interc_271_out;
  wire [0:0] direct_interc_272_out;
  wire [0:0] direct_interc_273_out;
  wire [0:0] direct_interc_274_out;
  wire [0:0] direct_interc_27_out;
  wire [0:0] direct_interc_28_out;
  wire [0:0] direct_interc_29_out;
  wire [0:0] direct_interc_2_out;
  wire [0:0] direct_interc_30_out;
  wire [0:0] direct_interc_31_out;
  wire [0:0] direct_interc_32_out;
  wire [0:0] direct_interc_33_out;
  wire [0:0] direct_interc_34_out;
  wire [0:0] direct_interc_35_out;
  wire [0:0] direct_interc_36_out;
  wire [0:0] direct_interc_37_out;
  wire [0:0] direct_interc_38_out;
  wire [0:0] direct_interc_39_out;
  wire [0:0] direct_interc_3_out;
  wire [0:0] direct_interc_40_out;
  wire [0:0] direct_interc_41_out;
  wire [0:0] direct_interc_42_out;
  wire [0:0] direct_interc_43_out;
  wire [0:0] direct_interc_44_out;
  wire [0:0] direct_interc_45_out;
  wire [0:0] direct_interc_46_out;
  wire [0:0] direct_interc_47_out;
  wire [0:0] direct_interc_48_out;
  wire [0:0] direct_interc_49_out;
  wire [0:0] direct_interc_4_out;
  wire [0:0] direct_interc_50_out;
  wire [0:0] direct_interc_51_out;
  wire [0:0] direct_interc_52_out;
  wire [0:0] direct_interc_53_out;
  wire [0:0] direct_interc_54_out;
  wire [0:0] direct_interc_55_out;
  wire [0:0] direct_interc_56_out;
  wire [0:0] direct_interc_57_out;
  wire [0:0] direct_interc_58_out;
  wire [0:0] direct_interc_59_out;
  wire [0:0] direct_interc_5_out;
  wire [0:0] direct_interc_60_out;
  wire [0:0] direct_interc_61_out;
  wire [0:0] direct_interc_62_out;
  wire [0:0] direct_interc_63_out;
  wire [0:0] direct_interc_64_out;
  wire [0:0] direct_interc_65_out;
  wire [0:0] direct_interc_66_out;
  wire [0:0] direct_interc_67_out;
  wire [0:0] direct_interc_68_out;
  wire [0:0] direct_interc_69_out;
  wire [0:0] direct_interc_6_out;
  wire [0:0] direct_interc_70_out;
  wire [0:0] direct_interc_71_out;
  wire [0:0] direct_interc_72_out;
  wire [0:0] direct_interc_73_out;
  wire [0:0] direct_interc_74_out;
  wire [0:0] direct_interc_75_out;
  wire [0:0] direct_interc_76_out;
  wire [0:0] direct_interc_77_out;
  wire [0:0] direct_interc_78_out;
  wire [0:0] direct_interc_79_out;
  wire [0:0] direct_interc_7_out;
  wire [0:0] direct_interc_80_out;
  wire [0:0] direct_interc_81_out;
  wire [0:0] direct_interc_82_out;
  wire [0:0] direct_interc_83_out;
  wire [0:0] direct_interc_84_out;
  wire [0:0] direct_interc_85_out;
  wire [0:0] direct_interc_86_out;
  wire [0:0] direct_interc_87_out;
  wire [0:0] direct_interc_88_out;
  wire [0:0] direct_interc_89_out;
  wire [0:0] direct_interc_8_out;
  wire [0:0] direct_interc_90_out;
  wire [0:0] direct_interc_91_out;
  wire [0:0] direct_interc_92_out;
  wire [0:0] direct_interc_93_out;
  wire [0:0] direct_interc_94_out;
  wire [0:0] direct_interc_95_out;
  wire [0:0] direct_interc_96_out;
  wire [0:0] direct_interc_97_out;
  wire [0:0] direct_interc_98_out;
  wire [0:0] direct_interc_99_out;
  wire [0:0] direct_interc_9_out;
  wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_0_ccff_tail;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_100_ccff_tail;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_101_ccff_tail;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_102_ccff_tail;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_103_ccff_tail;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_104_ccff_tail;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_105_ccff_tail;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_106_ccff_tail;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_107_ccff_tail;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_108_ccff_tail;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_109_ccff_tail;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_10__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_10__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_10_ccff_tail;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_110_ccff_tail;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_111_ccff_tail;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_112_ccff_tail;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_113_ccff_tail;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_114_ccff_tail;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_115_ccff_tail;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_116_ccff_tail;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_117_ccff_tail;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_118_ccff_tail;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_119_ccff_tail;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_11__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_11__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_11_ccff_tail;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_120_ccff_tail;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_121_ccff_tail;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_122_ccff_tail;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_123_ccff_tail;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_124_ccff_tail;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_125_ccff_tail;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_126_ccff_tail;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_127_ccff_tail;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_128_ccff_tail;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_129_ccff_tail;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_12__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_12_ccff_tail;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_130_ccff_tail;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_131_ccff_tail;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_132_ccff_tail;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_133_ccff_tail;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_134_ccff_tail;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_135_ccff_tail;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_136_ccff_tail;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_137_ccff_tail;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_138_ccff_tail;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_139_ccff_tail;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_13_ccff_tail;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_140_ccff_tail;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_141_ccff_tail;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_142_ccff_tail;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_143_ccff_tail;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_14_ccff_tail;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_15_ccff_tail;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_16_ccff_tail;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_17_ccff_tail;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_18_ccff_tail;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_19_ccff_tail;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_1__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_1__12__undriven_top_width_0_height_0__pin_33_;
  wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_1_ccff_tail;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_20_ccff_tail;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_21_ccff_tail;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_22_ccff_tail;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_23_ccff_tail;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_24_ccff_tail;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_25_ccff_tail;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_26_ccff_tail;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_27_ccff_tail;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_28_ccff_tail;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_29_ccff_tail;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_2__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_2_ccff_tail;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_30_ccff_tail;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_31_ccff_tail;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_32_ccff_tail;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_33_ccff_tail;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_34_ccff_tail;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_35_ccff_tail;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_36_ccff_tail;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_37_ccff_tail;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_38_ccff_tail;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_39_ccff_tail;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_3__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_3_ccff_tail;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_40_ccff_tail;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_41_ccff_tail;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_42_ccff_tail;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_43_ccff_tail;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_44_ccff_tail;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_45_ccff_tail;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_46_ccff_tail;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_47_ccff_tail;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_48_ccff_tail;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_49_ccff_tail;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_4__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_4_ccff_tail;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_50_ccff_tail;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_51_ccff_tail;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_52_ccff_tail;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_53_ccff_tail;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_54_ccff_tail;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_55_ccff_tail;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_56_ccff_tail;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_57_ccff_tail;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_58_ccff_tail;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_59_ccff_tail;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_5__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_5_ccff_tail;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_60_ccff_tail;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_61_ccff_tail;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_62_ccff_tail;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_63_ccff_tail;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_64_ccff_tail;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_65_ccff_tail;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_66_ccff_tail;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_67_ccff_tail;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_68_ccff_tail;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_69_ccff_tail;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_6__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_6__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_6_ccff_tail;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_70_ccff_tail;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_71_ccff_tail;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_72_ccff_tail;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_73_ccff_tail;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_74_ccff_tail;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_75_ccff_tail;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_76_ccff_tail;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_77_ccff_tail;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_78_ccff_tail;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_79_ccff_tail;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_7__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_7_ccff_tail;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_80_ccff_tail;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_81_ccff_tail;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_82_ccff_tail;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_83_ccff_tail;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_84_ccff_tail;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_85_ccff_tail;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_86_ccff_tail;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_87_ccff_tail;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_88_ccff_tail;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_89_ccff_tail;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_8__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_8__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_8_ccff_tail;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_90_ccff_tail;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_91_ccff_tail;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_92_ccff_tail;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_93_ccff_tail;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_94_ccff_tail;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_95_ccff_tail;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_96_ccff_tail;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_97_ccff_tail;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_98_ccff_tail;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_99_ccff_tail;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_9__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_9__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_9_ccff_tail;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_io_bottom_0_ccff_tail;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_10_ccff_tail;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_11_ccff_tail;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_1_ccff_tail;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_2_ccff_tail;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_3_ccff_tail;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_4_ccff_tail;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_5_ccff_tail;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_6_ccff_tail;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_7_ccff_tail;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_8_ccff_tail;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_9_ccff_tail;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_left_0_ccff_tail;
  wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_10_ccff_tail;
  wire [0:0] grid_io_left_10_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_10_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_11_ccff_tail;
  wire [0:0] grid_io_left_11_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_11_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_1_ccff_tail;
  wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_2_ccff_tail;
  wire [0:0] grid_io_left_2_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_2_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_3_ccff_tail;
  wire [0:0] grid_io_left_3_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_3_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_4_ccff_tail;
  wire [0:0] grid_io_left_4_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_4_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_5_ccff_tail;
  wire [0:0] grid_io_left_5_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_5_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_6_ccff_tail;
  wire [0:0] grid_io_left_6_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_6_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_7_ccff_tail;
  wire [0:0] grid_io_left_7_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_7_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_8_ccff_tail;
  wire [0:0] grid_io_left_8_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_8_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_9_ccff_tail;
  wire [0:0] grid_io_left_9_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_9_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_0_ccff_tail;
  wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_10_ccff_tail;
  wire [0:0] grid_io_right_10_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_10_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_11_ccff_tail;
  wire [0:0] grid_io_right_11_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_11_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_1_ccff_tail;
  wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_2_ccff_tail;
  wire [0:0] grid_io_right_2_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_2_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_3_ccff_tail;
  wire [0:0] grid_io_right_3_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_3_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_4_ccff_tail;
  wire [0:0] grid_io_right_4_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_4_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_5_ccff_tail;
  wire [0:0] grid_io_right_5_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_5_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_6_ccff_tail;
  wire [0:0] grid_io_right_6_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_6_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_7_ccff_tail;
  wire [0:0] grid_io_right_7_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_7_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_8_ccff_tail;
  wire [0:0] grid_io_right_8_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_8_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_9_ccff_tail;
  wire [0:0] grid_io_right_9_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_9_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_0_ccff_tail;
  wire [0:0] grid_io_top_10_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_10_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_10_ccff_tail;
  wire [0:0] grid_io_top_11_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_11_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_11_ccff_tail;
  wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_1_ccff_tail;
  wire [0:0] grid_io_top_2_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_2_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_2_ccff_tail;
  wire [0:0] grid_io_top_3_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_3_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_3_ccff_tail;
  wire [0:0] grid_io_top_4_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_4_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_4_ccff_tail;
  wire [0:0] grid_io_top_5_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_5_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_5_ccff_tail;
  wire [0:0] grid_io_top_6_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_6_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_6_ccff_tail;
  wire [0:0] grid_io_top_7_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_7_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_7_ccff_tail;
  wire [0:0] grid_io_top_8_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_8_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_8_ccff_tail;
  wire [0:0] grid_io_top_9_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_9_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_9_ccff_tail;
  wire [0:19] sb_0__0__0_chanx_right_out;
  wire [0:19] sb_0__0__0_chany_top_out;
  wire [0:0] sb_0__12__0_ccff_tail;
  wire [0:19] sb_0__12__0_chanx_right_out;
  wire [0:19] sb_0__12__0_chany_bottom_out;
  wire [0:0] sb_0__1__0_ccff_tail;
  wire [0:19] sb_0__1__0_chanx_right_out;
  wire [0:19] sb_0__1__0_chany_bottom_out;
  wire [0:19] sb_0__1__0_chany_top_out;
  wire [0:0] sb_0__1__10_ccff_tail;
  wire [0:19] sb_0__1__10_chanx_right_out;
  wire [0:19] sb_0__1__10_chany_bottom_out;
  wire [0:19] sb_0__1__10_chany_top_out;
  wire [0:0] sb_0__1__1_ccff_tail;
  wire [0:19] sb_0__1__1_chanx_right_out;
  wire [0:19] sb_0__1__1_chany_bottom_out;
  wire [0:19] sb_0__1__1_chany_top_out;
  wire [0:0] sb_0__1__2_ccff_tail;
  wire [0:19] sb_0__1__2_chanx_right_out;
  wire [0:19] sb_0__1__2_chany_bottom_out;
  wire [0:19] sb_0__1__2_chany_top_out;
  wire [0:0] sb_0__1__3_ccff_tail;
  wire [0:19] sb_0__1__3_chanx_right_out;
  wire [0:19] sb_0__1__3_chany_bottom_out;
  wire [0:19] sb_0__1__3_chany_top_out;
  wire [0:0] sb_0__1__4_ccff_tail;
  wire [0:19] sb_0__1__4_chanx_right_out;
  wire [0:19] sb_0__1__4_chany_bottom_out;
  wire [0:19] sb_0__1__4_chany_top_out;
  wire [0:0] sb_0__1__5_ccff_tail;
  wire [0:19] sb_0__1__5_chanx_right_out;
  wire [0:19] sb_0__1__5_chany_bottom_out;
  wire [0:19] sb_0__1__5_chany_top_out;
  wire [0:0] sb_0__1__6_ccff_tail;
  wire [0:19] sb_0__1__6_chanx_right_out;
  wire [0:19] sb_0__1__6_chany_bottom_out;
  wire [0:19] sb_0__1__6_chany_top_out;
  wire [0:0] sb_0__1__7_ccff_tail;
  wire [0:19] sb_0__1__7_chanx_right_out;
  wire [0:19] sb_0__1__7_chany_bottom_out;
  wire [0:19] sb_0__1__7_chany_top_out;
  wire [0:0] sb_0__1__8_ccff_tail;
  wire [0:19] sb_0__1__8_chanx_right_out;
  wire [0:19] sb_0__1__8_chany_bottom_out;
  wire [0:19] sb_0__1__8_chany_top_out;
  wire [0:0] sb_0__1__9_ccff_tail;
  wire [0:19] sb_0__1__9_chanx_right_out;
  wire [0:19] sb_0__1__9_chany_bottom_out;
  wire [0:19] sb_0__1__9_chany_top_out;
  wire [0:0] sb_12__0__0_ccff_tail;
  wire [0:19] sb_12__0__0_chanx_left_out;
  wire [0:19] sb_12__0__0_chany_top_out;
  wire [0:0] sb_12__12__0_ccff_tail;
  wire [0:19] sb_12__12__0_chanx_left_out;
  wire [0:19] sb_12__12__0_chany_bottom_out;
  wire [0:0] sb_12__1__0_ccff_tail;
  wire [0:19] sb_12__1__0_chanx_left_out;
  wire [0:19] sb_12__1__0_chany_bottom_out;
  wire [0:19] sb_12__1__0_chany_top_out;
  wire [0:0] sb_12__1__10_ccff_tail;
  wire [0:19] sb_12__1__10_chanx_left_out;
  wire [0:19] sb_12__1__10_chany_bottom_out;
  wire [0:19] sb_12__1__10_chany_top_out;
  wire [0:0] sb_12__1__1_ccff_tail;
  wire [0:19] sb_12__1__1_chanx_left_out;
  wire [0:19] sb_12__1__1_chany_bottom_out;
  wire [0:19] sb_12__1__1_chany_top_out;
  wire [0:0] sb_12__1__2_ccff_tail;
  wire [0:19] sb_12__1__2_chanx_left_out;
  wire [0:19] sb_12__1__2_chany_bottom_out;
  wire [0:19] sb_12__1__2_chany_top_out;
  wire [0:0] sb_12__1__3_ccff_tail;
  wire [0:19] sb_12__1__3_chanx_left_out;
  wire [0:19] sb_12__1__3_chany_bottom_out;
  wire [0:19] sb_12__1__3_chany_top_out;
  wire [0:0] sb_12__1__4_ccff_tail;
  wire [0:19] sb_12__1__4_chanx_left_out;
  wire [0:19] sb_12__1__4_chany_bottom_out;
  wire [0:19] sb_12__1__4_chany_top_out;
  wire [0:0] sb_12__1__5_ccff_tail;
  wire [0:19] sb_12__1__5_chanx_left_out;
  wire [0:19] sb_12__1__5_chany_bottom_out;
  wire [0:19] sb_12__1__5_chany_top_out;
  wire [0:0] sb_12__1__6_ccff_tail;
  wire [0:19] sb_12__1__6_chanx_left_out;
  wire [0:19] sb_12__1__6_chany_bottom_out;
  wire [0:19] sb_12__1__6_chany_top_out;
  wire [0:0] sb_12__1__7_ccff_tail;
  wire [0:19] sb_12__1__7_chanx_left_out;
  wire [0:19] sb_12__1__7_chany_bottom_out;
  wire [0:19] sb_12__1__7_chany_top_out;
  wire [0:0] sb_12__1__8_ccff_tail;
  wire [0:19] sb_12__1__8_chanx_left_out;
  wire [0:19] sb_12__1__8_chany_bottom_out;
  wire [0:19] sb_12__1__8_chany_top_out;
  wire [0:0] sb_12__1__9_ccff_tail;
  wire [0:19] sb_12__1__9_chanx_left_out;
  wire [0:19] sb_12__1__9_chany_bottom_out;
  wire [0:19] sb_12__1__9_chany_top_out;
  wire [0:0] sb_1__0__0_ccff_tail;
  wire [0:19] sb_1__0__0_chanx_left_out;
  wire [0:19] sb_1__0__0_chanx_right_out;
  wire [0:19] sb_1__0__0_chany_top_out;
  wire [0:0] sb_1__0__10_ccff_tail;
  wire [0:19] sb_1__0__10_chanx_left_out;
  wire [0:19] sb_1__0__10_chanx_right_out;
  wire [0:19] sb_1__0__10_chany_top_out;
  wire [0:0] sb_1__0__1_ccff_tail;
  wire [0:19] sb_1__0__1_chanx_left_out;
  wire [0:19] sb_1__0__1_chanx_right_out;
  wire [0:19] sb_1__0__1_chany_top_out;
  wire [0:0] sb_1__0__2_ccff_tail;
  wire [0:19] sb_1__0__2_chanx_left_out;
  wire [0:19] sb_1__0__2_chanx_right_out;
  wire [0:19] sb_1__0__2_chany_top_out;
  wire [0:0] sb_1__0__3_ccff_tail;
  wire [0:19] sb_1__0__3_chanx_left_out;
  wire [0:19] sb_1__0__3_chanx_right_out;
  wire [0:19] sb_1__0__3_chany_top_out;
  wire [0:0] sb_1__0__4_ccff_tail;
  wire [0:19] sb_1__0__4_chanx_left_out;
  wire [0:19] sb_1__0__4_chanx_right_out;
  wire [0:19] sb_1__0__4_chany_top_out;
  wire [0:0] sb_1__0__5_ccff_tail;
  wire [0:19] sb_1__0__5_chanx_left_out;
  wire [0:19] sb_1__0__5_chanx_right_out;
  wire [0:19] sb_1__0__5_chany_top_out;
  wire [0:0] sb_1__0__6_ccff_tail;
  wire [0:19] sb_1__0__6_chanx_left_out;
  wire [0:19] sb_1__0__6_chanx_right_out;
  wire [0:19] sb_1__0__6_chany_top_out;
  wire [0:0] sb_1__0__7_ccff_tail;
  wire [0:19] sb_1__0__7_chanx_left_out;
  wire [0:19] sb_1__0__7_chanx_right_out;
  wire [0:19] sb_1__0__7_chany_top_out;
  wire [0:0] sb_1__0__8_ccff_tail;
  wire [0:19] sb_1__0__8_chanx_left_out;
  wire [0:19] sb_1__0__8_chanx_right_out;
  wire [0:19] sb_1__0__8_chany_top_out;
  wire [0:0] sb_1__0__9_ccff_tail;
  wire [0:19] sb_1__0__9_chanx_left_out;
  wire [0:19] sb_1__0__9_chanx_right_out;
  wire [0:19] sb_1__0__9_chany_top_out;
  wire [0:0] sb_1__12__0_ccff_tail;
  wire [0:19] sb_1__12__0_chanx_left_out;
  wire [0:19] sb_1__12__0_chanx_right_out;
  wire [0:19] sb_1__12__0_chany_bottom_out;
  wire [0:0] sb_1__12__10_ccff_tail;
  wire [0:19] sb_1__12__10_chanx_left_out;
  wire [0:19] sb_1__12__10_chanx_right_out;
  wire [0:19] sb_1__12__10_chany_bottom_out;
  wire [0:0] sb_1__12__1_ccff_tail;
  wire [0:19] sb_1__12__1_chanx_left_out;
  wire [0:19] sb_1__12__1_chanx_right_out;
  wire [0:19] sb_1__12__1_chany_bottom_out;
  wire [0:0] sb_1__12__2_ccff_tail;
  wire [0:19] sb_1__12__2_chanx_left_out;
  wire [0:19] sb_1__12__2_chanx_right_out;
  wire [0:19] sb_1__12__2_chany_bottom_out;
  wire [0:0] sb_1__12__3_ccff_tail;
  wire [0:19] sb_1__12__3_chanx_left_out;
  wire [0:19] sb_1__12__3_chanx_right_out;
  wire [0:19] sb_1__12__3_chany_bottom_out;
  wire [0:0] sb_1__12__4_ccff_tail;
  wire [0:19] sb_1__12__4_chanx_left_out;
  wire [0:19] sb_1__12__4_chanx_right_out;
  wire [0:19] sb_1__12__4_chany_bottom_out;
  wire [0:0] sb_1__12__5_ccff_tail;
  wire [0:19] sb_1__12__5_chanx_left_out;
  wire [0:19] sb_1__12__5_chanx_right_out;
  wire [0:19] sb_1__12__5_chany_bottom_out;
  wire [0:0] sb_1__12__6_ccff_tail;
  wire [0:19] sb_1__12__6_chanx_left_out;
  wire [0:19] sb_1__12__6_chanx_right_out;
  wire [0:19] sb_1__12__6_chany_bottom_out;
  wire [0:0] sb_1__12__7_ccff_tail;
  wire [0:19] sb_1__12__7_chanx_left_out;
  wire [0:19] sb_1__12__7_chanx_right_out;
  wire [0:19] sb_1__12__7_chany_bottom_out;
  wire [0:0] sb_1__12__8_ccff_tail;
  wire [0:19] sb_1__12__8_chanx_left_out;
  wire [0:19] sb_1__12__8_chanx_right_out;
  wire [0:19] sb_1__12__8_chany_bottom_out;
  wire [0:0] sb_1__12__9_ccff_tail;
  wire [0:19] sb_1__12__9_chanx_left_out;
  wire [0:19] sb_1__12__9_chanx_right_out;
  wire [0:19] sb_1__12__9_chany_bottom_out;
  wire [0:0] sb_1__1__0_ccff_tail;
  wire [0:19] sb_1__1__0_chanx_left_out;
  wire [0:19] sb_1__1__0_chanx_right_out;
  wire [0:19] sb_1__1__0_chany_bottom_out;
  wire [0:19] sb_1__1__0_chany_top_out;
  wire [0:0] sb_1__1__100_ccff_tail;
  wire [0:19] sb_1__1__100_chanx_left_out;
  wire [0:19] sb_1__1__100_chanx_right_out;
  wire [0:19] sb_1__1__100_chany_bottom_out;
  wire [0:19] sb_1__1__100_chany_top_out;
  wire [0:0] sb_1__1__101_ccff_tail;
  wire [0:19] sb_1__1__101_chanx_left_out;
  wire [0:19] sb_1__1__101_chanx_right_out;
  wire [0:19] sb_1__1__101_chany_bottom_out;
  wire [0:19] sb_1__1__101_chany_top_out;
  wire [0:0] sb_1__1__102_ccff_tail;
  wire [0:19] sb_1__1__102_chanx_left_out;
  wire [0:19] sb_1__1__102_chanx_right_out;
  wire [0:19] sb_1__1__102_chany_bottom_out;
  wire [0:19] sb_1__1__102_chany_top_out;
  wire [0:0] sb_1__1__103_ccff_tail;
  wire [0:19] sb_1__1__103_chanx_left_out;
  wire [0:19] sb_1__1__103_chanx_right_out;
  wire [0:19] sb_1__1__103_chany_bottom_out;
  wire [0:19] sb_1__1__103_chany_top_out;
  wire [0:0] sb_1__1__104_ccff_tail;
  wire [0:19] sb_1__1__104_chanx_left_out;
  wire [0:19] sb_1__1__104_chanx_right_out;
  wire [0:19] sb_1__1__104_chany_bottom_out;
  wire [0:19] sb_1__1__104_chany_top_out;
  wire [0:0] sb_1__1__105_ccff_tail;
  wire [0:19] sb_1__1__105_chanx_left_out;
  wire [0:19] sb_1__1__105_chanx_right_out;
  wire [0:19] sb_1__1__105_chany_bottom_out;
  wire [0:19] sb_1__1__105_chany_top_out;
  wire [0:0] sb_1__1__106_ccff_tail;
  wire [0:19] sb_1__1__106_chanx_left_out;
  wire [0:19] sb_1__1__106_chanx_right_out;
  wire [0:19] sb_1__1__106_chany_bottom_out;
  wire [0:19] sb_1__1__106_chany_top_out;
  wire [0:0] sb_1__1__107_ccff_tail;
  wire [0:19] sb_1__1__107_chanx_left_out;
  wire [0:19] sb_1__1__107_chanx_right_out;
  wire [0:19] sb_1__1__107_chany_bottom_out;
  wire [0:19] sb_1__1__107_chany_top_out;
  wire [0:0] sb_1__1__108_ccff_tail;
  wire [0:19] sb_1__1__108_chanx_left_out;
  wire [0:19] sb_1__1__108_chanx_right_out;
  wire [0:19] sb_1__1__108_chany_bottom_out;
  wire [0:19] sb_1__1__108_chany_top_out;
  wire [0:0] sb_1__1__109_ccff_tail;
  wire [0:19] sb_1__1__109_chanx_left_out;
  wire [0:19] sb_1__1__109_chanx_right_out;
  wire [0:19] sb_1__1__109_chany_bottom_out;
  wire [0:19] sb_1__1__109_chany_top_out;
  wire [0:0] sb_1__1__10_ccff_tail;
  wire [0:19] sb_1__1__10_chanx_left_out;
  wire [0:19] sb_1__1__10_chanx_right_out;
  wire [0:19] sb_1__1__10_chany_bottom_out;
  wire [0:19] sb_1__1__10_chany_top_out;
  wire [0:0] sb_1__1__110_ccff_tail;
  wire [0:19] sb_1__1__110_chanx_left_out;
  wire [0:19] sb_1__1__110_chanx_right_out;
  wire [0:19] sb_1__1__110_chany_bottom_out;
  wire [0:19] sb_1__1__110_chany_top_out;
  wire [0:0] sb_1__1__111_ccff_tail;
  wire [0:19] sb_1__1__111_chanx_left_out;
  wire [0:19] sb_1__1__111_chanx_right_out;
  wire [0:19] sb_1__1__111_chany_bottom_out;
  wire [0:19] sb_1__1__111_chany_top_out;
  wire [0:0] sb_1__1__112_ccff_tail;
  wire [0:19] sb_1__1__112_chanx_left_out;
  wire [0:19] sb_1__1__112_chanx_right_out;
  wire [0:19] sb_1__1__112_chany_bottom_out;
  wire [0:19] sb_1__1__112_chany_top_out;
  wire [0:0] sb_1__1__113_ccff_tail;
  wire [0:19] sb_1__1__113_chanx_left_out;
  wire [0:19] sb_1__1__113_chanx_right_out;
  wire [0:19] sb_1__1__113_chany_bottom_out;
  wire [0:19] sb_1__1__113_chany_top_out;
  wire [0:0] sb_1__1__114_ccff_tail;
  wire [0:19] sb_1__1__114_chanx_left_out;
  wire [0:19] sb_1__1__114_chanx_right_out;
  wire [0:19] sb_1__1__114_chany_bottom_out;
  wire [0:19] sb_1__1__114_chany_top_out;
  wire [0:0] sb_1__1__115_ccff_tail;
  wire [0:19] sb_1__1__115_chanx_left_out;
  wire [0:19] sb_1__1__115_chanx_right_out;
  wire [0:19] sb_1__1__115_chany_bottom_out;
  wire [0:19] sb_1__1__115_chany_top_out;
  wire [0:0] sb_1__1__116_ccff_tail;
  wire [0:19] sb_1__1__116_chanx_left_out;
  wire [0:19] sb_1__1__116_chanx_right_out;
  wire [0:19] sb_1__1__116_chany_bottom_out;
  wire [0:19] sb_1__1__116_chany_top_out;
  wire [0:0] sb_1__1__117_ccff_tail;
  wire [0:19] sb_1__1__117_chanx_left_out;
  wire [0:19] sb_1__1__117_chanx_right_out;
  wire [0:19] sb_1__1__117_chany_bottom_out;
  wire [0:19] sb_1__1__117_chany_top_out;
  wire [0:0] sb_1__1__118_ccff_tail;
  wire [0:19] sb_1__1__118_chanx_left_out;
  wire [0:19] sb_1__1__118_chanx_right_out;
  wire [0:19] sb_1__1__118_chany_bottom_out;
  wire [0:19] sb_1__1__118_chany_top_out;
  wire [0:0] sb_1__1__119_ccff_tail;
  wire [0:19] sb_1__1__119_chanx_left_out;
  wire [0:19] sb_1__1__119_chanx_right_out;
  wire [0:19] sb_1__1__119_chany_bottom_out;
  wire [0:19] sb_1__1__119_chany_top_out;
  wire [0:0] sb_1__1__11_ccff_tail;
  wire [0:19] sb_1__1__11_chanx_left_out;
  wire [0:19] sb_1__1__11_chanx_right_out;
  wire [0:19] sb_1__1__11_chany_bottom_out;
  wire [0:19] sb_1__1__11_chany_top_out;
  wire [0:0] sb_1__1__120_ccff_tail;
  wire [0:19] sb_1__1__120_chanx_left_out;
  wire [0:19] sb_1__1__120_chanx_right_out;
  wire [0:19] sb_1__1__120_chany_bottom_out;
  wire [0:19] sb_1__1__120_chany_top_out;
  wire [0:0] sb_1__1__12_ccff_tail;
  wire [0:19] sb_1__1__12_chanx_left_out;
  wire [0:19] sb_1__1__12_chanx_right_out;
  wire [0:19] sb_1__1__12_chany_bottom_out;
  wire [0:19] sb_1__1__12_chany_top_out;
  wire [0:0] sb_1__1__13_ccff_tail;
  wire [0:19] sb_1__1__13_chanx_left_out;
  wire [0:19] sb_1__1__13_chanx_right_out;
  wire [0:19] sb_1__1__13_chany_bottom_out;
  wire [0:19] sb_1__1__13_chany_top_out;
  wire [0:0] sb_1__1__14_ccff_tail;
  wire [0:19] sb_1__1__14_chanx_left_out;
  wire [0:19] sb_1__1__14_chanx_right_out;
  wire [0:19] sb_1__1__14_chany_bottom_out;
  wire [0:19] sb_1__1__14_chany_top_out;
  wire [0:0] sb_1__1__15_ccff_tail;
  wire [0:19] sb_1__1__15_chanx_left_out;
  wire [0:19] sb_1__1__15_chanx_right_out;
  wire [0:19] sb_1__1__15_chany_bottom_out;
  wire [0:19] sb_1__1__15_chany_top_out;
  wire [0:0] sb_1__1__16_ccff_tail;
  wire [0:19] sb_1__1__16_chanx_left_out;
  wire [0:19] sb_1__1__16_chanx_right_out;
  wire [0:19] sb_1__1__16_chany_bottom_out;
  wire [0:19] sb_1__1__16_chany_top_out;
  wire [0:0] sb_1__1__17_ccff_tail;
  wire [0:19] sb_1__1__17_chanx_left_out;
  wire [0:19] sb_1__1__17_chanx_right_out;
  wire [0:19] sb_1__1__17_chany_bottom_out;
  wire [0:19] sb_1__1__17_chany_top_out;
  wire [0:0] sb_1__1__18_ccff_tail;
  wire [0:19] sb_1__1__18_chanx_left_out;
  wire [0:19] sb_1__1__18_chanx_right_out;
  wire [0:19] sb_1__1__18_chany_bottom_out;
  wire [0:19] sb_1__1__18_chany_top_out;
  wire [0:0] sb_1__1__19_ccff_tail;
  wire [0:19] sb_1__1__19_chanx_left_out;
  wire [0:19] sb_1__1__19_chanx_right_out;
  wire [0:19] sb_1__1__19_chany_bottom_out;
  wire [0:19] sb_1__1__19_chany_top_out;
  wire [0:0] sb_1__1__1_ccff_tail;
  wire [0:19] sb_1__1__1_chanx_left_out;
  wire [0:19] sb_1__1__1_chanx_right_out;
  wire [0:19] sb_1__1__1_chany_bottom_out;
  wire [0:19] sb_1__1__1_chany_top_out;
  wire [0:0] sb_1__1__20_ccff_tail;
  wire [0:19] sb_1__1__20_chanx_left_out;
  wire [0:19] sb_1__1__20_chanx_right_out;
  wire [0:19] sb_1__1__20_chany_bottom_out;
  wire [0:19] sb_1__1__20_chany_top_out;
  wire [0:0] sb_1__1__21_ccff_tail;
  wire [0:19] sb_1__1__21_chanx_left_out;
  wire [0:19] sb_1__1__21_chanx_right_out;
  wire [0:19] sb_1__1__21_chany_bottom_out;
  wire [0:19] sb_1__1__21_chany_top_out;
  wire [0:0] sb_1__1__22_ccff_tail;
  wire [0:19] sb_1__1__22_chanx_left_out;
  wire [0:19] sb_1__1__22_chanx_right_out;
  wire [0:19] sb_1__1__22_chany_bottom_out;
  wire [0:19] sb_1__1__22_chany_top_out;
  wire [0:0] sb_1__1__23_ccff_tail;
  wire [0:19] sb_1__1__23_chanx_left_out;
  wire [0:19] sb_1__1__23_chanx_right_out;
  wire [0:19] sb_1__1__23_chany_bottom_out;
  wire [0:19] sb_1__1__23_chany_top_out;
  wire [0:0] sb_1__1__24_ccff_tail;
  wire [0:19] sb_1__1__24_chanx_left_out;
  wire [0:19] sb_1__1__24_chanx_right_out;
  wire [0:19] sb_1__1__24_chany_bottom_out;
  wire [0:19] sb_1__1__24_chany_top_out;
  wire [0:0] sb_1__1__25_ccff_tail;
  wire [0:19] sb_1__1__25_chanx_left_out;
  wire [0:19] sb_1__1__25_chanx_right_out;
  wire [0:19] sb_1__1__25_chany_bottom_out;
  wire [0:19] sb_1__1__25_chany_top_out;
  wire [0:0] sb_1__1__26_ccff_tail;
  wire [0:19] sb_1__1__26_chanx_left_out;
  wire [0:19] sb_1__1__26_chanx_right_out;
  wire [0:19] sb_1__1__26_chany_bottom_out;
  wire [0:19] sb_1__1__26_chany_top_out;
  wire [0:0] sb_1__1__27_ccff_tail;
  wire [0:19] sb_1__1__27_chanx_left_out;
  wire [0:19] sb_1__1__27_chanx_right_out;
  wire [0:19] sb_1__1__27_chany_bottom_out;
  wire [0:19] sb_1__1__27_chany_top_out;
  wire [0:0] sb_1__1__28_ccff_tail;
  wire [0:19] sb_1__1__28_chanx_left_out;
  wire [0:19] sb_1__1__28_chanx_right_out;
  wire [0:19] sb_1__1__28_chany_bottom_out;
  wire [0:19] sb_1__1__28_chany_top_out;
  wire [0:0] sb_1__1__29_ccff_tail;
  wire [0:19] sb_1__1__29_chanx_left_out;
  wire [0:19] sb_1__1__29_chanx_right_out;
  wire [0:19] sb_1__1__29_chany_bottom_out;
  wire [0:19] sb_1__1__29_chany_top_out;
  wire [0:0] sb_1__1__2_ccff_tail;
  wire [0:19] sb_1__1__2_chanx_left_out;
  wire [0:19] sb_1__1__2_chanx_right_out;
  wire [0:19] sb_1__1__2_chany_bottom_out;
  wire [0:19] sb_1__1__2_chany_top_out;
  wire [0:0] sb_1__1__30_ccff_tail;
  wire [0:19] sb_1__1__30_chanx_left_out;
  wire [0:19] sb_1__1__30_chanx_right_out;
  wire [0:19] sb_1__1__30_chany_bottom_out;
  wire [0:19] sb_1__1__30_chany_top_out;
  wire [0:0] sb_1__1__31_ccff_tail;
  wire [0:19] sb_1__1__31_chanx_left_out;
  wire [0:19] sb_1__1__31_chanx_right_out;
  wire [0:19] sb_1__1__31_chany_bottom_out;
  wire [0:19] sb_1__1__31_chany_top_out;
  wire [0:0] sb_1__1__32_ccff_tail;
  wire [0:19] sb_1__1__32_chanx_left_out;
  wire [0:19] sb_1__1__32_chanx_right_out;
  wire [0:19] sb_1__1__32_chany_bottom_out;
  wire [0:19] sb_1__1__32_chany_top_out;
  wire [0:0] sb_1__1__33_ccff_tail;
  wire [0:19] sb_1__1__33_chanx_left_out;
  wire [0:19] sb_1__1__33_chanx_right_out;
  wire [0:19] sb_1__1__33_chany_bottom_out;
  wire [0:19] sb_1__1__33_chany_top_out;
  wire [0:0] sb_1__1__34_ccff_tail;
  wire [0:19] sb_1__1__34_chanx_left_out;
  wire [0:19] sb_1__1__34_chanx_right_out;
  wire [0:19] sb_1__1__34_chany_bottom_out;
  wire [0:19] sb_1__1__34_chany_top_out;
  wire [0:0] sb_1__1__35_ccff_tail;
  wire [0:19] sb_1__1__35_chanx_left_out;
  wire [0:19] sb_1__1__35_chanx_right_out;
  wire [0:19] sb_1__1__35_chany_bottom_out;
  wire [0:19] sb_1__1__35_chany_top_out;
  wire [0:0] sb_1__1__36_ccff_tail;
  wire [0:19] sb_1__1__36_chanx_left_out;
  wire [0:19] sb_1__1__36_chanx_right_out;
  wire [0:19] sb_1__1__36_chany_bottom_out;
  wire [0:19] sb_1__1__36_chany_top_out;
  wire [0:0] sb_1__1__37_ccff_tail;
  wire [0:19] sb_1__1__37_chanx_left_out;
  wire [0:19] sb_1__1__37_chanx_right_out;
  wire [0:19] sb_1__1__37_chany_bottom_out;
  wire [0:19] sb_1__1__37_chany_top_out;
  wire [0:0] sb_1__1__38_ccff_tail;
  wire [0:19] sb_1__1__38_chanx_left_out;
  wire [0:19] sb_1__1__38_chanx_right_out;
  wire [0:19] sb_1__1__38_chany_bottom_out;
  wire [0:19] sb_1__1__38_chany_top_out;
  wire [0:0] sb_1__1__39_ccff_tail;
  wire [0:19] sb_1__1__39_chanx_left_out;
  wire [0:19] sb_1__1__39_chanx_right_out;
  wire [0:19] sb_1__1__39_chany_bottom_out;
  wire [0:19] sb_1__1__39_chany_top_out;
  wire [0:0] sb_1__1__3_ccff_tail;
  wire [0:19] sb_1__1__3_chanx_left_out;
  wire [0:19] sb_1__1__3_chanx_right_out;
  wire [0:19] sb_1__1__3_chany_bottom_out;
  wire [0:19] sb_1__1__3_chany_top_out;
  wire [0:0] sb_1__1__40_ccff_tail;
  wire [0:19] sb_1__1__40_chanx_left_out;
  wire [0:19] sb_1__1__40_chanx_right_out;
  wire [0:19] sb_1__1__40_chany_bottom_out;
  wire [0:19] sb_1__1__40_chany_top_out;
  wire [0:0] sb_1__1__41_ccff_tail;
  wire [0:19] sb_1__1__41_chanx_left_out;
  wire [0:19] sb_1__1__41_chanx_right_out;
  wire [0:19] sb_1__1__41_chany_bottom_out;
  wire [0:19] sb_1__1__41_chany_top_out;
  wire [0:0] sb_1__1__42_ccff_tail;
  wire [0:19] sb_1__1__42_chanx_left_out;
  wire [0:19] sb_1__1__42_chanx_right_out;
  wire [0:19] sb_1__1__42_chany_bottom_out;
  wire [0:19] sb_1__1__42_chany_top_out;
  wire [0:0] sb_1__1__43_ccff_tail;
  wire [0:19] sb_1__1__43_chanx_left_out;
  wire [0:19] sb_1__1__43_chanx_right_out;
  wire [0:19] sb_1__1__43_chany_bottom_out;
  wire [0:19] sb_1__1__43_chany_top_out;
  wire [0:0] sb_1__1__44_ccff_tail;
  wire [0:19] sb_1__1__44_chanx_left_out;
  wire [0:19] sb_1__1__44_chanx_right_out;
  wire [0:19] sb_1__1__44_chany_bottom_out;
  wire [0:19] sb_1__1__44_chany_top_out;
  wire [0:0] sb_1__1__45_ccff_tail;
  wire [0:19] sb_1__1__45_chanx_left_out;
  wire [0:19] sb_1__1__45_chanx_right_out;
  wire [0:19] sb_1__1__45_chany_bottom_out;
  wire [0:19] sb_1__1__45_chany_top_out;
  wire [0:0] sb_1__1__46_ccff_tail;
  wire [0:19] sb_1__1__46_chanx_left_out;
  wire [0:19] sb_1__1__46_chanx_right_out;
  wire [0:19] sb_1__1__46_chany_bottom_out;
  wire [0:19] sb_1__1__46_chany_top_out;
  wire [0:0] sb_1__1__47_ccff_tail;
  wire [0:19] sb_1__1__47_chanx_left_out;
  wire [0:19] sb_1__1__47_chanx_right_out;
  wire [0:19] sb_1__1__47_chany_bottom_out;
  wire [0:19] sb_1__1__47_chany_top_out;
  wire [0:0] sb_1__1__48_ccff_tail;
  wire [0:19] sb_1__1__48_chanx_left_out;
  wire [0:19] sb_1__1__48_chanx_right_out;
  wire [0:19] sb_1__1__48_chany_bottom_out;
  wire [0:19] sb_1__1__48_chany_top_out;
  wire [0:0] sb_1__1__49_ccff_tail;
  wire [0:19] sb_1__1__49_chanx_left_out;
  wire [0:19] sb_1__1__49_chanx_right_out;
  wire [0:19] sb_1__1__49_chany_bottom_out;
  wire [0:19] sb_1__1__49_chany_top_out;
  wire [0:0] sb_1__1__4_ccff_tail;
  wire [0:19] sb_1__1__4_chanx_left_out;
  wire [0:19] sb_1__1__4_chanx_right_out;
  wire [0:19] sb_1__1__4_chany_bottom_out;
  wire [0:19] sb_1__1__4_chany_top_out;
  wire [0:0] sb_1__1__50_ccff_tail;
  wire [0:19] sb_1__1__50_chanx_left_out;
  wire [0:19] sb_1__1__50_chanx_right_out;
  wire [0:19] sb_1__1__50_chany_bottom_out;
  wire [0:19] sb_1__1__50_chany_top_out;
  wire [0:0] sb_1__1__51_ccff_tail;
  wire [0:19] sb_1__1__51_chanx_left_out;
  wire [0:19] sb_1__1__51_chanx_right_out;
  wire [0:19] sb_1__1__51_chany_bottom_out;
  wire [0:19] sb_1__1__51_chany_top_out;
  wire [0:0] sb_1__1__52_ccff_tail;
  wire [0:19] sb_1__1__52_chanx_left_out;
  wire [0:19] sb_1__1__52_chanx_right_out;
  wire [0:19] sb_1__1__52_chany_bottom_out;
  wire [0:19] sb_1__1__52_chany_top_out;
  wire [0:0] sb_1__1__53_ccff_tail;
  wire [0:19] sb_1__1__53_chanx_left_out;
  wire [0:19] sb_1__1__53_chanx_right_out;
  wire [0:19] sb_1__1__53_chany_bottom_out;
  wire [0:19] sb_1__1__53_chany_top_out;
  wire [0:0] sb_1__1__54_ccff_tail;
  wire [0:19] sb_1__1__54_chanx_left_out;
  wire [0:19] sb_1__1__54_chanx_right_out;
  wire [0:19] sb_1__1__54_chany_bottom_out;
  wire [0:19] sb_1__1__54_chany_top_out;
  wire [0:0] sb_1__1__55_ccff_tail;
  wire [0:19] sb_1__1__55_chanx_left_out;
  wire [0:19] sb_1__1__55_chanx_right_out;
  wire [0:19] sb_1__1__55_chany_bottom_out;
  wire [0:19] sb_1__1__55_chany_top_out;
  wire [0:0] sb_1__1__56_ccff_tail;
  wire [0:19] sb_1__1__56_chanx_left_out;
  wire [0:19] sb_1__1__56_chanx_right_out;
  wire [0:19] sb_1__1__56_chany_bottom_out;
  wire [0:19] sb_1__1__56_chany_top_out;
  wire [0:0] sb_1__1__57_ccff_tail;
  wire [0:19] sb_1__1__57_chanx_left_out;
  wire [0:19] sb_1__1__57_chanx_right_out;
  wire [0:19] sb_1__1__57_chany_bottom_out;
  wire [0:19] sb_1__1__57_chany_top_out;
  wire [0:0] sb_1__1__58_ccff_tail;
  wire [0:19] sb_1__1__58_chanx_left_out;
  wire [0:19] sb_1__1__58_chanx_right_out;
  wire [0:19] sb_1__1__58_chany_bottom_out;
  wire [0:19] sb_1__1__58_chany_top_out;
  wire [0:0] sb_1__1__59_ccff_tail;
  wire [0:19] sb_1__1__59_chanx_left_out;
  wire [0:19] sb_1__1__59_chanx_right_out;
  wire [0:19] sb_1__1__59_chany_bottom_out;
  wire [0:19] sb_1__1__59_chany_top_out;
  wire [0:0] sb_1__1__5_ccff_tail;
  wire [0:19] sb_1__1__5_chanx_left_out;
  wire [0:19] sb_1__1__5_chanx_right_out;
  wire [0:19] sb_1__1__5_chany_bottom_out;
  wire [0:19] sb_1__1__5_chany_top_out;
  wire [0:0] sb_1__1__60_ccff_tail;
  wire [0:19] sb_1__1__60_chanx_left_out;
  wire [0:19] sb_1__1__60_chanx_right_out;
  wire [0:19] sb_1__1__60_chany_bottom_out;
  wire [0:19] sb_1__1__60_chany_top_out;
  wire [0:0] sb_1__1__61_ccff_tail;
  wire [0:19] sb_1__1__61_chanx_left_out;
  wire [0:19] sb_1__1__61_chanx_right_out;
  wire [0:19] sb_1__1__61_chany_bottom_out;
  wire [0:19] sb_1__1__61_chany_top_out;
  wire [0:0] sb_1__1__62_ccff_tail;
  wire [0:19] sb_1__1__62_chanx_left_out;
  wire [0:19] sb_1__1__62_chanx_right_out;
  wire [0:19] sb_1__1__62_chany_bottom_out;
  wire [0:19] sb_1__1__62_chany_top_out;
  wire [0:0] sb_1__1__63_ccff_tail;
  wire [0:19] sb_1__1__63_chanx_left_out;
  wire [0:19] sb_1__1__63_chanx_right_out;
  wire [0:19] sb_1__1__63_chany_bottom_out;
  wire [0:19] sb_1__1__63_chany_top_out;
  wire [0:0] sb_1__1__64_ccff_tail;
  wire [0:19] sb_1__1__64_chanx_left_out;
  wire [0:19] sb_1__1__64_chanx_right_out;
  wire [0:19] sb_1__1__64_chany_bottom_out;
  wire [0:19] sb_1__1__64_chany_top_out;
  wire [0:0] sb_1__1__65_ccff_tail;
  wire [0:19] sb_1__1__65_chanx_left_out;
  wire [0:19] sb_1__1__65_chanx_right_out;
  wire [0:19] sb_1__1__65_chany_bottom_out;
  wire [0:19] sb_1__1__65_chany_top_out;
  wire [0:0] sb_1__1__66_ccff_tail;
  wire [0:19] sb_1__1__66_chanx_left_out;
  wire [0:19] sb_1__1__66_chanx_right_out;
  wire [0:19] sb_1__1__66_chany_bottom_out;
  wire [0:19] sb_1__1__66_chany_top_out;
  wire [0:0] sb_1__1__67_ccff_tail;
  wire [0:19] sb_1__1__67_chanx_left_out;
  wire [0:19] sb_1__1__67_chanx_right_out;
  wire [0:19] sb_1__1__67_chany_bottom_out;
  wire [0:19] sb_1__1__67_chany_top_out;
  wire [0:0] sb_1__1__68_ccff_tail;
  wire [0:19] sb_1__1__68_chanx_left_out;
  wire [0:19] sb_1__1__68_chanx_right_out;
  wire [0:19] sb_1__1__68_chany_bottom_out;
  wire [0:19] sb_1__1__68_chany_top_out;
  wire [0:0] sb_1__1__69_ccff_tail;
  wire [0:19] sb_1__1__69_chanx_left_out;
  wire [0:19] sb_1__1__69_chanx_right_out;
  wire [0:19] sb_1__1__69_chany_bottom_out;
  wire [0:19] sb_1__1__69_chany_top_out;
  wire [0:0] sb_1__1__6_ccff_tail;
  wire [0:19] sb_1__1__6_chanx_left_out;
  wire [0:19] sb_1__1__6_chanx_right_out;
  wire [0:19] sb_1__1__6_chany_bottom_out;
  wire [0:19] sb_1__1__6_chany_top_out;
  wire [0:0] sb_1__1__70_ccff_tail;
  wire [0:19] sb_1__1__70_chanx_left_out;
  wire [0:19] sb_1__1__70_chanx_right_out;
  wire [0:19] sb_1__1__70_chany_bottom_out;
  wire [0:19] sb_1__1__70_chany_top_out;
  wire [0:0] sb_1__1__71_ccff_tail;
  wire [0:19] sb_1__1__71_chanx_left_out;
  wire [0:19] sb_1__1__71_chanx_right_out;
  wire [0:19] sb_1__1__71_chany_bottom_out;
  wire [0:19] sb_1__1__71_chany_top_out;
  wire [0:0] sb_1__1__72_ccff_tail;
  wire [0:19] sb_1__1__72_chanx_left_out;
  wire [0:19] sb_1__1__72_chanx_right_out;
  wire [0:19] sb_1__1__72_chany_bottom_out;
  wire [0:19] sb_1__1__72_chany_top_out;
  wire [0:0] sb_1__1__73_ccff_tail;
  wire [0:19] sb_1__1__73_chanx_left_out;
  wire [0:19] sb_1__1__73_chanx_right_out;
  wire [0:19] sb_1__1__73_chany_bottom_out;
  wire [0:19] sb_1__1__73_chany_top_out;
  wire [0:0] sb_1__1__74_ccff_tail;
  wire [0:19] sb_1__1__74_chanx_left_out;
  wire [0:19] sb_1__1__74_chanx_right_out;
  wire [0:19] sb_1__1__74_chany_bottom_out;
  wire [0:19] sb_1__1__74_chany_top_out;
  wire [0:0] sb_1__1__75_ccff_tail;
  wire [0:19] sb_1__1__75_chanx_left_out;
  wire [0:19] sb_1__1__75_chanx_right_out;
  wire [0:19] sb_1__1__75_chany_bottom_out;
  wire [0:19] sb_1__1__75_chany_top_out;
  wire [0:0] sb_1__1__76_ccff_tail;
  wire [0:19] sb_1__1__76_chanx_left_out;
  wire [0:19] sb_1__1__76_chanx_right_out;
  wire [0:19] sb_1__1__76_chany_bottom_out;
  wire [0:19] sb_1__1__76_chany_top_out;
  wire [0:0] sb_1__1__77_ccff_tail;
  wire [0:19] sb_1__1__77_chanx_left_out;
  wire [0:19] sb_1__1__77_chanx_right_out;
  wire [0:19] sb_1__1__77_chany_bottom_out;
  wire [0:19] sb_1__1__77_chany_top_out;
  wire [0:0] sb_1__1__78_ccff_tail;
  wire [0:19] sb_1__1__78_chanx_left_out;
  wire [0:19] sb_1__1__78_chanx_right_out;
  wire [0:19] sb_1__1__78_chany_bottom_out;
  wire [0:19] sb_1__1__78_chany_top_out;
  wire [0:0] sb_1__1__79_ccff_tail;
  wire [0:19] sb_1__1__79_chanx_left_out;
  wire [0:19] sb_1__1__79_chanx_right_out;
  wire [0:19] sb_1__1__79_chany_bottom_out;
  wire [0:19] sb_1__1__79_chany_top_out;
  wire [0:0] sb_1__1__7_ccff_tail;
  wire [0:19] sb_1__1__7_chanx_left_out;
  wire [0:19] sb_1__1__7_chanx_right_out;
  wire [0:19] sb_1__1__7_chany_bottom_out;
  wire [0:19] sb_1__1__7_chany_top_out;
  wire [0:0] sb_1__1__80_ccff_tail;
  wire [0:19] sb_1__1__80_chanx_left_out;
  wire [0:19] sb_1__1__80_chanx_right_out;
  wire [0:19] sb_1__1__80_chany_bottom_out;
  wire [0:19] sb_1__1__80_chany_top_out;
  wire [0:0] sb_1__1__81_ccff_tail;
  wire [0:19] sb_1__1__81_chanx_left_out;
  wire [0:19] sb_1__1__81_chanx_right_out;
  wire [0:19] sb_1__1__81_chany_bottom_out;
  wire [0:19] sb_1__1__81_chany_top_out;
  wire [0:0] sb_1__1__82_ccff_tail;
  wire [0:19] sb_1__1__82_chanx_left_out;
  wire [0:19] sb_1__1__82_chanx_right_out;
  wire [0:19] sb_1__1__82_chany_bottom_out;
  wire [0:19] sb_1__1__82_chany_top_out;
  wire [0:0] sb_1__1__83_ccff_tail;
  wire [0:19] sb_1__1__83_chanx_left_out;
  wire [0:19] sb_1__1__83_chanx_right_out;
  wire [0:19] sb_1__1__83_chany_bottom_out;
  wire [0:19] sb_1__1__83_chany_top_out;
  wire [0:0] sb_1__1__84_ccff_tail;
  wire [0:19] sb_1__1__84_chanx_left_out;
  wire [0:19] sb_1__1__84_chanx_right_out;
  wire [0:19] sb_1__1__84_chany_bottom_out;
  wire [0:19] sb_1__1__84_chany_top_out;
  wire [0:0] sb_1__1__85_ccff_tail;
  wire [0:19] sb_1__1__85_chanx_left_out;
  wire [0:19] sb_1__1__85_chanx_right_out;
  wire [0:19] sb_1__1__85_chany_bottom_out;
  wire [0:19] sb_1__1__85_chany_top_out;
  wire [0:0] sb_1__1__86_ccff_tail;
  wire [0:19] sb_1__1__86_chanx_left_out;
  wire [0:19] sb_1__1__86_chanx_right_out;
  wire [0:19] sb_1__1__86_chany_bottom_out;
  wire [0:19] sb_1__1__86_chany_top_out;
  wire [0:0] sb_1__1__87_ccff_tail;
  wire [0:19] sb_1__1__87_chanx_left_out;
  wire [0:19] sb_1__1__87_chanx_right_out;
  wire [0:19] sb_1__1__87_chany_bottom_out;
  wire [0:19] sb_1__1__87_chany_top_out;
  wire [0:0] sb_1__1__88_ccff_tail;
  wire [0:19] sb_1__1__88_chanx_left_out;
  wire [0:19] sb_1__1__88_chanx_right_out;
  wire [0:19] sb_1__1__88_chany_bottom_out;
  wire [0:19] sb_1__1__88_chany_top_out;
  wire [0:0] sb_1__1__89_ccff_tail;
  wire [0:19] sb_1__1__89_chanx_left_out;
  wire [0:19] sb_1__1__89_chanx_right_out;
  wire [0:19] sb_1__1__89_chany_bottom_out;
  wire [0:19] sb_1__1__89_chany_top_out;
  wire [0:0] sb_1__1__8_ccff_tail;
  wire [0:19] sb_1__1__8_chanx_left_out;
  wire [0:19] sb_1__1__8_chanx_right_out;
  wire [0:19] sb_1__1__8_chany_bottom_out;
  wire [0:19] sb_1__1__8_chany_top_out;
  wire [0:0] sb_1__1__90_ccff_tail;
  wire [0:19] sb_1__1__90_chanx_left_out;
  wire [0:19] sb_1__1__90_chanx_right_out;
  wire [0:19] sb_1__1__90_chany_bottom_out;
  wire [0:19] sb_1__1__90_chany_top_out;
  wire [0:0] sb_1__1__91_ccff_tail;
  wire [0:19] sb_1__1__91_chanx_left_out;
  wire [0:19] sb_1__1__91_chanx_right_out;
  wire [0:19] sb_1__1__91_chany_bottom_out;
  wire [0:19] sb_1__1__91_chany_top_out;
  wire [0:0] sb_1__1__92_ccff_tail;
  wire [0:19] sb_1__1__92_chanx_left_out;
  wire [0:19] sb_1__1__92_chanx_right_out;
  wire [0:19] sb_1__1__92_chany_bottom_out;
  wire [0:19] sb_1__1__92_chany_top_out;
  wire [0:0] sb_1__1__93_ccff_tail;
  wire [0:19] sb_1__1__93_chanx_left_out;
  wire [0:19] sb_1__1__93_chanx_right_out;
  wire [0:19] sb_1__1__93_chany_bottom_out;
  wire [0:19] sb_1__1__93_chany_top_out;
  wire [0:0] sb_1__1__94_ccff_tail;
  wire [0:19] sb_1__1__94_chanx_left_out;
  wire [0:19] sb_1__1__94_chanx_right_out;
  wire [0:19] sb_1__1__94_chany_bottom_out;
  wire [0:19] sb_1__1__94_chany_top_out;
  wire [0:0] sb_1__1__95_ccff_tail;
  wire [0:19] sb_1__1__95_chanx_left_out;
  wire [0:19] sb_1__1__95_chanx_right_out;
  wire [0:19] sb_1__1__95_chany_bottom_out;
  wire [0:19] sb_1__1__95_chany_top_out;
  wire [0:0] sb_1__1__96_ccff_tail;
  wire [0:19] sb_1__1__96_chanx_left_out;
  wire [0:19] sb_1__1__96_chanx_right_out;
  wire [0:19] sb_1__1__96_chany_bottom_out;
  wire [0:19] sb_1__1__96_chany_top_out;
  wire [0:0] sb_1__1__97_ccff_tail;
  wire [0:19] sb_1__1__97_chanx_left_out;
  wire [0:19] sb_1__1__97_chanx_right_out;
  wire [0:19] sb_1__1__97_chany_bottom_out;
  wire [0:19] sb_1__1__97_chany_top_out;
  wire [0:0] sb_1__1__98_ccff_tail;
  wire [0:19] sb_1__1__98_chanx_left_out;
  wire [0:19] sb_1__1__98_chanx_right_out;
  wire [0:19] sb_1__1__98_chany_bottom_out;
  wire [0:19] sb_1__1__98_chany_top_out;
  wire [0:0] sb_1__1__99_ccff_tail;
  wire [0:19] sb_1__1__99_chanx_left_out;
  wire [0:19] sb_1__1__99_chanx_right_out;
  wire [0:19] sb_1__1__99_chany_bottom_out;
  wire [0:19] sb_1__1__99_chany_top_out;
  wire [0:0] sb_1__1__9_ccff_tail;
  wire [0:19] sb_1__1__9_chanx_left_out;
  wire [0:19] sb_1__1__9_chanx_right_out;
  wire [0:19] sb_1__1__9_chany_bottom_out;
  wire [0:19] sb_1__1__9_chany_top_out;
  wire [1:0] UNCONN;
  wire [317:0] scff_Wires;
  wire [132:0] regin_feedthrough_wires;
  wire [132:0] regout_feedthrough_wires;
  wire [287:0] Test_enWires;
  wire [624:0] prog_clk_0_wires;
  wire [251:0] prog_clk_1_wires;
  wire [135:0] prog_clk_2_wires;
  wire [100:0] prog_clk_3_wires;
  wire [251:0] clk_1_wires;
  wire [135:0] clk_2_wires;
  wire [100:0] clk_3_wires;

  grid_clb
  grid_clb_1__1_
  (
    .clk_0_N_in(clk_1_wires[4]),
    .prog_clk_0_N_in(prog_clk_1_wires[4]),
    .prog_clk_0_W_out(prog_clk_0_wires[3]),
    .prog_clk_0_E_out(prog_clk_0_wires[1]),
    .prog_clk_0_S_out(prog_clk_0_wires[0]),
    .Test_en_E_in(Test_enWires[24]),
    .SC_OUT_BOT(scff_Wires[25]),
    .SC_IN_TOP(scff_Wires[23]),
    .top_width_0_height_0__pin_0_(cbx_1__1__0_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__0_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__0_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__0_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__0_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__0_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__0_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__0_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__0_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__0_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__0_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__0_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__0_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__0_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__0_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__0_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__0_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__0_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__0_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__0_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__0_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__0_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__0_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__0_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__0_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__0_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__0_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__0_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__0_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__0_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__0_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__0_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_0_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_0_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_0_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_0_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_0_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_0_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_0_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_0_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_0_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_0_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_0_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_0_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_0_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_0_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_0_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_0_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_0_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_0_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_0_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_0_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_0_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_0_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_0_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_0_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_0_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_0_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_0_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_0_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_0_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_0_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_0_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_0_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_0_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_1__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_0_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__2_
  (
    .clk_0_S_in(clk_1_wires[3]),
    .prog_clk_0_S_in(prog_clk_1_wires[3]),
    .prog_clk_0_W_out(prog_clk_0_wires[9]),
    .prog_clk_0_E_out(prog_clk_0_wires[7]),
    .prog_clk_0_S_out(prog_clk_0_wires[6]),
    .Test_en_E_in(Test_enWires[46]),
    .SC_OUT_BOT(scff_Wires[22]),
    .SC_IN_TOP(scff_Wires[21]),
    .top_width_0_height_0__pin_0_(cbx_1__1__1_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__1_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__1_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__1_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__1_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__1_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__1_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__1_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__1_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__1_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__1_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__1_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__1_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__1_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__1_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__1_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[1]),
    .right_width_0_height_0__pin_16_(cby_1__1__1_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__1_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__1_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__1_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__1_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__1_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__1_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__1_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__1_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__1_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__1_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__1_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__1_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__1_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__1_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__1_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_1_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_1_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_1_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_1_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_1_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_1_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_1_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_1_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_1_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_1_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_1_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_1_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_1_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_1_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_1_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_1_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_1_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_1_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_1_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_1_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_1_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_1_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_1_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_1_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_1_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_1_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_1_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_1_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_1_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_1_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_1_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_1_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_1_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[0]),
    .ccff_tail(grid_clb_1_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__3_
  (
    .clk_0_N_in(clk_1_wires[11]),
    .prog_clk_0_N_in(prog_clk_1_wires[11]),
    .prog_clk_0_W_out(prog_clk_0_wires[14]),
    .prog_clk_0_E_out(prog_clk_0_wires[12]),
    .prog_clk_0_S_out(prog_clk_0_wires[11]),
    .Test_en_E_in(Test_enWires[68]),
    .SC_OUT_BOT(scff_Wires[20]),
    .SC_IN_TOP(scff_Wires[19]),
    .top_width_0_height_0__pin_0_(cbx_1__1__2_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__2_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__2_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__2_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__2_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__2_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__2_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__2_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__2_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__2_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__2_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__2_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__2_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__2_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__2_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__2_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[2]),
    .right_width_0_height_0__pin_16_(cby_1__1__2_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__2_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__2_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__2_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__2_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__2_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__2_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__2_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__2_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__2_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__2_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__2_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__2_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__2_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__2_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__2_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_2_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_2_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_2_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_2_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_2_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_2_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_2_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_2_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_2_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_2_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_2_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_2_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_2_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_2_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_2_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_2_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_2_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_2_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_2_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_2_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_2_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_2_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_2_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_2_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_2_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_2_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_2_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_2_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_2_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_2_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_2_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_2_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_2_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[1]),
    .ccff_tail(grid_clb_2_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__4_
  (
    .clk_0_S_in(clk_1_wires[10]),
    .prog_clk_0_S_in(prog_clk_1_wires[10]),
    .prog_clk_0_W_out(prog_clk_0_wires[19]),
    .prog_clk_0_E_out(prog_clk_0_wires[17]),
    .prog_clk_0_S_out(prog_clk_0_wires[16]),
    .Test_en_E_in(Test_enWires[90]),
    .SC_OUT_BOT(scff_Wires[18]),
    .SC_IN_TOP(scff_Wires[17]),
    .top_width_0_height_0__pin_0_(cbx_1__1__3_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__3_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__3_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__3_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__3_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__3_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__3_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__3_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__3_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__3_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__3_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__3_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__3_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__3_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__3_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__3_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[3]),
    .right_width_0_height_0__pin_16_(cby_1__1__3_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__3_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__3_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__3_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__3_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__3_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__3_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__3_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__3_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__3_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__3_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__3_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__3_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__3_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__3_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__3_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_3_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_3_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_3_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_3_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_3_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_3_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_3_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_3_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_3_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_3_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_3_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_3_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_3_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_3_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_3_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_3_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_3_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_3_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_3_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_3_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_3_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_3_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_3_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_3_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_3_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_3_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_3_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_3_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_3_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_3_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_3_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_3_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_3_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[2]),
    .ccff_tail(grid_clb_3_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__5_
  (
    .clk_0_N_in(clk_1_wires[18]),
    .prog_clk_0_N_in(prog_clk_1_wires[18]),
    .prog_clk_0_W_out(prog_clk_0_wires[24]),
    .prog_clk_0_E_out(prog_clk_0_wires[22]),
    .prog_clk_0_S_out(prog_clk_0_wires[21]),
    .Test_en_E_in(Test_enWires[112]),
    .SC_OUT_BOT(scff_Wires[16]),
    .SC_IN_TOP(scff_Wires[15]),
    .top_width_0_height_0__pin_0_(cbx_1__1__4_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__4_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__4_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__4_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__4_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__4_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__4_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__4_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__4_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__4_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__4_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__4_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__4_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__4_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__4_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__4_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[4]),
    .right_width_0_height_0__pin_16_(cby_1__1__4_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__4_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__4_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__4_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__4_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__4_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__4_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__4_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__4_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__4_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__4_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__4_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__4_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__4_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__4_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__4_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_4_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_4_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_4_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_4_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_4_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_4_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_4_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_4_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_4_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_4_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_4_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_4_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_4_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_4_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_4_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_4_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_4_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_4_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_4_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_4_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_4_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_4_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_4_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_4_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_4_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_4_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_4_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_4_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_4_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_4_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_4_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_4_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_4_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[3]),
    .ccff_tail(grid_clb_4_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__6_
  (
    .clk_0_S_in(clk_1_wires[17]),
    .prog_clk_0_S_in(prog_clk_1_wires[17]),
    .prog_clk_0_W_out(prog_clk_0_wires[29]),
    .prog_clk_0_E_out(prog_clk_0_wires[27]),
    .prog_clk_0_S_out(prog_clk_0_wires[26]),
    .Test_en_E_in(Test_enWires[134]),
    .SC_OUT_BOT(scff_Wires[14]),
    .SC_IN_TOP(scff_Wires[13]),
    .top_width_0_height_0__pin_0_(cbx_1__1__5_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__5_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__5_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__5_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__5_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__5_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__5_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__5_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__5_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__5_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__5_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__5_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__5_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__5_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__5_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__5_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[5]),
    .right_width_0_height_0__pin_16_(cby_1__1__5_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__5_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__5_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__5_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__5_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__5_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__5_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__5_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__5_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__5_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__5_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__5_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__5_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__5_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__5_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__5_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_5_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_5_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_5_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_5_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_5_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_5_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_5_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_5_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_5_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_5_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_5_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_5_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_5_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_5_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_5_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_5_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_5_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_5_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_5_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_5_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_5_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_5_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_5_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_5_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_5_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_5_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_5_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_5_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_5_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_5_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_5_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_5_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_5_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[4]),
    .ccff_tail(grid_clb_5_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__7_
  (
    .clk_0_N_in(clk_1_wires[25]),
    .prog_clk_0_N_in(prog_clk_1_wires[25]),
    .prog_clk_0_W_out(prog_clk_0_wires[34]),
    .prog_clk_0_E_out(prog_clk_0_wires[32]),
    .prog_clk_0_S_out(prog_clk_0_wires[31]),
    .Test_en_E_in(Test_enWires[156]),
    .SC_OUT_BOT(scff_Wires[12]),
    .SC_IN_TOP(scff_Wires[11]),
    .top_width_0_height_0__pin_0_(cbx_1__1__6_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__6_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__6_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__6_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__6_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__6_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__6_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__6_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__6_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__6_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__6_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__6_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__6_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__6_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__6_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__6_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[6]),
    .right_width_0_height_0__pin_16_(cby_1__1__6_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__6_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__6_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__6_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__6_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__6_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__6_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__6_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__6_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__6_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__6_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__6_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__6_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__6_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__6_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__6_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_6_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_6_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_6_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_6_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_6_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_6_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_6_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_6_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_6_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_6_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_6_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_6_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_6_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_6_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_6_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_6_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_6_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_6_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_6_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_6_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_6_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_6_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_6_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_6_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_6_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_6_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_6_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_6_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_6_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_6_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_6_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_6_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_6_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[5]),
    .ccff_tail(grid_clb_6_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__8_
  (
    .clk_0_S_in(clk_1_wires[24]),
    .prog_clk_0_S_in(prog_clk_1_wires[24]),
    .prog_clk_0_W_out(prog_clk_0_wires[39]),
    .prog_clk_0_E_out(prog_clk_0_wires[37]),
    .prog_clk_0_S_out(prog_clk_0_wires[36]),
    .Test_en_E_in(Test_enWires[178]),
    .SC_OUT_BOT(scff_Wires[10]),
    .SC_IN_TOP(scff_Wires[9]),
    .top_width_0_height_0__pin_0_(cbx_1__1__7_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__7_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__7_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__7_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__7_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__7_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__7_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__7_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__7_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__7_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__7_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__7_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__7_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__7_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__7_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__7_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[7]),
    .right_width_0_height_0__pin_16_(cby_1__1__7_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__7_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__7_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__7_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__7_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__7_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__7_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__7_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__7_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__7_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__7_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__7_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__7_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__7_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__7_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__7_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_7_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_7_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_7_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_7_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_7_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_7_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_7_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_7_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_7_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_7_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_7_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_7_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_7_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_7_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_7_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_7_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_7_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_7_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_7_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_7_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_7_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_7_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_7_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_7_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_7_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_7_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_7_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_7_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_7_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_7_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_7_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_7_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_7_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[6]),
    .ccff_tail(grid_clb_7_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__9_
  (
    .clk_0_N_in(clk_1_wires[32]),
    .prog_clk_0_N_in(prog_clk_1_wires[32]),
    .prog_clk_0_W_out(prog_clk_0_wires[44]),
    .prog_clk_0_E_out(prog_clk_0_wires[42]),
    .prog_clk_0_S_out(prog_clk_0_wires[41]),
    .Test_en_E_in(Test_enWires[200]),
    .SC_OUT_BOT(scff_Wires[8]),
    .SC_IN_TOP(scff_Wires[7]),
    .top_width_0_height_0__pin_0_(cbx_1__1__8_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__8_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__8_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__8_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__8_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__8_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__8_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__8_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__8_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__8_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__8_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__8_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__8_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__8_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__8_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__8_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[8]),
    .right_width_0_height_0__pin_16_(cby_1__1__8_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__8_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__8_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__8_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__8_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__8_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__8_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__8_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__8_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__8_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__8_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__8_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__8_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__8_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__8_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__8_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_8_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_8_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_8_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_8_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_8_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_8_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_8_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_8_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_8_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_8_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_8_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_8_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_8_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_8_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_8_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_8_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_8_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_8_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_8_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_8_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_8_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_8_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_8_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_8_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_8_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_8_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_8_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_8_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_8_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_8_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_8_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_8_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_8_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[7]),
    .ccff_tail(grid_clb_8_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__10_
  (
    .clk_0_S_in(clk_1_wires[31]),
    .prog_clk_0_S_in(prog_clk_1_wires[31]),
    .prog_clk_0_W_out(prog_clk_0_wires[49]),
    .prog_clk_0_E_out(prog_clk_0_wires[47]),
    .prog_clk_0_S_out(prog_clk_0_wires[46]),
    .Test_en_E_in(Test_enWires[222]),
    .SC_OUT_BOT(scff_Wires[6]),
    .SC_IN_TOP(scff_Wires[5]),
    .top_width_0_height_0__pin_0_(cbx_1__1__9_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__9_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__9_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__9_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__9_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__9_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__9_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__9_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__9_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__9_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__9_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__9_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__9_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__9_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__9_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__9_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[9]),
    .right_width_0_height_0__pin_16_(cby_1__1__9_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__9_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__9_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__9_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__9_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__9_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__9_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__9_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__9_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__9_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__9_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__9_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__9_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__9_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__9_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__9_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_9_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_9_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_9_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_9_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_9_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_9_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_9_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_9_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_9_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_9_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_9_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_9_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_9_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_9_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_9_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_9_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_9_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_9_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_9_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_9_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_9_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_9_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_9_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_9_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_9_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_9_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_9_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_9_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_9_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_9_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_9_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_9_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_9_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[8]),
    .ccff_tail(grid_clb_9_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__11_
  (
    .clk_0_N_in(clk_1_wires[39]),
    .prog_clk_0_N_in(prog_clk_1_wires[39]),
    .prog_clk_0_W_out(prog_clk_0_wires[54]),
    .prog_clk_0_E_out(prog_clk_0_wires[52]),
    .prog_clk_0_S_out(prog_clk_0_wires[51]),
    .Test_en_E_in(Test_enWires[244]),
    .SC_OUT_BOT(scff_Wires[4]),
    .SC_IN_TOP(scff_Wires[3]),
    .top_width_0_height_0__pin_0_(cbx_1__1__10_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__10_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__10_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__10_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__10_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__10_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__10_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__10_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__10_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__10_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__10_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__10_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__10_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__10_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__10_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__10_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[10]),
    .right_width_0_height_0__pin_16_(cby_1__1__10_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__10_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__10_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__10_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__10_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__10_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__10_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__10_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__10_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__10_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__10_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__10_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__10_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__10_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__10_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__10_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_10_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_10_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_10_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_10_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_10_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_10_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_10_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_10_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_10_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_10_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_10_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_10_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_10_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_10_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_10_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_10_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_10_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_10_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_10_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_10_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_10_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_10_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_10_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_10_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_10_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_10_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_10_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_10_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_10_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_10_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_10_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_10_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_10_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[9]),
    .ccff_tail(grid_clb_10_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__12_
  (
    .clk_0_S_in(clk_1_wires[38]),
    .prog_clk_0_S_in(prog_clk_1_wires[38]),
    .prog_clk_0_W_out(prog_clk_0_wires[61]),
    .prog_clk_0_N_out(prog_clk_0_wires[59]),
    .prog_clk_0_E_out(prog_clk_0_wires[57]),
    .prog_clk_0_S_out(prog_clk_0_wires[56]),
    .Test_en_E_in(Test_enWires[266]),
    .SC_OUT_BOT(scff_Wires[2]),
    .SC_IN_TOP(scff_Wires[1]),
    .top_width_0_height_0__pin_0_(cbx_1__12__0_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__0_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__0_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__0_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__0_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__0_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__0_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__0_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__0_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__0_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__0_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__0_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__0_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__0_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__0_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__0_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_1__12__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__11_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__11_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__11_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__11_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__11_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__11_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__11_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__11_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__11_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__11_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__11_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__11_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__11_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__11_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__11_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__11_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_11_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_11_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_11_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_11_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_11_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_11_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_11_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_11_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_11_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_11_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_11_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_11_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_11_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_11_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_11_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_11_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_11_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_11_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_11_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_11_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_11_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_11_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_11_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_11_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_11_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_11_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_11_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_11_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_11_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_11_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_11_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_11_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_11_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[10]),
    .ccff_tail(grid_clb_11_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__1_
  (
    .clk_0_N_in(clk_1_wires[6]),
    .prog_clk_0_N_in(prog_clk_1_wires[6]),
    .prog_clk_0_E_out(prog_clk_0_wires[64]),
    .prog_clk_0_S_out(prog_clk_0_wires[63]),
    .Test_en_W_out(Test_enWires[26]),
    .Test_en_E_in(Test_enWires[25]),
    .SC_OUT_TOP(scff_Wires[29]),
    .SC_IN_BOT(scff_Wires[28]),
    .top_width_0_height_0__pin_0_(cbx_1__1__11_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__11_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__11_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__11_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__11_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__11_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__11_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__11_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__11_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__11_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__11_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__11_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__11_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__11_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__11_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__11_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[11]),
    .right_width_0_height_0__pin_16_(cby_1__1__12_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__12_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__12_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__12_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__12_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__12_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__12_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__12_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__12_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__12_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__12_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__12_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__12_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__12_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__12_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__12_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__0_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_12_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_12_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_12_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_12_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_12_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_12_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_12_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_12_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_12_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_12_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_12_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_12_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_12_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_12_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_12_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_12_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_12_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_12_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_12_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_12_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_12_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_12_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_12_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_12_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_12_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_12_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_12_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_12_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_12_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_12_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_12_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_12_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_2__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_12_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__2_
  (
    .clk_0_S_in(clk_1_wires[5]),
    .prog_clk_0_S_in(prog_clk_1_wires[5]),
    .prog_clk_0_E_out(prog_clk_0_wires[67]),
    .prog_clk_0_S_out(prog_clk_0_wires[66]),
    .Test_en_W_out(Test_enWires[48]),
    .Test_en_E_in(Test_enWires[47]),
    .SC_OUT_TOP(scff_Wires[31]),
    .SC_IN_BOT(scff_Wires[30]),
    .top_width_0_height_0__pin_0_(cbx_1__1__12_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__12_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__12_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__12_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__12_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__12_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__12_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__12_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__12_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__12_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__12_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__12_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__12_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__12_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__12_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__12_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[12]),
    .right_width_0_height_0__pin_16_(cby_1__1__13_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__13_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__13_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__13_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__13_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__13_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__13_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__13_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__13_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__13_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__13_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__13_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__13_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__13_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__13_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__13_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__1_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_13_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_13_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_13_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_13_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_13_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_13_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_13_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_13_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_13_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_13_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_13_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_13_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_13_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_13_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_13_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_13_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_13_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_13_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_13_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_13_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_13_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_13_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_13_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_13_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_13_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_13_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_13_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_13_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_13_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_13_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_13_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_13_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[11]),
    .ccff_tail(grid_clb_13_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__3_
  (
    .clk_0_N_in(clk_1_wires[13]),
    .prog_clk_0_N_in(prog_clk_1_wires[13]),
    .prog_clk_0_E_out(prog_clk_0_wires[70]),
    .prog_clk_0_S_out(prog_clk_0_wires[69]),
    .Test_en_W_out(Test_enWires[70]),
    .Test_en_E_in(Test_enWires[69]),
    .SC_OUT_TOP(scff_Wires[33]),
    .SC_IN_BOT(scff_Wires[32]),
    .top_width_0_height_0__pin_0_(cbx_1__1__13_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__13_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__13_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__13_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__13_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__13_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__13_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__13_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__13_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__13_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__13_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__13_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__13_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__13_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__13_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__13_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[13]),
    .right_width_0_height_0__pin_16_(cby_1__1__14_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__14_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__14_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__14_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__14_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__14_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__14_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__14_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__14_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__14_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__14_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__14_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__14_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__14_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__14_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__14_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__2_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_14_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_14_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_14_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_14_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_14_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_14_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_14_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_14_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_14_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_14_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_14_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_14_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_14_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_14_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_14_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_14_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_14_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_14_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_14_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_14_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_14_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_14_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_14_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_14_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_14_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_14_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_14_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_14_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_14_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_14_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_14_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_14_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[12]),
    .ccff_tail(grid_clb_14_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__4_
  (
    .clk_0_S_in(clk_1_wires[12]),
    .prog_clk_0_S_in(prog_clk_1_wires[12]),
    .prog_clk_0_E_out(prog_clk_0_wires[73]),
    .prog_clk_0_S_out(prog_clk_0_wires[72]),
    .Test_en_W_out(Test_enWires[92]),
    .Test_en_E_in(Test_enWires[91]),
    .SC_OUT_TOP(scff_Wires[35]),
    .SC_IN_BOT(scff_Wires[34]),
    .top_width_0_height_0__pin_0_(cbx_1__1__14_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__14_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__14_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__14_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__14_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__14_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__14_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__14_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__14_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__14_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__14_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__14_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__14_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__14_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__14_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__14_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[14]),
    .right_width_0_height_0__pin_16_(cby_1__1__15_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__15_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__15_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__15_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__15_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__15_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__15_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__15_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__15_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__15_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__15_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__15_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__15_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__15_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__15_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__15_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__3_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_15_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_15_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_15_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_15_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_15_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_15_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_15_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_15_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_15_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_15_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_15_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_15_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_15_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_15_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_15_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_15_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_15_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_15_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_15_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_15_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_15_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_15_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_15_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_15_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_15_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_15_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_15_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_15_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_15_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_15_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_15_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_15_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[13]),
    .ccff_tail(grid_clb_15_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__5_
  (
    .clk_0_N_in(clk_1_wires[20]),
    .prog_clk_0_N_in(prog_clk_1_wires[20]),
    .prog_clk_0_E_out(prog_clk_0_wires[76]),
    .prog_clk_0_S_out(prog_clk_0_wires[75]),
    .Test_en_W_out(Test_enWires[114]),
    .Test_en_E_in(Test_enWires[113]),
    .SC_OUT_TOP(scff_Wires[37]),
    .SC_IN_BOT(scff_Wires[36]),
    .top_width_0_height_0__pin_0_(cbx_1__1__15_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__15_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__15_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__15_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__15_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__15_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__15_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__15_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__15_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__15_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__15_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__15_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__15_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__15_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__15_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__15_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[15]),
    .right_width_0_height_0__pin_16_(cby_1__1__16_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__16_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__16_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__16_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__16_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__16_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__16_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__16_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__16_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__16_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__16_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__16_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__16_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__16_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__16_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__16_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__4_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_16_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_16_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_16_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_16_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_16_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_16_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_16_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_16_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_16_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_16_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_16_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_16_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_16_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_16_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_16_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_16_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_16_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_16_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_16_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_16_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_16_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_16_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_16_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_16_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_16_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_16_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_16_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_16_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_16_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_16_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_16_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_16_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[14]),
    .ccff_tail(grid_clb_16_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__6_
  (
    .clk_0_S_in(clk_1_wires[19]),
    .prog_clk_0_S_in(prog_clk_1_wires[19]),
    .prog_clk_0_E_out(prog_clk_0_wires[79]),
    .prog_clk_0_S_out(prog_clk_0_wires[78]),
    .Test_en_W_out(Test_enWires[136]),
    .Test_en_E_in(Test_enWires[135]),
    .SC_OUT_TOP(scff_Wires[39]),
    .SC_IN_BOT(scff_Wires[38]),
    .top_width_0_height_0__pin_0_(cbx_1__1__16_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__16_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__16_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__16_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__16_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__16_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__16_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__16_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__16_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__16_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__16_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__16_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__16_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__16_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__16_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__16_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[16]),
    .right_width_0_height_0__pin_16_(cby_1__1__17_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__17_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__17_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__17_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__17_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__17_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__17_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__17_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__17_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__17_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__17_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__17_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__17_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__17_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__17_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__17_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__5_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_17_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_17_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_17_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_17_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_17_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_17_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_17_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_17_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_17_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_17_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_17_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_17_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_17_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_17_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_17_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_17_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_17_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_17_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_17_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_17_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_17_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_17_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_17_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_17_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_17_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_17_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_17_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_17_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_17_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_17_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_17_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_17_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[15]),
    .ccff_tail(grid_clb_17_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__7_
  (
    .clk_0_N_in(clk_1_wires[27]),
    .prog_clk_0_N_in(prog_clk_1_wires[27]),
    .prog_clk_0_E_out(prog_clk_0_wires[82]),
    .prog_clk_0_S_out(prog_clk_0_wires[81]),
    .Test_en_W_out(Test_enWires[158]),
    .Test_en_E_in(Test_enWires[157]),
    .SC_OUT_TOP(scff_Wires[41]),
    .SC_IN_BOT(scff_Wires[40]),
    .top_width_0_height_0__pin_0_(cbx_1__1__17_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__17_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__17_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__17_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__17_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__17_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__17_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__17_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__17_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__17_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__17_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__17_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__17_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__17_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__17_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__17_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[17]),
    .right_width_0_height_0__pin_16_(cby_1__1__18_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__18_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__18_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__18_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__18_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__18_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__18_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__18_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__18_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__18_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__18_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__18_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__18_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__18_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__18_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__18_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__6_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_18_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_18_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_18_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_18_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_18_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_18_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_18_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_18_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_18_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_18_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_18_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_18_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_18_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_18_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_18_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_18_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_18_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_18_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_18_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_18_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_18_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_18_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_18_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_18_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_18_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_18_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_18_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_18_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_18_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_18_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_18_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_18_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[16]),
    .ccff_tail(grid_clb_18_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__8_
  (
    .clk_0_S_in(clk_1_wires[26]),
    .prog_clk_0_S_in(prog_clk_1_wires[26]),
    .prog_clk_0_E_out(prog_clk_0_wires[85]),
    .prog_clk_0_S_out(prog_clk_0_wires[84]),
    .Test_en_W_out(Test_enWires[180]),
    .Test_en_E_in(Test_enWires[179]),
    .SC_OUT_TOP(scff_Wires[43]),
    .SC_IN_BOT(scff_Wires[42]),
    .top_width_0_height_0__pin_0_(cbx_1__1__18_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__18_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__18_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__18_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__18_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__18_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__18_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__18_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__18_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__18_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__18_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__18_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__18_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__18_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__18_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__18_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[18]),
    .right_width_0_height_0__pin_16_(cby_1__1__19_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__19_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__19_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__19_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__19_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__19_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__19_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__19_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__19_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__19_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__19_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__19_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__19_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__19_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__19_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__19_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__7_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_19_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_19_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_19_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_19_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_19_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_19_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_19_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_19_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_19_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_19_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_19_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_19_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_19_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_19_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_19_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_19_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_19_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_19_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_19_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_19_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_19_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_19_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_19_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_19_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_19_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_19_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_19_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_19_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_19_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_19_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_19_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_19_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[17]),
    .ccff_tail(grid_clb_19_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__9_
  (
    .clk_0_N_in(clk_1_wires[34]),
    .prog_clk_0_N_in(prog_clk_1_wires[34]),
    .prog_clk_0_E_out(prog_clk_0_wires[88]),
    .prog_clk_0_S_out(prog_clk_0_wires[87]),
    .Test_en_W_out(Test_enWires[202]),
    .Test_en_E_in(Test_enWires[201]),
    .SC_OUT_TOP(scff_Wires[45]),
    .SC_IN_BOT(scff_Wires[44]),
    .top_width_0_height_0__pin_0_(cbx_1__1__19_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__19_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__19_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__19_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__19_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__19_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__19_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__19_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__19_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__19_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__19_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__19_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__19_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__19_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__19_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__19_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[19]),
    .right_width_0_height_0__pin_16_(cby_1__1__20_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__20_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__20_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__20_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__20_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__20_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__20_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__20_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__20_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__20_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__20_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__20_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__20_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__20_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__20_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__20_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__8_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_20_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_20_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_20_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_20_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_20_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_20_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_20_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_20_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_20_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_20_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_20_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_20_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_20_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_20_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_20_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_20_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_20_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_20_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_20_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_20_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_20_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_20_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_20_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_20_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_20_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_20_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_20_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_20_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_20_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_20_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_20_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_20_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[18]),
    .ccff_tail(grid_clb_20_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__10_
  (
    .clk_0_S_in(clk_1_wires[33]),
    .prog_clk_0_S_in(prog_clk_1_wires[33]),
    .prog_clk_0_E_out(prog_clk_0_wires[91]),
    .prog_clk_0_S_out(prog_clk_0_wires[90]),
    .Test_en_W_out(Test_enWires[224]),
    .Test_en_E_in(Test_enWires[223]),
    .SC_OUT_TOP(scff_Wires[47]),
    .SC_IN_BOT(scff_Wires[46]),
    .top_width_0_height_0__pin_0_(cbx_1__1__20_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__20_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__20_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__20_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__20_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__20_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__20_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__20_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__20_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__20_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__20_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__20_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__20_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__20_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__20_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__20_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[20]),
    .right_width_0_height_0__pin_16_(cby_1__1__21_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__21_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__21_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__21_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__21_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__21_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__21_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__21_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__21_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__21_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__21_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__21_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__21_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__21_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__21_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__21_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__9_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_21_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_21_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_21_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_21_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_21_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_21_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_21_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_21_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_21_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_21_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_21_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_21_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_21_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_21_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_21_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_21_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_21_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_21_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_21_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_21_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_21_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_21_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_21_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_21_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_21_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_21_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_21_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_21_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_21_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_21_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_21_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_21_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[19]),
    .ccff_tail(grid_clb_21_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__11_
  (
    .clk_0_N_in(clk_1_wires[41]),
    .prog_clk_0_N_in(prog_clk_1_wires[41]),
    .prog_clk_0_E_out(prog_clk_0_wires[94]),
    .prog_clk_0_S_out(prog_clk_0_wires[93]),
    .Test_en_W_out(Test_enWires[246]),
    .Test_en_E_in(Test_enWires[245]),
    .SC_OUT_TOP(scff_Wires[49]),
    .SC_IN_BOT(scff_Wires[48]),
    .top_width_0_height_0__pin_0_(cbx_1__1__21_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__21_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__21_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__21_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__21_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__21_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__21_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__21_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__21_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__21_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__21_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__21_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__21_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__21_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__21_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__21_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[21]),
    .right_width_0_height_0__pin_16_(cby_1__1__22_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__22_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__22_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__22_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__22_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__22_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__22_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__22_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__22_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__22_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__22_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__22_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__22_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__22_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__22_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__22_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__10_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_22_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_22_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_22_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_22_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_22_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_22_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_22_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_22_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_22_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_22_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_22_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_22_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_22_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_22_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_22_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_22_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_22_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_22_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_22_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_22_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_22_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_22_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_22_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_22_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_22_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_22_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_22_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_22_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_22_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_22_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_22_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_22_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[20]),
    .ccff_tail(grid_clb_22_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__12_
  (
    .clk_0_S_in(clk_1_wires[40]),
    .prog_clk_0_S_in(prog_clk_1_wires[40]),
    .prog_clk_0_N_out(prog_clk_0_wires[99]),
    .prog_clk_0_E_out(prog_clk_0_wires[97]),
    .prog_clk_0_S_out(prog_clk_0_wires[96]),
    .Test_en_W_out(Test_enWires[268]),
    .Test_en_E_in(Test_enWires[267]),
    .SC_OUT_TOP(scff_Wires[51]),
    .SC_IN_BOT(scff_Wires[50]),
    .top_width_0_height_0__pin_0_(cbx_1__12__1_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__1_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__1_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__1_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__1_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__1_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__1_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__1_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__1_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__1_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__1_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__1_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__1_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__1_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__1_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__1_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_2__12__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__23_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__23_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__23_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__23_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__23_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__23_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__23_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__23_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__23_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__23_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__23_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__23_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__23_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__23_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__23_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__23_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__11_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_23_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_23_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_23_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_23_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_23_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_23_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_23_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_23_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_23_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_23_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_23_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_23_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_23_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_23_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_23_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_23_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_23_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_23_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_23_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_23_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_23_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_23_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_23_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_23_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_23_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_23_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_23_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_23_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_23_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_23_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_23_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_23_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[21]),
    .ccff_tail(grid_clb_23_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__1_
  (
    .clk_0_N_in(clk_1_wires[46]),
    .prog_clk_0_N_in(prog_clk_1_wires[46]),
    .prog_clk_0_E_out(prog_clk_0_wires[102]),
    .prog_clk_0_S_out(prog_clk_0_wires[101]),
    .Test_en_W_out(Test_enWires[28]),
    .Test_en_E_in(Test_enWires[27]),
    .SC_OUT_BOT(scff_Wires[78]),
    .SC_IN_TOP(scff_Wires[76]),
    .top_width_0_height_0__pin_0_(cbx_1__1__22_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__22_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__22_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__22_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__22_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__22_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__22_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__22_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__22_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__22_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__22_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__22_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__22_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__22_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__22_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__22_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[22]),
    .right_width_0_height_0__pin_16_(cby_1__1__24_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__24_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__24_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__24_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__24_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__24_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__24_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__24_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__24_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__24_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__24_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__24_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__24_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__24_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__24_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__24_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__12_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_24_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_24_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_24_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_24_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_24_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_24_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_24_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_24_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_24_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_24_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_24_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_24_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_24_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_24_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_24_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_24_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_24_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_24_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_24_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_24_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_24_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_24_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_24_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_24_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_24_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_24_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_24_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_24_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_24_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_24_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_24_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_24_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_3__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_24_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__2_
  (
    .clk_0_S_in(clk_1_wires[45]),
    .prog_clk_0_S_in(prog_clk_1_wires[45]),
    .prog_clk_0_E_out(prog_clk_0_wires[105]),
    .prog_clk_0_S_out(prog_clk_0_wires[104]),
    .Test_en_W_out(Test_enWires[50]),
    .Test_en_E_in(Test_enWires[49]),
    .SC_OUT_BOT(scff_Wires[75]),
    .SC_IN_TOP(scff_Wires[74]),
    .top_width_0_height_0__pin_0_(cbx_1__1__23_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__23_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__23_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__23_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__23_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__23_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__23_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__23_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__23_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__23_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__23_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__23_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__23_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__23_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__23_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__23_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[23]),
    .right_width_0_height_0__pin_16_(cby_1__1__25_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__25_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__25_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__25_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__25_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__25_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__25_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__25_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__25_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__25_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__25_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__25_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__25_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__25_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__25_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__25_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__13_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_25_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_25_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_25_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_25_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_25_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_25_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_25_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_25_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_25_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_25_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_25_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_25_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_25_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_25_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_25_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_25_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_25_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_25_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_25_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_25_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_25_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_25_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_25_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_25_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_25_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_25_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_25_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_25_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_25_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_25_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_25_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_25_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[22]),
    .ccff_tail(grid_clb_25_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__3_
  (
    .clk_0_N_in(clk_1_wires[53]),
    .prog_clk_0_N_in(prog_clk_1_wires[53]),
    .prog_clk_0_E_out(prog_clk_0_wires[108]),
    .prog_clk_0_S_out(prog_clk_0_wires[107]),
    .Test_en_W_out(Test_enWires[72]),
    .Test_en_E_in(Test_enWires[71]),
    .SC_OUT_BOT(scff_Wires[73]),
    .SC_IN_TOP(scff_Wires[72]),
    .top_width_0_height_0__pin_0_(cbx_1__1__24_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__24_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__24_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__24_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__24_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__24_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__24_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__24_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__24_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__24_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__24_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__24_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__24_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__24_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__24_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__24_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[24]),
    .right_width_0_height_0__pin_16_(cby_1__1__26_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__26_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__26_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__26_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__26_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__26_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__26_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__26_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__26_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__26_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__26_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__26_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__26_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__26_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__26_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__26_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__14_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_26_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_26_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_26_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_26_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_26_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_26_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_26_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_26_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_26_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_26_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_26_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_26_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_26_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_26_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_26_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_26_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_26_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_26_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_26_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_26_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_26_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_26_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_26_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_26_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_26_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_26_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_26_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_26_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_26_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_26_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_26_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_26_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[23]),
    .ccff_tail(grid_clb_26_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__4_
  (
    .clk_0_S_in(clk_1_wires[52]),
    .prog_clk_0_S_in(prog_clk_1_wires[52]),
    .prog_clk_0_E_out(prog_clk_0_wires[111]),
    .prog_clk_0_S_out(prog_clk_0_wires[110]),
    .Test_en_W_out(Test_enWires[94]),
    .Test_en_E_in(Test_enWires[93]),
    .SC_OUT_BOT(scff_Wires[71]),
    .SC_IN_TOP(scff_Wires[70]),
    .top_width_0_height_0__pin_0_(cbx_1__1__25_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__25_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__25_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__25_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__25_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__25_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__25_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__25_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__25_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__25_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__25_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__25_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__25_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__25_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__25_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__25_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[25]),
    .right_width_0_height_0__pin_16_(cby_1__1__27_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__27_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__27_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__27_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__27_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__27_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__27_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__27_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__27_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__27_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__27_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__27_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__27_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__27_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__27_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__27_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__15_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_27_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_27_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_27_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_27_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_27_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_27_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_27_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_27_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_27_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_27_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_27_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_27_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_27_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_27_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_27_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_27_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_27_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_27_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_27_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_27_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_27_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_27_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_27_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_27_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_27_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_27_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_27_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_27_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_27_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_27_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_27_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_27_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[24]),
    .ccff_tail(grid_clb_27_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__5_
  (
    .clk_0_N_in(clk_1_wires[60]),
    .prog_clk_0_N_in(prog_clk_1_wires[60]),
    .prog_clk_0_E_out(prog_clk_0_wires[114]),
    .prog_clk_0_S_out(prog_clk_0_wires[113]),
    .Test_en_W_out(Test_enWires[116]),
    .Test_en_E_in(Test_enWires[115]),
    .SC_OUT_BOT(scff_Wires[69]),
    .SC_IN_TOP(scff_Wires[68]),
    .top_width_0_height_0__pin_0_(cbx_1__1__26_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__26_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__26_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__26_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__26_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__26_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__26_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__26_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__26_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__26_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__26_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__26_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__26_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__26_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__26_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__26_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[26]),
    .right_width_0_height_0__pin_16_(cby_1__1__28_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__28_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__28_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__28_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__28_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__28_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__28_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__28_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__28_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__28_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__28_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__28_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__28_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__28_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__28_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__28_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__16_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_28_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_28_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_28_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_28_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_28_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_28_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_28_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_28_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_28_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_28_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_28_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_28_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_28_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_28_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_28_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_28_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_28_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_28_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_28_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_28_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_28_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_28_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_28_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_28_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_28_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_28_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_28_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_28_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_28_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_28_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_28_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_28_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[25]),
    .ccff_tail(grid_clb_28_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__6_
  (
    .clk_0_S_in(clk_1_wires[59]),
    .prog_clk_0_S_in(prog_clk_1_wires[59]),
    .prog_clk_0_E_out(prog_clk_0_wires[117]),
    .prog_clk_0_S_out(prog_clk_0_wires[116]),
    .Test_en_W_out(Test_enWires[138]),
    .Test_en_E_in(Test_enWires[137]),
    .SC_OUT_BOT(scff_Wires[67]),
    .SC_IN_TOP(scff_Wires[66]),
    .top_width_0_height_0__pin_0_(cbx_1__1__27_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__27_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__27_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__27_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__27_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__27_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__27_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__27_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__27_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__27_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__27_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__27_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__27_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__27_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__27_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__27_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[27]),
    .right_width_0_height_0__pin_16_(cby_1__1__29_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__29_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__29_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__29_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__29_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__29_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__29_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__29_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__29_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__29_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__29_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__29_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__29_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__29_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__29_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__29_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__17_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_29_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_29_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_29_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_29_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_29_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_29_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_29_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_29_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_29_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_29_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_29_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_29_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_29_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_29_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_29_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_29_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_29_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_29_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_29_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_29_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_29_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_29_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_29_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_29_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_29_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_29_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_29_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_29_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_29_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_29_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_29_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_29_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[26]),
    .ccff_tail(grid_clb_29_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__7_
  (
    .clk_0_N_in(clk_1_wires[67]),
    .prog_clk_0_N_in(prog_clk_1_wires[67]),
    .prog_clk_0_E_out(prog_clk_0_wires[120]),
    .prog_clk_0_S_out(prog_clk_0_wires[119]),
    .Test_en_W_out(Test_enWires[160]),
    .Test_en_E_in(Test_enWires[159]),
    .SC_OUT_BOT(scff_Wires[65]),
    .SC_IN_TOP(scff_Wires[64]),
    .top_width_0_height_0__pin_0_(cbx_1__1__28_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__28_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__28_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__28_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__28_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__28_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__28_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__28_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__28_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__28_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__28_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__28_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__28_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__28_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__28_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__28_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[28]),
    .right_width_0_height_0__pin_16_(cby_1__1__30_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__30_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__30_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__30_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__30_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__30_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__30_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__30_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__30_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__30_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__30_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__30_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__30_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__30_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__30_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__30_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__18_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_30_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_30_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_30_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_30_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_30_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_30_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_30_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_30_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_30_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_30_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_30_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_30_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_30_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_30_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_30_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_30_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_30_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_30_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_30_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_30_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_30_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_30_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_30_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_30_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_30_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_30_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_30_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_30_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_30_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_30_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_30_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_30_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[27]),
    .ccff_tail(grid_clb_30_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__8_
  (
    .clk_0_S_in(clk_1_wires[66]),
    .prog_clk_0_S_in(prog_clk_1_wires[66]),
    .prog_clk_0_E_out(prog_clk_0_wires[123]),
    .prog_clk_0_S_out(prog_clk_0_wires[122]),
    .Test_en_W_out(Test_enWires[182]),
    .Test_en_E_in(Test_enWires[181]),
    .SC_OUT_BOT(scff_Wires[63]),
    .SC_IN_TOP(scff_Wires[62]),
    .top_width_0_height_0__pin_0_(cbx_1__1__29_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__29_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__29_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__29_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__29_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__29_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__29_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__29_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__29_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__29_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__29_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__29_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__29_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__29_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__29_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__29_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[29]),
    .right_width_0_height_0__pin_16_(cby_1__1__31_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__31_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__31_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__31_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__31_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__31_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__31_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__31_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__31_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__31_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__31_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__31_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__31_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__31_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__31_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__31_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__19_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_31_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_31_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_31_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_31_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_31_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_31_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_31_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_31_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_31_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_31_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_31_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_31_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_31_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_31_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_31_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_31_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_31_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_31_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_31_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_31_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_31_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_31_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_31_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_31_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_31_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_31_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_31_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_31_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_31_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_31_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_31_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_31_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[28]),
    .ccff_tail(grid_clb_31_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__9_
  (
    .clk_0_N_in(clk_1_wires[74]),
    .prog_clk_0_N_in(prog_clk_1_wires[74]),
    .prog_clk_0_E_out(prog_clk_0_wires[126]),
    .prog_clk_0_S_out(prog_clk_0_wires[125]),
    .Test_en_W_out(Test_enWires[204]),
    .Test_en_E_in(Test_enWires[203]),
    .SC_OUT_BOT(scff_Wires[61]),
    .SC_IN_TOP(scff_Wires[60]),
    .top_width_0_height_0__pin_0_(cbx_1__1__30_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__30_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__30_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__30_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__30_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__30_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__30_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__30_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__30_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__30_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__30_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__30_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__30_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__30_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__30_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__30_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[30]),
    .right_width_0_height_0__pin_16_(cby_1__1__32_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__32_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__32_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__32_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__32_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__32_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__32_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__32_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__32_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__32_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__32_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__32_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__32_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__32_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__32_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__32_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__20_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_32_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_32_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_32_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_32_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_32_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_32_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_32_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_32_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_32_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_32_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_32_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_32_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_32_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_32_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_32_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_32_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_32_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_32_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_32_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_32_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_32_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_32_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_32_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_32_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_32_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_32_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_32_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_32_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_32_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_32_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_32_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_32_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[29]),
    .ccff_tail(grid_clb_32_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__10_
  (
    .clk_0_S_in(clk_1_wires[73]),
    .prog_clk_0_S_in(prog_clk_1_wires[73]),
    .prog_clk_0_E_out(prog_clk_0_wires[129]),
    .prog_clk_0_S_out(prog_clk_0_wires[128]),
    .Test_en_W_out(Test_enWires[226]),
    .Test_en_E_in(Test_enWires[225]),
    .SC_OUT_BOT(scff_Wires[59]),
    .SC_IN_TOP(scff_Wires[58]),
    .top_width_0_height_0__pin_0_(cbx_1__1__31_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__31_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__31_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__31_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__31_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__31_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__31_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__31_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__31_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__31_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__31_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__31_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__31_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__31_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__31_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__31_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[31]),
    .right_width_0_height_0__pin_16_(cby_1__1__33_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__33_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__33_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__33_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__33_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__33_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__33_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__33_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__33_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__33_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__33_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__33_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__33_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__33_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__33_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__33_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__21_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_33_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_33_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_33_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_33_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_33_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_33_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_33_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_33_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_33_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_33_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_33_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_33_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_33_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_33_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_33_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_33_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_33_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_33_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_33_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_33_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_33_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_33_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_33_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_33_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_33_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_33_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_33_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_33_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_33_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_33_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_33_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_33_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[30]),
    .ccff_tail(grid_clb_33_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__11_
  (
    .clk_0_N_in(clk_1_wires[81]),
    .prog_clk_0_N_in(prog_clk_1_wires[81]),
    .prog_clk_0_E_out(prog_clk_0_wires[132]),
    .prog_clk_0_S_out(prog_clk_0_wires[131]),
    .Test_en_W_out(Test_enWires[248]),
    .Test_en_E_in(Test_enWires[247]),
    .SC_OUT_BOT(scff_Wires[57]),
    .SC_IN_TOP(scff_Wires[56]),
    .top_width_0_height_0__pin_0_(cbx_1__1__32_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__32_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__32_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__32_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__32_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__32_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__32_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__32_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__32_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__32_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__32_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__32_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__32_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__32_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__32_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__32_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[32]),
    .right_width_0_height_0__pin_16_(cby_1__1__34_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__34_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__34_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__34_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__34_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__34_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__34_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__34_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__34_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__34_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__34_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__34_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__34_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__34_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__34_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__34_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__22_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_34_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_34_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_34_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_34_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_34_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_34_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_34_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_34_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_34_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_34_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_34_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_34_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_34_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_34_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_34_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_34_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_34_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_34_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_34_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_34_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_34_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_34_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_34_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_34_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_34_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_34_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_34_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_34_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_34_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_34_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_34_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_34_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[31]),
    .ccff_tail(grid_clb_34_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__12_
  (
    .clk_0_S_in(clk_1_wires[80]),
    .prog_clk_0_S_in(prog_clk_1_wires[80]),
    .prog_clk_0_N_out(prog_clk_0_wires[137]),
    .prog_clk_0_E_out(prog_clk_0_wires[135]),
    .prog_clk_0_S_out(prog_clk_0_wires[134]),
    .Test_en_W_out(Test_enWires[270]),
    .Test_en_E_in(Test_enWires[269]),
    .SC_OUT_BOT(scff_Wires[55]),
    .SC_IN_TOP(scff_Wires[54]),
    .top_width_0_height_0__pin_0_(cbx_1__12__2_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__2_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__2_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__2_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__2_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__2_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__2_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__2_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__2_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__2_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__2_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__2_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__2_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__2_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__2_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__2_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_3__12__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__35_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__35_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__35_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__35_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__35_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__35_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__35_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__35_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__35_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__35_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__35_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__35_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__35_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__35_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__35_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__35_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__23_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_35_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_35_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_35_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_35_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_35_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_35_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_35_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_35_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_35_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_35_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_35_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_35_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_35_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_35_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_35_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_35_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_35_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_35_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_35_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_35_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_35_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_35_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_35_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_35_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_35_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_35_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_35_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_35_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_35_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_35_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_35_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_35_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[32]),
    .ccff_tail(grid_clb_35_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__1_
  (
    .clk_0_N_in(clk_1_wires[48]),
    .prog_clk_0_N_in(prog_clk_1_wires[48]),
    .prog_clk_0_E_out(prog_clk_0_wires[140]),
    .prog_clk_0_S_out(prog_clk_0_wires[139]),
    .Test_en_W_out(Test_enWires[30]),
    .Test_en_E_in(Test_enWires[29]),
    .SC_OUT_TOP(scff_Wires[82]),
    .SC_IN_BOT(scff_Wires[81]),
    .top_width_0_height_0__pin_0_(cbx_1__1__33_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__33_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__33_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__33_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__33_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__33_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__33_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__33_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__33_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__33_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__33_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__33_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__33_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__33_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__33_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__33_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[33]),
    .right_width_0_height_0__pin_16_(cby_1__1__36_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__36_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__36_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__36_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__36_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__36_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__36_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__36_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__36_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__36_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__36_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__36_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__36_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__36_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__36_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__36_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__24_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_36_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_36_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_36_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_36_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_36_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_36_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_36_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_36_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_36_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_36_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_36_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_36_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_36_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_36_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_36_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_36_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_36_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_36_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_36_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_36_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_36_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_36_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_36_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_36_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_36_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_36_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_36_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_36_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_36_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_36_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_36_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_36_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_4__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_36_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__2_
  (
    .clk_0_S_in(clk_1_wires[47]),
    .prog_clk_0_S_in(prog_clk_1_wires[47]),
    .prog_clk_0_E_out(prog_clk_0_wires[143]),
    .prog_clk_0_S_out(prog_clk_0_wires[142]),
    .Test_en_W_out(Test_enWires[52]),
    .Test_en_E_in(Test_enWires[51]),
    .SC_OUT_TOP(scff_Wires[84]),
    .SC_IN_BOT(scff_Wires[83]),
    .top_width_0_height_0__pin_0_(cbx_1__1__34_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__34_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__34_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__34_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__34_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__34_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__34_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__34_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__34_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__34_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__34_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__34_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__34_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__34_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__34_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__34_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[34]),
    .right_width_0_height_0__pin_16_(cby_1__1__37_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__37_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__37_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__37_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__37_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__37_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__37_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__37_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__37_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__37_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__37_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__37_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__37_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__37_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__37_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__37_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__25_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_37_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_37_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_37_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_37_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_37_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_37_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_37_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_37_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_37_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_37_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_37_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_37_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_37_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_37_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_37_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_37_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_37_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_37_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_37_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_37_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_37_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_37_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_37_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_37_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_37_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_37_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_37_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_37_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_37_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_37_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_37_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_37_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[33]),
    .ccff_tail(grid_clb_37_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__3_
  (
    .clk_0_N_in(clk_1_wires[55]),
    .prog_clk_0_N_in(prog_clk_1_wires[55]),
    .prog_clk_0_E_out(prog_clk_0_wires[146]),
    .prog_clk_0_S_out(prog_clk_0_wires[145]),
    .Test_en_W_out(Test_enWires[74]),
    .Test_en_E_in(Test_enWires[73]),
    .SC_OUT_TOP(scff_Wires[86]),
    .SC_IN_BOT(scff_Wires[85]),
    .top_width_0_height_0__pin_0_(cbx_1__1__35_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__35_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__35_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__35_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__35_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__35_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__35_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__35_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__35_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__35_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__35_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__35_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__35_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__35_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__35_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__35_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[35]),
    .right_width_0_height_0__pin_16_(cby_1__1__38_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__38_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__38_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__38_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__38_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__38_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__38_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__38_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__38_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__38_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__38_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__38_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__38_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__38_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__38_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__38_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__26_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_38_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_38_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_38_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_38_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_38_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_38_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_38_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_38_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_38_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_38_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_38_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_38_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_38_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_38_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_38_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_38_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_38_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_38_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_38_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_38_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_38_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_38_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_38_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_38_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_38_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_38_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_38_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_38_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_38_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_38_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_38_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_38_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[34]),
    .ccff_tail(grid_clb_38_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__4_
  (
    .clk_0_S_in(clk_1_wires[54]),
    .prog_clk_0_S_in(prog_clk_1_wires[54]),
    .prog_clk_0_E_out(prog_clk_0_wires[149]),
    .prog_clk_0_S_out(prog_clk_0_wires[148]),
    .Test_en_W_out(Test_enWires[96]),
    .Test_en_E_in(Test_enWires[95]),
    .SC_OUT_TOP(scff_Wires[88]),
    .SC_IN_BOT(scff_Wires[87]),
    .top_width_0_height_0__pin_0_(cbx_1__1__36_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__36_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__36_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__36_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__36_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__36_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__36_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__36_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__36_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__36_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__36_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__36_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__36_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__36_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__36_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__36_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[36]),
    .right_width_0_height_0__pin_16_(cby_1__1__39_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__39_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__39_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__39_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__39_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__39_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__39_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__39_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__39_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__39_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__39_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__39_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__39_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__39_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__39_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__39_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__27_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_39_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_39_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_39_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_39_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_39_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_39_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_39_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_39_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_39_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_39_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_39_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_39_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_39_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_39_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_39_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_39_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_39_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_39_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_39_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_39_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_39_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_39_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_39_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_39_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_39_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_39_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_39_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_39_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_39_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_39_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_39_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_39_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[35]),
    .ccff_tail(grid_clb_39_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__5_
  (
    .clk_0_N_in(clk_1_wires[62]),
    .prog_clk_0_N_in(prog_clk_1_wires[62]),
    .prog_clk_0_E_out(prog_clk_0_wires[152]),
    .prog_clk_0_S_out(prog_clk_0_wires[151]),
    .Test_en_W_out(Test_enWires[118]),
    .Test_en_E_in(Test_enWires[117]),
    .SC_OUT_TOP(scff_Wires[90]),
    .SC_IN_BOT(scff_Wires[89]),
    .top_width_0_height_0__pin_0_(cbx_1__1__37_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__37_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__37_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__37_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__37_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__37_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__37_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__37_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__37_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__37_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__37_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__37_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__37_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__37_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__37_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__37_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[37]),
    .right_width_0_height_0__pin_16_(cby_1__1__40_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__40_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__40_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__40_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__40_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__40_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__40_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__40_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__40_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__40_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__40_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__40_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__40_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__40_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__40_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__40_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__28_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_40_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_40_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_40_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_40_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_40_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_40_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_40_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_40_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_40_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_40_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_40_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_40_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_40_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_40_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_40_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_40_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_40_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_40_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_40_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_40_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_40_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_40_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_40_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_40_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_40_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_40_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_40_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_40_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_40_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_40_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_40_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_40_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[36]),
    .ccff_tail(grid_clb_40_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__6_
  (
    .clk_0_S_in(clk_1_wires[61]),
    .prog_clk_0_S_in(prog_clk_1_wires[61]),
    .prog_clk_0_E_out(prog_clk_0_wires[155]),
    .prog_clk_0_S_out(prog_clk_0_wires[154]),
    .Test_en_W_out(Test_enWires[140]),
    .Test_en_E_in(Test_enWires[139]),
    .SC_OUT_TOP(scff_Wires[92]),
    .SC_IN_BOT(scff_Wires[91]),
    .top_width_0_height_0__pin_0_(cbx_1__1__38_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__38_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__38_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__38_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__38_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__38_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__38_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__38_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__38_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__38_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__38_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__38_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__38_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__38_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__38_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__38_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[38]),
    .right_width_0_height_0__pin_16_(cby_1__1__41_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__41_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__41_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__41_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__41_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__41_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__41_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__41_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__41_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__41_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__41_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__41_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__41_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__41_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__41_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__41_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__29_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_41_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_41_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_41_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_41_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_41_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_41_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_41_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_41_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_41_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_41_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_41_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_41_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_41_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_41_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_41_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_41_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_41_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_41_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_41_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_41_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_41_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_41_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_41_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_41_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_41_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_41_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_41_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_41_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_41_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_41_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_41_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_41_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[37]),
    .ccff_tail(grid_clb_41_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__7_
  (
    .clk_0_N_in(clk_1_wires[69]),
    .prog_clk_0_N_in(prog_clk_1_wires[69]),
    .prog_clk_0_E_out(prog_clk_0_wires[158]),
    .prog_clk_0_S_out(prog_clk_0_wires[157]),
    .Test_en_W_out(Test_enWires[162]),
    .Test_en_E_in(Test_enWires[161]),
    .SC_OUT_TOP(scff_Wires[94]),
    .SC_IN_BOT(scff_Wires[93]),
    .top_width_0_height_0__pin_0_(cbx_1__1__39_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__39_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__39_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__39_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__39_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__39_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__39_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__39_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__39_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__39_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__39_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__39_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__39_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__39_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__39_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__39_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[39]),
    .right_width_0_height_0__pin_16_(cby_1__1__42_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__42_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__42_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__42_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__42_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__42_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__42_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__42_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__42_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__42_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__42_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__42_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__42_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__42_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__42_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__42_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__30_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_42_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_42_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_42_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_42_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_42_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_42_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_42_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_42_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_42_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_42_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_42_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_42_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_42_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_42_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_42_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_42_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_42_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_42_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_42_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_42_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_42_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_42_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_42_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_42_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_42_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_42_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_42_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_42_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_42_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_42_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_42_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_42_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[38]),
    .ccff_tail(grid_clb_42_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__8_
  (
    .clk_0_S_in(clk_1_wires[68]),
    .prog_clk_0_S_in(prog_clk_1_wires[68]),
    .prog_clk_0_E_out(prog_clk_0_wires[161]),
    .prog_clk_0_S_out(prog_clk_0_wires[160]),
    .Test_en_W_out(Test_enWires[184]),
    .Test_en_E_in(Test_enWires[183]),
    .SC_OUT_TOP(scff_Wires[96]),
    .SC_IN_BOT(scff_Wires[95]),
    .top_width_0_height_0__pin_0_(cbx_1__1__40_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__40_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__40_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__40_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__40_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__40_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__40_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__40_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__40_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__40_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__40_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__40_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__40_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__40_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__40_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__40_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[40]),
    .right_width_0_height_0__pin_16_(cby_1__1__43_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__43_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__43_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__43_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__43_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__43_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__43_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__43_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__43_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__43_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__43_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__43_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__43_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__43_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__43_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__43_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__31_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_43_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_43_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_43_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_43_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_43_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_43_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_43_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_43_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_43_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_43_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_43_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_43_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_43_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_43_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_43_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_43_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_43_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_43_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_43_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_43_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_43_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_43_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_43_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_43_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_43_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_43_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_43_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_43_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_43_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_43_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_43_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_43_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[39]),
    .ccff_tail(grid_clb_43_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__9_
  (
    .clk_0_N_in(clk_1_wires[76]),
    .prog_clk_0_N_in(prog_clk_1_wires[76]),
    .prog_clk_0_E_out(prog_clk_0_wires[164]),
    .prog_clk_0_S_out(prog_clk_0_wires[163]),
    .Test_en_W_out(Test_enWires[206]),
    .Test_en_E_in(Test_enWires[205]),
    .SC_OUT_TOP(scff_Wires[98]),
    .SC_IN_BOT(scff_Wires[97]),
    .top_width_0_height_0__pin_0_(cbx_1__1__41_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__41_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__41_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__41_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__41_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__41_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__41_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__41_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__41_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__41_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__41_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__41_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__41_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__41_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__41_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__41_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[41]),
    .right_width_0_height_0__pin_16_(cby_1__1__44_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__44_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__44_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__44_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__44_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__44_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__44_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__44_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__44_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__44_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__44_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__44_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__44_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__44_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__44_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__44_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__32_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_44_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_44_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_44_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_44_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_44_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_44_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_44_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_44_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_44_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_44_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_44_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_44_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_44_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_44_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_44_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_44_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_44_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_44_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_44_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_44_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_44_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_44_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_44_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_44_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_44_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_44_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_44_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_44_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_44_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_44_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_44_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_44_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[40]),
    .ccff_tail(grid_clb_44_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__10_
  (
    .clk_0_S_in(clk_1_wires[75]),
    .prog_clk_0_S_in(prog_clk_1_wires[75]),
    .prog_clk_0_E_out(prog_clk_0_wires[167]),
    .prog_clk_0_S_out(prog_clk_0_wires[166]),
    .Test_en_W_out(Test_enWires[228]),
    .Test_en_E_in(Test_enWires[227]),
    .SC_OUT_TOP(scff_Wires[100]),
    .SC_IN_BOT(scff_Wires[99]),
    .top_width_0_height_0__pin_0_(cbx_1__1__42_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__42_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__42_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__42_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__42_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__42_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__42_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__42_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__42_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__42_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__42_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__42_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__42_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__42_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__42_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__42_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[42]),
    .right_width_0_height_0__pin_16_(cby_1__1__45_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__45_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__45_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__45_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__45_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__45_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__45_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__45_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__45_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__45_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__45_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__45_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__45_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__45_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__45_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__45_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__33_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_45_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_45_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_45_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_45_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_45_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_45_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_45_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_45_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_45_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_45_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_45_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_45_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_45_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_45_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_45_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_45_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_45_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_45_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_45_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_45_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_45_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_45_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_45_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_45_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_45_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_45_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_45_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_45_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_45_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_45_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_45_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_45_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[41]),
    .ccff_tail(grid_clb_45_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__11_
  (
    .clk_0_N_in(clk_1_wires[83]),
    .prog_clk_0_N_in(prog_clk_1_wires[83]),
    .prog_clk_0_E_out(prog_clk_0_wires[170]),
    .prog_clk_0_S_out(prog_clk_0_wires[169]),
    .Test_en_W_out(Test_enWires[250]),
    .Test_en_E_in(Test_enWires[249]),
    .SC_OUT_TOP(scff_Wires[102]),
    .SC_IN_BOT(scff_Wires[101]),
    .top_width_0_height_0__pin_0_(cbx_1__1__43_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__43_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__43_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__43_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__43_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__43_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__43_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__43_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__43_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__43_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__43_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__43_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__43_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__43_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__43_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__43_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[43]),
    .right_width_0_height_0__pin_16_(cby_1__1__46_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__46_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__46_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__46_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__46_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__46_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__46_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__46_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__46_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__46_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__46_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__46_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__46_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__46_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__46_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__46_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__34_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_46_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_46_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_46_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_46_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_46_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_46_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_46_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_46_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_46_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_46_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_46_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_46_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_46_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_46_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_46_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_46_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_46_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_46_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_46_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_46_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_46_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_46_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_46_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_46_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_46_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_46_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_46_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_46_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_46_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_46_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_46_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_46_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[42]),
    .ccff_tail(grid_clb_46_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__12_
  (
    .clk_0_S_in(clk_1_wires[82]),
    .prog_clk_0_S_in(prog_clk_1_wires[82]),
    .prog_clk_0_N_out(prog_clk_0_wires[175]),
    .prog_clk_0_E_out(prog_clk_0_wires[173]),
    .prog_clk_0_S_out(prog_clk_0_wires[172]),
    .Test_en_W_out(Test_enWires[272]),
    .Test_en_E_in(Test_enWires[271]),
    .SC_OUT_TOP(scff_Wires[104]),
    .SC_IN_BOT(scff_Wires[103]),
    .top_width_0_height_0__pin_0_(cbx_1__12__3_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__3_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__3_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__3_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__3_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__3_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__3_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__3_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__3_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__3_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__3_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__3_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__3_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__3_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__3_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__3_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_4__12__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__47_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__47_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__47_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__47_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__47_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__47_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__47_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__47_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__47_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__47_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__47_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__47_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__47_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__47_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__47_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__47_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__35_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_47_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_47_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_47_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_47_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_47_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_47_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_47_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_47_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_47_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_47_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_47_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_47_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_47_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_47_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_47_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_47_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_47_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_47_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_47_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_47_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_47_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_47_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_47_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_47_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_47_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_47_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_47_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_47_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_47_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_47_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_47_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_47_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[43]),
    .ccff_tail(grid_clb_47_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__1_
  (
    .clk_0_N_in(clk_1_wires[88]),
    .prog_clk_0_N_in(prog_clk_1_wires[88]),
    .prog_clk_0_E_out(prog_clk_0_wires[178]),
    .prog_clk_0_S_out(prog_clk_0_wires[177]),
    .Test_en_W_out(Test_enWires[32]),
    .Test_en_E_in(Test_enWires[31]),
    .SC_OUT_BOT(scff_Wires[131]),
    .SC_IN_TOP(scff_Wires[129]),
    .top_width_0_height_0__pin_0_(cbx_1__1__44_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__44_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__44_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__44_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__44_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__44_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__44_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__44_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__44_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__44_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__44_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__44_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__44_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__44_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__44_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__44_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[44]),
    .right_width_0_height_0__pin_16_(cby_1__1__48_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__48_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__48_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__48_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__48_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__48_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__48_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__48_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__48_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__48_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__48_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__48_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__48_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__48_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__48_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__48_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__36_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_48_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_48_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_48_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_48_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_48_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_48_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_48_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_48_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_48_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_48_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_48_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_48_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_48_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_48_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_48_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_48_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_48_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_48_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_48_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_48_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_48_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_48_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_48_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_48_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_48_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_48_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_48_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_48_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_48_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_48_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_48_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_48_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_5__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_48_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__2_
  (
    .clk_0_S_in(clk_1_wires[87]),
    .prog_clk_0_S_in(prog_clk_1_wires[87]),
    .prog_clk_0_E_out(prog_clk_0_wires[181]),
    .prog_clk_0_S_out(prog_clk_0_wires[180]),
    .Test_en_W_out(Test_enWires[54]),
    .Test_en_E_in(Test_enWires[53]),
    .SC_OUT_BOT(scff_Wires[128]),
    .SC_IN_TOP(scff_Wires[127]),
    .top_width_0_height_0__pin_0_(cbx_1__1__45_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__45_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__45_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__45_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__45_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__45_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__45_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__45_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__45_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__45_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__45_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__45_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__45_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__45_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__45_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__45_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[45]),
    .right_width_0_height_0__pin_16_(cby_1__1__49_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__49_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__49_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__49_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__49_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__49_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__49_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__49_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__49_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__49_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__49_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__49_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__49_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__49_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__49_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__49_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__37_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_49_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_49_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_49_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_49_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_49_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_49_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_49_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_49_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_49_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_49_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_49_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_49_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_49_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_49_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_49_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_49_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_49_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_49_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_49_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_49_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_49_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_49_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_49_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_49_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_49_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_49_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_49_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_49_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_49_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_49_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_49_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_49_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[44]),
    .ccff_tail(grid_clb_49_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__3_
  (
    .clk_0_N_in(clk_1_wires[95]),
    .prog_clk_0_N_in(prog_clk_1_wires[95]),
    .prog_clk_0_E_out(prog_clk_0_wires[184]),
    .prog_clk_0_S_out(prog_clk_0_wires[183]),
    .Test_en_W_out(Test_enWires[76]),
    .Test_en_E_in(Test_enWires[75]),
    .SC_OUT_BOT(scff_Wires[126]),
    .SC_IN_TOP(scff_Wires[125]),
    .top_width_0_height_0__pin_0_(cbx_1__1__46_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__46_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__46_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__46_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__46_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__46_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__46_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__46_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__46_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__46_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__46_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__46_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__46_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__46_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__46_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__46_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[46]),
    .right_width_0_height_0__pin_16_(cby_1__1__50_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__50_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__50_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__50_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__50_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__50_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__50_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__50_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__50_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__50_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__50_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__50_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__50_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__50_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__50_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__50_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__38_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_50_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_50_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_50_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_50_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_50_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_50_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_50_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_50_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_50_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_50_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_50_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_50_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_50_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_50_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_50_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_50_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_50_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_50_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_50_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_50_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_50_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_50_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_50_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_50_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_50_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_50_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_50_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_50_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_50_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_50_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_50_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_50_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[45]),
    .ccff_tail(grid_clb_50_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__4_
  (
    .clk_0_S_in(clk_1_wires[94]),
    .prog_clk_0_S_in(prog_clk_1_wires[94]),
    .prog_clk_0_E_out(prog_clk_0_wires[187]),
    .prog_clk_0_S_out(prog_clk_0_wires[186]),
    .Test_en_W_out(Test_enWires[98]),
    .Test_en_E_in(Test_enWires[97]),
    .SC_OUT_BOT(scff_Wires[124]),
    .SC_IN_TOP(scff_Wires[123]),
    .top_width_0_height_0__pin_0_(cbx_1__1__47_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__47_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__47_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__47_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__47_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__47_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__47_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__47_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__47_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__47_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__47_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__47_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__47_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__47_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__47_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__47_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[47]),
    .right_width_0_height_0__pin_16_(cby_1__1__51_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__51_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__51_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__51_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__51_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__51_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__51_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__51_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__51_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__51_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__51_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__51_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__51_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__51_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__51_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__51_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__39_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_51_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_51_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_51_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_51_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_51_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_51_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_51_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_51_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_51_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_51_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_51_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_51_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_51_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_51_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_51_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_51_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_51_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_51_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_51_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_51_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_51_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_51_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_51_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_51_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_51_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_51_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_51_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_51_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_51_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_51_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_51_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_51_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[46]),
    .ccff_tail(grid_clb_51_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__5_
  (
    .clk_0_N_in(clk_1_wires[102]),
    .prog_clk_0_N_in(prog_clk_1_wires[102]),
    .prog_clk_0_E_out(prog_clk_0_wires[190]),
    .prog_clk_0_S_out(prog_clk_0_wires[189]),
    .Test_en_W_out(Test_enWires[120]),
    .Test_en_E_in(Test_enWires[119]),
    .SC_OUT_BOT(scff_Wires[122]),
    .SC_IN_TOP(scff_Wires[121]),
    .top_width_0_height_0__pin_0_(cbx_1__1__48_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__48_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__48_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__48_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__48_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__48_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__48_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__48_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__48_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__48_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__48_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__48_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__48_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__48_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__48_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__48_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[48]),
    .right_width_0_height_0__pin_16_(cby_1__1__52_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__52_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__52_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__52_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__52_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__52_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__52_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__52_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__52_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__52_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__52_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__52_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__52_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__52_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__52_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__52_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__40_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_52_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_52_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_52_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_52_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_52_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_52_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_52_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_52_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_52_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_52_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_52_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_52_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_52_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_52_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_52_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_52_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_52_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_52_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_52_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_52_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_52_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_52_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_52_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_52_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_52_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_52_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_52_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_52_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_52_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_52_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_52_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_52_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[47]),
    .ccff_tail(grid_clb_52_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__6_
  (
    .clk_0_S_in(clk_1_wires[101]),
    .prog_clk_0_S_in(prog_clk_1_wires[101]),
    .prog_clk_0_E_out(prog_clk_0_wires[193]),
    .prog_clk_0_S_out(prog_clk_0_wires[192]),
    .Test_en_W_out(Test_enWires[142]),
    .Test_en_E_in(Test_enWires[141]),
    .SC_OUT_BOT(scff_Wires[120]),
    .SC_IN_TOP(scff_Wires[119]),
    .top_width_0_height_0__pin_0_(cbx_1__1__49_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__49_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__49_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__49_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__49_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__49_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__49_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__49_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__49_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__49_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__49_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__49_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__49_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__49_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__49_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__49_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[49]),
    .right_width_0_height_0__pin_16_(cby_1__1__53_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__53_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__53_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__53_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__53_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__53_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__53_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__53_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__53_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__53_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__53_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__53_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__53_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__53_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__53_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__53_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__41_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_53_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_53_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_53_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_53_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_53_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_53_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_53_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_53_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_53_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_53_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_53_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_53_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_53_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_53_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_53_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_53_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_53_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_53_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_53_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_53_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_53_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_53_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_53_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_53_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_53_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_53_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_53_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_53_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_53_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_53_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_53_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_53_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[48]),
    .ccff_tail(grid_clb_53_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__7_
  (
    .clk_0_N_in(clk_1_wires[109]),
    .prog_clk_0_N_in(prog_clk_1_wires[109]),
    .prog_clk_0_E_out(prog_clk_0_wires[196]),
    .prog_clk_0_S_out(prog_clk_0_wires[195]),
    .Test_en_W_out(Test_enWires[164]),
    .Test_en_E_in(Test_enWires[163]),
    .SC_OUT_BOT(scff_Wires[118]),
    .SC_IN_TOP(scff_Wires[117]),
    .top_width_0_height_0__pin_0_(cbx_1__1__50_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__50_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__50_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__50_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__50_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__50_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__50_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__50_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__50_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__50_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__50_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__50_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__50_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__50_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__50_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__50_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[50]),
    .right_width_0_height_0__pin_16_(cby_1__1__54_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__54_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__54_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__54_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__54_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__54_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__54_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__54_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__54_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__54_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__54_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__54_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__54_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__54_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__54_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__54_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__42_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_54_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_54_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_54_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_54_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_54_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_54_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_54_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_54_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_54_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_54_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_54_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_54_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_54_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_54_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_54_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_54_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_54_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_54_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_54_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_54_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_54_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_54_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_54_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_54_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_54_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_54_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_54_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_54_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_54_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_54_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_54_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_54_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[49]),
    .ccff_tail(grid_clb_54_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__8_
  (
    .clk_0_S_in(clk_1_wires[108]),
    .prog_clk_0_S_in(prog_clk_1_wires[108]),
    .prog_clk_0_E_out(prog_clk_0_wires[199]),
    .prog_clk_0_S_out(prog_clk_0_wires[198]),
    .Test_en_W_out(Test_enWires[186]),
    .Test_en_E_in(Test_enWires[185]),
    .SC_OUT_BOT(scff_Wires[116]),
    .SC_IN_TOP(scff_Wires[115]),
    .top_width_0_height_0__pin_0_(cbx_1__1__51_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__51_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__51_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__51_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__51_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__51_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__51_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__51_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__51_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__51_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__51_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__51_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__51_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__51_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__51_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__51_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[51]),
    .right_width_0_height_0__pin_16_(cby_1__1__55_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__55_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__55_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__55_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__55_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__55_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__55_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__55_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__55_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__55_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__55_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__55_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__55_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__55_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__55_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__55_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__43_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_55_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_55_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_55_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_55_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_55_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_55_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_55_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_55_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_55_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_55_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_55_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_55_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_55_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_55_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_55_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_55_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_55_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_55_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_55_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_55_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_55_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_55_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_55_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_55_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_55_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_55_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_55_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_55_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_55_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_55_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_55_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_55_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[50]),
    .ccff_tail(grid_clb_55_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__9_
  (
    .clk_0_N_in(clk_1_wires[116]),
    .prog_clk_0_N_in(prog_clk_1_wires[116]),
    .prog_clk_0_E_out(prog_clk_0_wires[202]),
    .prog_clk_0_S_out(prog_clk_0_wires[201]),
    .Test_en_W_out(Test_enWires[208]),
    .Test_en_E_in(Test_enWires[207]),
    .SC_OUT_BOT(scff_Wires[114]),
    .SC_IN_TOP(scff_Wires[113]),
    .top_width_0_height_0__pin_0_(cbx_1__1__52_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__52_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__52_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__52_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__52_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__52_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__52_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__52_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__52_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__52_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__52_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__52_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__52_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__52_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__52_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__52_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[52]),
    .right_width_0_height_0__pin_16_(cby_1__1__56_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__56_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__56_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__56_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__56_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__56_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__56_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__56_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__56_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__56_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__56_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__56_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__56_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__56_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__56_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__56_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__44_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_56_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_56_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_56_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_56_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_56_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_56_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_56_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_56_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_56_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_56_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_56_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_56_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_56_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_56_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_56_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_56_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_56_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_56_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_56_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_56_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_56_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_56_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_56_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_56_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_56_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_56_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_56_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_56_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_56_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_56_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_56_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_56_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[51]),
    .ccff_tail(grid_clb_56_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__10_
  (
    .clk_0_S_in(clk_1_wires[115]),
    .prog_clk_0_S_in(prog_clk_1_wires[115]),
    .prog_clk_0_E_out(prog_clk_0_wires[205]),
    .prog_clk_0_S_out(prog_clk_0_wires[204]),
    .Test_en_W_out(Test_enWires[230]),
    .Test_en_E_in(Test_enWires[229]),
    .SC_OUT_BOT(scff_Wires[112]),
    .SC_IN_TOP(scff_Wires[111]),
    .top_width_0_height_0__pin_0_(cbx_1__1__53_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__53_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__53_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__53_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__53_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__53_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__53_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__53_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__53_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__53_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__53_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__53_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__53_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__53_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__53_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__53_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[53]),
    .right_width_0_height_0__pin_16_(cby_1__1__57_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__57_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__57_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__57_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__57_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__57_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__57_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__57_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__57_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__57_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__57_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__57_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__57_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__57_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__57_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__57_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__45_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_57_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_57_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_57_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_57_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_57_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_57_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_57_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_57_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_57_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_57_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_57_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_57_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_57_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_57_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_57_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_57_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_57_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_57_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_57_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_57_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_57_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_57_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_57_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_57_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_57_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_57_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_57_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_57_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_57_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_57_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_57_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_57_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[52]),
    .ccff_tail(grid_clb_57_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__11_
  (
    .clk_0_N_in(clk_1_wires[123]),
    .prog_clk_0_N_in(prog_clk_1_wires[123]),
    .prog_clk_0_E_out(prog_clk_0_wires[208]),
    .prog_clk_0_S_out(prog_clk_0_wires[207]),
    .Test_en_W_out(Test_enWires[252]),
    .Test_en_E_in(Test_enWires[251]),
    .SC_OUT_BOT(scff_Wires[110]),
    .SC_IN_TOP(scff_Wires[109]),
    .top_width_0_height_0__pin_0_(cbx_1__1__54_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__54_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__54_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__54_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__54_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__54_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__54_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__54_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__54_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__54_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__54_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__54_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__54_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__54_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__54_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__54_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[54]),
    .right_width_0_height_0__pin_16_(cby_1__1__58_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__58_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__58_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__58_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__58_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__58_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__58_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__58_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__58_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__58_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__58_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__58_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__58_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__58_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__58_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__58_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__46_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_58_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_58_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_58_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_58_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_58_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_58_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_58_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_58_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_58_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_58_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_58_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_58_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_58_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_58_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_58_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_58_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_58_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_58_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_58_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_58_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_58_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_58_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_58_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_58_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_58_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_58_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_58_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_58_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_58_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_58_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_58_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_58_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[53]),
    .ccff_tail(grid_clb_58_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__12_
  (
    .clk_0_S_in(clk_1_wires[122]),
    .prog_clk_0_S_in(prog_clk_1_wires[122]),
    .prog_clk_0_N_out(prog_clk_0_wires[213]),
    .prog_clk_0_E_out(prog_clk_0_wires[211]),
    .prog_clk_0_S_out(prog_clk_0_wires[210]),
    .Test_en_W_out(Test_enWires[274]),
    .Test_en_E_in(Test_enWires[273]),
    .SC_OUT_BOT(scff_Wires[108]),
    .SC_IN_TOP(scff_Wires[107]),
    .top_width_0_height_0__pin_0_(cbx_1__12__4_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__4_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__4_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__4_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__4_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__4_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__4_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__4_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__4_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__4_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__4_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__4_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__4_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__4_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__4_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__4_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_5__12__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__59_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__59_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__59_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__59_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__59_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__59_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__59_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__59_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__59_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__59_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__59_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__59_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__59_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__59_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__59_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__59_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__47_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_59_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_59_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_59_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_59_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_59_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_59_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_59_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_59_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_59_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_59_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_59_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_59_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_59_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_59_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_59_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_59_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_59_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_59_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_59_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_59_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_59_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_59_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_59_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_59_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_59_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_59_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_59_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_59_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_59_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_59_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_59_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_59_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[54]),
    .ccff_tail(grid_clb_59_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__1_
  (
    .clk_0_N_in(clk_1_wires[90]),
    .prog_clk_0_N_in(prog_clk_1_wires[90]),
    .prog_clk_0_E_out(prog_clk_0_wires[216]),
    .prog_clk_0_S_out(prog_clk_0_wires[215]),
    .Test_en_W_out(Test_enWires[34]),
    .Test_en_E_in(Test_enWires[33]),
    .SC_OUT_TOP(scff_Wires[135]),
    .SC_IN_BOT(scff_Wires[134]),
    .top_width_0_height_0__pin_0_(cbx_1__1__55_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__55_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__55_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__55_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__55_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__55_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__55_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__55_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__55_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__55_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__55_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__55_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__55_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__55_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__55_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__55_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[55]),
    .right_width_0_height_0__pin_16_(cby_1__1__60_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__60_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__60_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__60_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__60_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__60_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__60_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__60_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__60_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__60_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__60_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__60_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__60_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__60_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__60_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__60_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__48_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_60_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_60_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_60_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_60_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_60_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_60_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_60_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_60_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_60_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_60_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_60_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_60_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_60_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_60_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_60_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_60_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_60_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_60_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_60_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_60_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_60_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_60_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_60_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_60_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_60_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_60_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_60_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_60_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_60_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_60_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_60_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_60_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_6__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_60_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__2_
  (
    .clk_0_S_in(clk_1_wires[89]),
    .prog_clk_0_S_in(prog_clk_1_wires[89]),
    .prog_clk_0_E_out(prog_clk_0_wires[219]),
    .prog_clk_0_S_out(prog_clk_0_wires[218]),
    .Test_en_W_out(Test_enWires[56]),
    .Test_en_E_in(Test_enWires[55]),
    .SC_OUT_TOP(scff_Wires[137]),
    .SC_IN_BOT(scff_Wires[136]),
    .top_width_0_height_0__pin_0_(cbx_1__1__56_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__56_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__56_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__56_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__56_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__56_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__56_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__56_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__56_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__56_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__56_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__56_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__56_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__56_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__56_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__56_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[56]),
    .right_width_0_height_0__pin_16_(cby_1__1__61_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__61_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__61_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__61_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__61_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__61_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__61_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__61_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__61_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__61_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__61_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__61_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__61_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__61_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__61_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__61_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__49_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_61_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_61_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_61_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_61_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_61_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_61_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_61_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_61_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_61_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_61_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_61_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_61_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_61_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_61_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_61_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_61_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_61_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_61_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_61_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_61_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_61_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_61_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_61_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_61_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_61_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_61_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_61_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_61_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_61_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_61_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_61_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_61_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[55]),
    .ccff_tail(grid_clb_61_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__3_
  (
    .clk_0_N_in(clk_1_wires[97]),
    .prog_clk_0_N_in(prog_clk_1_wires[97]),
    .prog_clk_0_E_out(prog_clk_0_wires[222]),
    .prog_clk_0_S_out(prog_clk_0_wires[221]),
    .Test_en_W_out(Test_enWires[78]),
    .Test_en_E_in(Test_enWires[77]),
    .SC_OUT_TOP(scff_Wires[139]),
    .SC_IN_BOT(scff_Wires[138]),
    .top_width_0_height_0__pin_0_(cbx_1__1__57_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__57_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__57_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__57_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__57_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__57_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__57_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__57_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__57_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__57_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__57_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__57_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__57_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__57_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__57_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__57_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[57]),
    .right_width_0_height_0__pin_16_(cby_1__1__62_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__62_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__62_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__62_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__62_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__62_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__62_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__62_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__62_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__62_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__62_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__62_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__62_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__62_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__62_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__62_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__50_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_62_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_62_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_62_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_62_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_62_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_62_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_62_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_62_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_62_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_62_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_62_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_62_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_62_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_62_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_62_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_62_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_62_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_62_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_62_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_62_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_62_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_62_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_62_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_62_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_62_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_62_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_62_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_62_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_62_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_62_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_62_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_62_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[56]),
    .ccff_tail(grid_clb_62_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__4_
  (
    .clk_0_S_in(clk_1_wires[96]),
    .prog_clk_0_S_in(prog_clk_1_wires[96]),
    .prog_clk_0_E_out(prog_clk_0_wires[225]),
    .prog_clk_0_S_out(prog_clk_0_wires[224]),
    .Test_en_W_out(Test_enWires[100]),
    .Test_en_E_in(Test_enWires[99]),
    .SC_OUT_TOP(scff_Wires[141]),
    .SC_IN_BOT(scff_Wires[140]),
    .top_width_0_height_0__pin_0_(cbx_1__1__58_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__58_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__58_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__58_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__58_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__58_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__58_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__58_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__58_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__58_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__58_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__58_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__58_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__58_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__58_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__58_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[58]),
    .right_width_0_height_0__pin_16_(cby_1__1__63_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__63_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__63_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__63_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__63_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__63_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__63_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__63_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__63_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__63_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__63_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__63_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__63_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__63_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__63_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__63_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__51_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_63_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_63_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_63_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_63_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_63_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_63_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_63_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_63_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_63_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_63_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_63_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_63_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_63_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_63_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_63_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_63_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_63_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_63_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_63_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_63_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_63_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_63_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_63_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_63_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_63_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_63_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_63_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_63_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_63_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_63_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_63_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_63_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[57]),
    .ccff_tail(grid_clb_63_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__5_
  (
    .clk_0_N_in(clk_1_wires[104]),
    .prog_clk_0_N_in(prog_clk_1_wires[104]),
    .prog_clk_0_E_out(prog_clk_0_wires[228]),
    .prog_clk_0_S_out(prog_clk_0_wires[227]),
    .Test_en_W_out(Test_enWires[122]),
    .Test_en_E_in(Test_enWires[121]),
    .SC_OUT_TOP(scff_Wires[143]),
    .SC_IN_BOT(scff_Wires[142]),
    .top_width_0_height_0__pin_0_(cbx_1__1__59_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__59_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__59_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__59_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__59_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__59_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__59_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__59_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__59_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__59_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__59_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__59_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__59_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__59_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__59_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__59_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[59]),
    .right_width_0_height_0__pin_16_(cby_1__1__64_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__64_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__64_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__64_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__64_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__64_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__64_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__64_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__64_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__64_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__64_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__64_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__64_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__64_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__64_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__64_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__52_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_64_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_64_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_64_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_64_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_64_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_64_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_64_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_64_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_64_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_64_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_64_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_64_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_64_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_64_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_64_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_64_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_64_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_64_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_64_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_64_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_64_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_64_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_64_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_64_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_64_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_64_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_64_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_64_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_64_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_64_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_64_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_64_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[58]),
    .ccff_tail(grid_clb_64_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__6_
  (
    .clk_0_S_in(clk_1_wires[103]),
    .prog_clk_0_S_in(prog_clk_1_wires[103]),
    .prog_clk_0_E_out(prog_clk_0_wires[231]),
    .prog_clk_0_S_out(prog_clk_0_wires[230]),
    .Test_en_W_out(Test_enWires[144]),
    .Test_en_E_in(Test_enWires[143]),
    .SC_OUT_TOP(scff_Wires[145]),
    .SC_IN_BOT(scff_Wires[144]),
    .top_width_0_height_0__pin_0_(cbx_1__1__60_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__60_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__60_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__60_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__60_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__60_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__60_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__60_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__60_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__60_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__60_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__60_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__60_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__60_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__60_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__60_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[60]),
    .right_width_0_height_0__pin_16_(cby_1__1__65_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__65_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__65_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__65_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__65_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__65_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__65_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__65_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__65_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__65_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__65_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__65_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__65_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__65_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__65_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__65_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__53_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_65_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_65_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_65_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_65_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_65_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_65_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_65_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_65_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_65_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_65_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_65_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_65_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_65_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_65_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_65_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_65_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_65_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_65_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_65_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_65_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_65_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_65_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_65_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_65_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_65_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_65_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_65_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_65_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_65_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_65_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_65_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_65_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[59]),
    .ccff_tail(grid_clb_65_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__7_
  (
    .clk_0_N_in(clk_1_wires[111]),
    .prog_clk_0_N_in(prog_clk_1_wires[111]),
    .prog_clk_0_E_out(prog_clk_0_wires[234]),
    .prog_clk_0_S_out(prog_clk_0_wires[233]),
    .Test_en_W_out(Test_enWires[166]),
    .Test_en_E_in(Test_enWires[165]),
    .SC_OUT_TOP(scff_Wires[147]),
    .SC_IN_BOT(scff_Wires[146]),
    .top_width_0_height_0__pin_0_(cbx_1__1__61_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__61_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__61_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__61_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__61_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__61_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__61_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__61_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__61_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__61_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__61_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__61_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__61_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__61_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__61_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__61_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[61]),
    .right_width_0_height_0__pin_16_(cby_1__1__66_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__66_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__66_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__66_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__66_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__66_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__66_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__66_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__66_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__66_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__66_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__66_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__66_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__66_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__66_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__66_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__54_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_66_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_66_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_66_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_66_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_66_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_66_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_66_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_66_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_66_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_66_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_66_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_66_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_66_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_66_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_66_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_66_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_66_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_66_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_66_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_66_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_66_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_66_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_66_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_66_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_66_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_66_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_66_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_66_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_66_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_66_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_66_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_66_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[60]),
    .ccff_tail(grid_clb_66_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__8_
  (
    .clk_0_S_in(clk_1_wires[110]),
    .prog_clk_0_S_in(prog_clk_1_wires[110]),
    .prog_clk_0_E_out(prog_clk_0_wires[237]),
    .prog_clk_0_S_out(prog_clk_0_wires[236]),
    .Test_en_W_out(Test_enWires[188]),
    .Test_en_E_in(Test_enWires[187]),
    .SC_OUT_TOP(scff_Wires[149]),
    .SC_IN_BOT(scff_Wires[148]),
    .top_width_0_height_0__pin_0_(cbx_1__1__62_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__62_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__62_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__62_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__62_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__62_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__62_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__62_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__62_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__62_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__62_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__62_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__62_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__62_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__62_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__62_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[62]),
    .right_width_0_height_0__pin_16_(cby_1__1__67_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__67_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__67_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__67_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__67_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__67_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__67_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__67_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__67_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__67_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__67_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__67_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__67_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__67_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__67_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__67_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__55_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_67_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_67_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_67_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_67_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_67_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_67_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_67_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_67_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_67_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_67_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_67_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_67_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_67_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_67_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_67_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_67_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_67_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_67_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_67_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_67_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_67_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_67_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_67_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_67_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_67_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_67_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_67_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_67_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_67_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_67_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_67_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_67_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[61]),
    .ccff_tail(grid_clb_67_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__9_
  (
    .clk_0_N_in(clk_1_wires[118]),
    .prog_clk_0_N_in(prog_clk_1_wires[118]),
    .prog_clk_0_E_out(prog_clk_0_wires[240]),
    .prog_clk_0_S_out(prog_clk_0_wires[239]),
    .Test_en_W_out(Test_enWires[210]),
    .Test_en_E_in(Test_enWires[209]),
    .SC_OUT_TOP(scff_Wires[151]),
    .SC_IN_BOT(scff_Wires[150]),
    .top_width_0_height_0__pin_0_(cbx_1__1__63_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__63_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__63_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__63_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__63_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__63_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__63_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__63_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__63_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__63_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__63_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__63_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__63_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__63_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__63_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__63_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[63]),
    .right_width_0_height_0__pin_16_(cby_1__1__68_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__68_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__68_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__68_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__68_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__68_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__68_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__68_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__68_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__68_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__68_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__68_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__68_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__68_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__68_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__68_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__56_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_68_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_68_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_68_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_68_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_68_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_68_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_68_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_68_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_68_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_68_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_68_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_68_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_68_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_68_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_68_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_68_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_68_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_68_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_68_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_68_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_68_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_68_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_68_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_68_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_68_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_68_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_68_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_68_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_68_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_68_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_68_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_68_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[62]),
    .ccff_tail(grid_clb_68_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__10_
  (
    .clk_0_S_in(clk_1_wires[117]),
    .prog_clk_0_S_in(prog_clk_1_wires[117]),
    .prog_clk_0_E_out(prog_clk_0_wires[243]),
    .prog_clk_0_S_out(prog_clk_0_wires[242]),
    .Test_en_W_out(Test_enWires[232]),
    .Test_en_E_in(Test_enWires[231]),
    .SC_OUT_TOP(scff_Wires[153]),
    .SC_IN_BOT(scff_Wires[152]),
    .top_width_0_height_0__pin_0_(cbx_1__1__64_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__64_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__64_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__64_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__64_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__64_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__64_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__64_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__64_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__64_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__64_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__64_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__64_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__64_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__64_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__64_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[64]),
    .right_width_0_height_0__pin_16_(cby_1__1__69_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__69_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__69_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__69_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__69_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__69_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__69_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__69_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__69_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__69_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__69_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__69_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__69_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__69_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__69_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__69_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__57_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_69_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_69_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_69_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_69_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_69_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_69_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_69_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_69_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_69_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_69_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_69_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_69_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_69_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_69_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_69_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_69_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_69_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_69_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_69_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_69_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_69_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_69_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_69_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_69_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_69_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_69_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_69_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_69_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_69_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_69_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_69_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_69_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[63]),
    .ccff_tail(grid_clb_69_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__11_
  (
    .clk_0_N_in(clk_1_wires[125]),
    .prog_clk_0_N_in(prog_clk_1_wires[125]),
    .prog_clk_0_E_out(prog_clk_0_wires[246]),
    .prog_clk_0_S_out(prog_clk_0_wires[245]),
    .Test_en_W_out(Test_enWires[254]),
    .Test_en_E_in(Test_enWires[253]),
    .SC_OUT_TOP(scff_Wires[155]),
    .SC_IN_BOT(scff_Wires[154]),
    .top_width_0_height_0__pin_0_(cbx_1__1__65_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__65_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__65_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__65_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__65_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__65_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__65_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__65_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__65_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__65_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__65_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__65_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__65_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__65_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__65_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__65_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[65]),
    .right_width_0_height_0__pin_16_(cby_1__1__70_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__70_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__70_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__70_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__70_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__70_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__70_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__70_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__70_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__70_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__70_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__70_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__70_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__70_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__70_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__70_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__58_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_70_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_70_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_70_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_70_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_70_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_70_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_70_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_70_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_70_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_70_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_70_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_70_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_70_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_70_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_70_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_70_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_70_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_70_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_70_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_70_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_70_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_70_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_70_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_70_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_70_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_70_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_70_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_70_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_70_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_70_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_70_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_70_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[64]),
    .ccff_tail(grid_clb_70_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__12_
  (
    .clk_0_S_in(clk_1_wires[124]),
    .prog_clk_0_S_in(prog_clk_1_wires[124]),
    .prog_clk_0_N_out(prog_clk_0_wires[251]),
    .prog_clk_0_E_out(prog_clk_0_wires[249]),
    .prog_clk_0_S_out(prog_clk_0_wires[248]),
    .Test_en_W_out(Test_enWires[276]),
    .Test_en_E_in(Test_enWires[275]),
    .SC_OUT_TOP(scff_Wires[157]),
    .SC_IN_BOT(scff_Wires[156]),
    .top_width_0_height_0__pin_0_(cbx_1__12__5_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__5_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__5_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__5_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__5_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__5_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__5_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__5_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__5_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__5_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__5_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__5_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__5_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__5_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__5_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__5_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_6__12__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__71_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__71_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__71_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__71_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__71_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__71_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__71_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__71_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__71_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__71_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__71_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__71_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__71_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__71_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__71_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__71_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__59_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_71_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_71_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_71_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_71_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_71_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_71_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_71_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_71_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_71_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_71_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_71_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_71_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_71_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_71_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_71_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_71_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_71_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_71_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_71_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_71_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_71_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_71_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_71_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_71_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_71_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_71_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_71_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_71_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_71_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_71_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_71_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_71_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[65]),
    .ccff_tail(grid_clb_71_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__1_
  (
    .clk_0_N_in(clk_1_wires[130]),
    .prog_clk_0_N_in(prog_clk_1_wires[130]),
    .prog_clk_0_E_out(prog_clk_0_wires[254]),
    .prog_clk_0_S_out(prog_clk_0_wires[253]),
    .Test_en_E_out(Test_enWires[36]),
    .Test_en_W_in(Test_enWires[35]),
    .SC_OUT_BOT(scff_Wires[184]),
    .SC_IN_TOP(scff_Wires[182]),
    .top_width_0_height_0__pin_0_(cbx_1__1__66_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__66_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__66_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__66_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__66_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__66_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__66_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__66_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__66_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__66_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__66_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__66_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__66_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__66_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__66_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__66_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[66]),
    .right_width_0_height_0__pin_16_(cby_1__1__72_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__72_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__72_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__72_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__72_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__72_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__72_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__72_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__72_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__72_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__72_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__72_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__72_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__72_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__72_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__72_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__60_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_72_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_72_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_72_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_72_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_72_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_72_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_72_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_72_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_72_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_72_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_72_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_72_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_72_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_72_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_72_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_72_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_72_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_72_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_72_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_72_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_72_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_72_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_72_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_72_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_72_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_72_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_72_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_72_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_72_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_72_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_72_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_72_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_7__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_72_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__2_
  (
    .clk_0_S_in(clk_1_wires[129]),
    .prog_clk_0_S_in(prog_clk_1_wires[129]),
    .prog_clk_0_E_out(prog_clk_0_wires[257]),
    .prog_clk_0_S_out(prog_clk_0_wires[256]),
    .Test_en_E_out(Test_enWires[58]),
    .Test_en_W_in(Test_enWires[57]),
    .SC_OUT_BOT(scff_Wires[181]),
    .SC_IN_TOP(scff_Wires[180]),
    .top_width_0_height_0__pin_0_(cbx_1__1__67_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__67_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__67_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__67_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__67_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__67_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__67_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__67_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__67_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__67_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__67_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__67_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__67_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__67_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__67_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__67_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[67]),
    .right_width_0_height_0__pin_16_(cby_1__1__73_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__73_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__73_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__73_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__73_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__73_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__73_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__73_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__73_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__73_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__73_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__73_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__73_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__73_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__73_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__73_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__61_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_73_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_73_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_73_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_73_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_73_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_73_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_73_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_73_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_73_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_73_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_73_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_73_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_73_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_73_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_73_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_73_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_73_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_73_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_73_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_73_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_73_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_73_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_73_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_73_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_73_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_73_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_73_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_73_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_73_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_73_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_73_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_73_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[66]),
    .ccff_tail(grid_clb_73_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__3_
  (
    .clk_0_N_in(clk_1_wires[137]),
    .prog_clk_0_N_in(prog_clk_1_wires[137]),
    .prog_clk_0_E_out(prog_clk_0_wires[260]),
    .prog_clk_0_S_out(prog_clk_0_wires[259]),
    .Test_en_E_out(Test_enWires[80]),
    .Test_en_W_in(Test_enWires[79]),
    .SC_OUT_BOT(scff_Wires[179]),
    .SC_IN_TOP(scff_Wires[178]),
    .top_width_0_height_0__pin_0_(cbx_1__1__68_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__68_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__68_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__68_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__68_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__68_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__68_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__68_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__68_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__68_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__68_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__68_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__68_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__68_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__68_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__68_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[68]),
    .right_width_0_height_0__pin_16_(cby_1__1__74_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__74_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__74_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__74_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__74_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__74_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__74_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__74_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__74_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__74_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__74_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__74_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__74_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__74_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__74_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__74_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__62_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_74_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_74_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_74_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_74_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_74_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_74_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_74_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_74_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_74_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_74_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_74_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_74_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_74_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_74_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_74_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_74_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_74_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_74_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_74_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_74_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_74_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_74_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_74_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_74_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_74_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_74_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_74_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_74_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_74_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_74_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_74_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_74_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[67]),
    .ccff_tail(grid_clb_74_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__4_
  (
    .clk_0_S_in(clk_1_wires[136]),
    .prog_clk_0_S_in(prog_clk_1_wires[136]),
    .prog_clk_0_E_out(prog_clk_0_wires[263]),
    .prog_clk_0_S_out(prog_clk_0_wires[262]),
    .Test_en_E_out(Test_enWires[102]),
    .Test_en_W_in(Test_enWires[101]),
    .SC_OUT_BOT(scff_Wires[177]),
    .SC_IN_TOP(scff_Wires[176]),
    .top_width_0_height_0__pin_0_(cbx_1__1__69_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__69_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__69_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__69_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__69_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__69_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__69_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__69_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__69_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__69_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__69_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__69_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__69_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__69_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__69_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__69_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[69]),
    .right_width_0_height_0__pin_16_(cby_1__1__75_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__75_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__75_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__75_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__75_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__75_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__75_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__75_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__75_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__75_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__75_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__75_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__75_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__75_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__75_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__75_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__63_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_75_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_75_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_75_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_75_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_75_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_75_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_75_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_75_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_75_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_75_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_75_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_75_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_75_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_75_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_75_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_75_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_75_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_75_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_75_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_75_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_75_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_75_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_75_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_75_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_75_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_75_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_75_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_75_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_75_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_75_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_75_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_75_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[68]),
    .ccff_tail(grid_clb_75_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__5_
  (
    .clk_0_N_in(clk_1_wires[144]),
    .prog_clk_0_N_in(prog_clk_1_wires[144]),
    .prog_clk_0_E_out(prog_clk_0_wires[266]),
    .prog_clk_0_S_out(prog_clk_0_wires[265]),
    .Test_en_E_out(Test_enWires[124]),
    .Test_en_W_in(Test_enWires[123]),
    .SC_OUT_BOT(scff_Wires[175]),
    .SC_IN_TOP(scff_Wires[174]),
    .top_width_0_height_0__pin_0_(cbx_1__1__70_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__70_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__70_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__70_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__70_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__70_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__70_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__70_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__70_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__70_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__70_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__70_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__70_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__70_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__70_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__70_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[70]),
    .right_width_0_height_0__pin_16_(cby_1__1__76_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__76_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__76_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__76_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__76_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__76_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__76_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__76_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__76_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__76_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__76_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__76_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__76_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__76_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__76_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__76_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__64_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_76_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_76_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_76_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_76_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_76_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_76_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_76_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_76_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_76_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_76_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_76_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_76_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_76_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_76_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_76_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_76_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_76_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_76_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_76_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_76_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_76_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_76_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_76_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_76_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_76_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_76_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_76_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_76_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_76_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_76_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_76_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_76_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[69]),
    .ccff_tail(grid_clb_76_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__6_
  (
    .clk_0_S_in(clk_1_wires[143]),
    .prog_clk_0_S_in(prog_clk_1_wires[143]),
    .prog_clk_0_E_out(prog_clk_0_wires[269]),
    .prog_clk_0_S_out(prog_clk_0_wires[268]),
    .Test_en_E_out(Test_enWires[146]),
    .Test_en_W_in(Test_enWires[145]),
    .SC_OUT_BOT(scff_Wires[173]),
    .SC_IN_TOP(scff_Wires[172]),
    .top_width_0_height_0__pin_0_(cbx_1__1__71_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__71_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__71_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__71_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__71_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__71_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__71_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__71_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__71_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__71_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__71_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__71_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__71_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__71_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__71_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__71_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[71]),
    .right_width_0_height_0__pin_16_(cby_1__1__77_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__77_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__77_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__77_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__77_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__77_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__77_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__77_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__77_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__77_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__77_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__77_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__77_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__77_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__77_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__77_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__65_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_77_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_77_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_77_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_77_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_77_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_77_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_77_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_77_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_77_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_77_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_77_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_77_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_77_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_77_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_77_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_77_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_77_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_77_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_77_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_77_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_77_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_77_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_77_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_77_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_77_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_77_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_77_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_77_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_77_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_77_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_77_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_77_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[70]),
    .ccff_tail(grid_clb_77_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__7_
  (
    .clk_0_N_in(clk_1_wires[151]),
    .prog_clk_0_N_in(prog_clk_1_wires[151]),
    .prog_clk_0_E_out(prog_clk_0_wires[272]),
    .prog_clk_0_S_out(prog_clk_0_wires[271]),
    .Test_en_E_out(Test_enWires[168]),
    .Test_en_W_in(Test_enWires[167]),
    .SC_OUT_BOT(scff_Wires[171]),
    .SC_IN_TOP(scff_Wires[170]),
    .top_width_0_height_0__pin_0_(cbx_1__1__72_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__72_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__72_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__72_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__72_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__72_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__72_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__72_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__72_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__72_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__72_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__72_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__72_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__72_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__72_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__72_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[72]),
    .right_width_0_height_0__pin_16_(cby_1__1__78_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__78_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__78_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__78_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__78_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__78_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__78_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__78_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__78_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__78_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__78_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__78_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__78_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__78_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__78_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__78_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__66_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_78_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_78_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_78_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_78_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_78_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_78_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_78_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_78_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_78_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_78_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_78_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_78_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_78_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_78_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_78_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_78_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_78_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_78_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_78_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_78_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_78_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_78_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_78_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_78_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_78_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_78_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_78_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_78_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_78_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_78_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_78_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_78_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[71]),
    .ccff_tail(grid_clb_78_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__8_
  (
    .clk_0_S_in(clk_1_wires[150]),
    .prog_clk_0_S_in(prog_clk_1_wires[150]),
    .prog_clk_0_E_out(prog_clk_0_wires[275]),
    .prog_clk_0_S_out(prog_clk_0_wires[274]),
    .Test_en_E_out(Test_enWires[190]),
    .Test_en_W_in(Test_enWires[189]),
    .SC_OUT_BOT(scff_Wires[169]),
    .SC_IN_TOP(scff_Wires[168]),
    .top_width_0_height_0__pin_0_(cbx_1__1__73_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__73_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__73_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__73_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__73_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__73_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__73_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__73_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__73_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__73_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__73_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__73_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__73_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__73_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__73_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__73_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[73]),
    .right_width_0_height_0__pin_16_(cby_1__1__79_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__79_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__79_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__79_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__79_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__79_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__79_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__79_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__79_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__79_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__79_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__79_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__79_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__79_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__79_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__79_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__67_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_79_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_79_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_79_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_79_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_79_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_79_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_79_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_79_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_79_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_79_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_79_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_79_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_79_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_79_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_79_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_79_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_79_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_79_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_79_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_79_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_79_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_79_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_79_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_79_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_79_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_79_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_79_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_79_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_79_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_79_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_79_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_79_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[72]),
    .ccff_tail(grid_clb_79_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__9_
  (
    .clk_0_N_in(clk_1_wires[158]),
    .prog_clk_0_N_in(prog_clk_1_wires[158]),
    .prog_clk_0_E_out(prog_clk_0_wires[278]),
    .prog_clk_0_S_out(prog_clk_0_wires[277]),
    .Test_en_E_out(Test_enWires[212]),
    .Test_en_W_in(Test_enWires[211]),
    .SC_OUT_BOT(scff_Wires[167]),
    .SC_IN_TOP(scff_Wires[166]),
    .top_width_0_height_0__pin_0_(cbx_1__1__74_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__74_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__74_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__74_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__74_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__74_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__74_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__74_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__74_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__74_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__74_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__74_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__74_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__74_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__74_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__74_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[74]),
    .right_width_0_height_0__pin_16_(cby_1__1__80_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__80_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__80_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__80_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__80_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__80_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__80_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__80_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__80_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__80_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__80_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__80_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__80_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__80_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__80_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__80_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__68_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_80_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_80_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_80_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_80_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_80_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_80_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_80_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_80_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_80_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_80_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_80_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_80_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_80_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_80_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_80_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_80_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_80_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_80_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_80_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_80_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_80_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_80_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_80_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_80_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_80_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_80_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_80_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_80_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_80_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_80_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_80_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_80_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[73]),
    .ccff_tail(grid_clb_80_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__10_
  (
    .clk_0_S_in(clk_1_wires[157]),
    .prog_clk_0_S_in(prog_clk_1_wires[157]),
    .prog_clk_0_E_out(prog_clk_0_wires[281]),
    .prog_clk_0_S_out(prog_clk_0_wires[280]),
    .Test_en_E_out(Test_enWires[234]),
    .Test_en_W_in(Test_enWires[233]),
    .SC_OUT_BOT(scff_Wires[165]),
    .SC_IN_TOP(scff_Wires[164]),
    .top_width_0_height_0__pin_0_(cbx_1__1__75_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__75_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__75_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__75_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__75_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__75_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__75_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__75_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__75_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__75_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__75_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__75_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__75_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__75_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__75_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__75_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[75]),
    .right_width_0_height_0__pin_16_(cby_1__1__81_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__81_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__81_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__81_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__81_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__81_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__81_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__81_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__81_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__81_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__81_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__81_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__81_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__81_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__81_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__81_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__69_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_81_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_81_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_81_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_81_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_81_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_81_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_81_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_81_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_81_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_81_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_81_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_81_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_81_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_81_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_81_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_81_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_81_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_81_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_81_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_81_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_81_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_81_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_81_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_81_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_81_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_81_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_81_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_81_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_81_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_81_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_81_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_81_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[74]),
    .ccff_tail(grid_clb_81_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__11_
  (
    .clk_0_N_in(clk_1_wires[165]),
    .prog_clk_0_N_in(prog_clk_1_wires[165]),
    .prog_clk_0_E_out(prog_clk_0_wires[284]),
    .prog_clk_0_S_out(prog_clk_0_wires[283]),
    .Test_en_E_out(Test_enWires[256]),
    .Test_en_W_in(Test_enWires[255]),
    .SC_OUT_BOT(scff_Wires[163]),
    .SC_IN_TOP(scff_Wires[162]),
    .top_width_0_height_0__pin_0_(cbx_1__1__76_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__76_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__76_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__76_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__76_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__76_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__76_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__76_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__76_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__76_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__76_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__76_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__76_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__76_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__76_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__76_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[76]),
    .right_width_0_height_0__pin_16_(cby_1__1__82_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__82_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__82_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__82_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__82_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__82_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__82_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__82_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__82_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__82_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__82_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__82_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__82_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__82_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__82_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__82_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__70_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_82_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_82_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_82_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_82_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_82_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_82_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_82_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_82_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_82_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_82_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_82_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_82_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_82_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_82_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_82_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_82_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_82_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_82_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_82_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_82_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_82_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_82_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_82_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_82_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_82_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_82_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_82_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_82_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_82_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_82_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_82_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_82_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[75]),
    .ccff_tail(grid_clb_82_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__12_
  (
    .clk_0_S_in(clk_1_wires[164]),
    .prog_clk_0_S_in(prog_clk_1_wires[164]),
    .prog_clk_0_N_out(prog_clk_0_wires[289]),
    .prog_clk_0_E_out(prog_clk_0_wires[287]),
    .prog_clk_0_S_out(prog_clk_0_wires[286]),
    .Test_en_E_out(Test_enWires[278]),
    .Test_en_W_in(Test_enWires[277]),
    .SC_OUT_BOT(scff_Wires[161]),
    .SC_IN_TOP(scff_Wires[160]),
    .top_width_0_height_0__pin_0_(cbx_1__12__6_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__6_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__6_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__6_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__6_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__6_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__6_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__6_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__6_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__6_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__6_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__6_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__6_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__6_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__6_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__6_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_7__12__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__83_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__83_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__83_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__83_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__83_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__83_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__83_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__83_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__83_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__83_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__83_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__83_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__83_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__83_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__83_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__83_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__71_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_83_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_83_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_83_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_83_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_83_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_83_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_83_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_83_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_83_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_83_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_83_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_83_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_83_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_83_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_83_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_83_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_83_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_83_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_83_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_83_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_83_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_83_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_83_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_83_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_83_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_83_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_83_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_83_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_83_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_83_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_83_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_83_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[76]),
    .ccff_tail(grid_clb_83_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__1_
  (
    .clk_0_N_in(clk_1_wires[132]),
    .prog_clk_0_N_in(prog_clk_1_wires[132]),
    .prog_clk_0_E_out(prog_clk_0_wires[292]),
    .prog_clk_0_S_out(prog_clk_0_wires[291]),
    .Test_en_E_out(Test_enWires[38]),
    .Test_en_W_in(Test_enWires[37]),
    .SC_OUT_TOP(scff_Wires[188]),
    .SC_IN_BOT(scff_Wires[187]),
    .top_width_0_height_0__pin_0_(cbx_1__1__77_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__77_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__77_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__77_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__77_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__77_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__77_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__77_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__77_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__77_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__77_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__77_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__77_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__77_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__77_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__77_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[77]),
    .right_width_0_height_0__pin_16_(cby_1__1__84_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__84_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__84_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__84_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__84_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__84_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__84_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__84_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__84_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__84_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__84_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__84_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__84_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__84_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__84_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__84_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__72_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_84_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_84_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_84_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_84_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_84_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_84_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_84_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_84_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_84_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_84_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_84_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_84_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_84_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_84_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_84_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_84_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_84_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_84_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_84_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_84_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_84_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_84_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_84_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_84_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_84_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_84_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_84_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_84_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_84_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_84_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_84_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_84_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_8__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_84_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__2_
  (
    .clk_0_S_in(clk_1_wires[131]),
    .prog_clk_0_S_in(prog_clk_1_wires[131]),
    .prog_clk_0_E_out(prog_clk_0_wires[295]),
    .prog_clk_0_S_out(prog_clk_0_wires[294]),
    .Test_en_E_out(Test_enWires[60]),
    .Test_en_W_in(Test_enWires[59]),
    .SC_OUT_TOP(scff_Wires[190]),
    .SC_IN_BOT(scff_Wires[189]),
    .top_width_0_height_0__pin_0_(cbx_1__1__78_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__78_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__78_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__78_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__78_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__78_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__78_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__78_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__78_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__78_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__78_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__78_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__78_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__78_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__78_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__78_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[78]),
    .right_width_0_height_0__pin_16_(cby_1__1__85_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__85_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__85_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__85_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__85_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__85_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__85_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__85_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__85_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__85_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__85_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__85_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__85_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__85_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__85_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__85_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__73_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_85_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_85_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_85_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_85_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_85_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_85_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_85_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_85_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_85_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_85_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_85_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_85_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_85_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_85_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_85_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_85_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_85_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_85_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_85_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_85_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_85_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_85_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_85_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_85_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_85_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_85_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_85_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_85_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_85_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_85_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_85_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_85_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[77]),
    .ccff_tail(grid_clb_85_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__3_
  (
    .clk_0_N_in(clk_1_wires[139]),
    .prog_clk_0_N_in(prog_clk_1_wires[139]),
    .prog_clk_0_E_out(prog_clk_0_wires[298]),
    .prog_clk_0_S_out(prog_clk_0_wires[297]),
    .Test_en_E_out(Test_enWires[82]),
    .Test_en_W_in(Test_enWires[81]),
    .SC_OUT_TOP(scff_Wires[192]),
    .SC_IN_BOT(scff_Wires[191]),
    .top_width_0_height_0__pin_0_(cbx_1__1__79_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__79_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__79_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__79_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__79_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__79_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__79_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__79_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__79_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__79_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__79_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__79_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__79_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__79_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__79_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__79_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[79]),
    .right_width_0_height_0__pin_16_(cby_1__1__86_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__86_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__86_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__86_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__86_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__86_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__86_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__86_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__86_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__86_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__86_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__86_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__86_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__86_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__86_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__86_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__74_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_86_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_86_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_86_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_86_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_86_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_86_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_86_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_86_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_86_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_86_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_86_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_86_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_86_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_86_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_86_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_86_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_86_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_86_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_86_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_86_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_86_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_86_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_86_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_86_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_86_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_86_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_86_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_86_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_86_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_86_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_86_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_86_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[78]),
    .ccff_tail(grid_clb_86_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__4_
  (
    .clk_0_S_in(clk_1_wires[138]),
    .prog_clk_0_S_in(prog_clk_1_wires[138]),
    .prog_clk_0_E_out(prog_clk_0_wires[301]),
    .prog_clk_0_S_out(prog_clk_0_wires[300]),
    .Test_en_E_out(Test_enWires[104]),
    .Test_en_W_in(Test_enWires[103]),
    .SC_OUT_TOP(scff_Wires[194]),
    .SC_IN_BOT(scff_Wires[193]),
    .top_width_0_height_0__pin_0_(cbx_1__1__80_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__80_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__80_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__80_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__80_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__80_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__80_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__80_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__80_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__80_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__80_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__80_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__80_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__80_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__80_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__80_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[80]),
    .right_width_0_height_0__pin_16_(cby_1__1__87_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__87_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__87_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__87_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__87_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__87_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__87_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__87_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__87_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__87_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__87_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__87_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__87_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__87_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__87_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__87_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__75_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_87_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_87_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_87_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_87_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_87_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_87_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_87_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_87_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_87_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_87_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_87_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_87_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_87_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_87_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_87_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_87_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_87_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_87_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_87_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_87_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_87_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_87_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_87_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_87_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_87_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_87_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_87_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_87_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_87_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_87_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_87_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_87_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[79]),
    .ccff_tail(grid_clb_87_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__5_
  (
    .clk_0_N_in(clk_1_wires[146]),
    .prog_clk_0_N_in(prog_clk_1_wires[146]),
    .prog_clk_0_E_out(prog_clk_0_wires[304]),
    .prog_clk_0_S_out(prog_clk_0_wires[303]),
    .Test_en_E_out(Test_enWires[126]),
    .Test_en_W_in(Test_enWires[125]),
    .SC_OUT_TOP(scff_Wires[196]),
    .SC_IN_BOT(scff_Wires[195]),
    .top_width_0_height_0__pin_0_(cbx_1__1__81_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__81_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__81_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__81_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__81_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__81_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__81_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__81_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__81_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__81_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__81_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__81_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__81_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__81_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__81_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__81_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[81]),
    .right_width_0_height_0__pin_16_(cby_1__1__88_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__88_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__88_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__88_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__88_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__88_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__88_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__88_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__88_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__88_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__88_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__88_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__88_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__88_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__88_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__88_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__76_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_88_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_88_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_88_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_88_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_88_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_88_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_88_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_88_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_88_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_88_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_88_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_88_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_88_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_88_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_88_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_88_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_88_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_88_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_88_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_88_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_88_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_88_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_88_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_88_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_88_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_88_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_88_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_88_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_88_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_88_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_88_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_88_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[80]),
    .ccff_tail(grid_clb_88_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__6_
  (
    .clk_0_S_in(clk_1_wires[145]),
    .prog_clk_0_S_in(prog_clk_1_wires[145]),
    .prog_clk_0_E_out(prog_clk_0_wires[307]),
    .prog_clk_0_S_out(prog_clk_0_wires[306]),
    .Test_en_E_out(Test_enWires[148]),
    .Test_en_W_in(Test_enWires[147]),
    .SC_OUT_TOP(scff_Wires[198]),
    .SC_IN_BOT(scff_Wires[197]),
    .top_width_0_height_0__pin_0_(cbx_1__1__82_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__82_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__82_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__82_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__82_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__82_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__82_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__82_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__82_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__82_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__82_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__82_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__82_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__82_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__82_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__82_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[82]),
    .right_width_0_height_0__pin_16_(cby_1__1__89_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__89_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__89_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__89_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__89_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__89_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__89_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__89_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__89_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__89_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__89_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__89_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__89_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__89_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__89_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__89_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__77_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_89_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_89_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_89_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_89_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_89_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_89_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_89_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_89_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_89_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_89_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_89_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_89_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_89_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_89_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_89_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_89_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_89_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_89_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_89_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_89_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_89_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_89_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_89_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_89_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_89_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_89_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_89_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_89_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_89_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_89_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_89_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_89_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[81]),
    .ccff_tail(grid_clb_89_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__7_
  (
    .clk_0_N_in(clk_1_wires[153]),
    .prog_clk_0_N_in(prog_clk_1_wires[153]),
    .prog_clk_0_E_out(prog_clk_0_wires[310]),
    .prog_clk_0_S_out(prog_clk_0_wires[309]),
    .Test_en_E_out(Test_enWires[170]),
    .Test_en_W_in(Test_enWires[169]),
    .SC_OUT_TOP(scff_Wires[200]),
    .SC_IN_BOT(scff_Wires[199]),
    .top_width_0_height_0__pin_0_(cbx_1__1__83_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__83_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__83_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__83_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__83_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__83_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__83_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__83_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__83_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__83_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__83_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__83_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__83_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__83_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__83_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__83_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[83]),
    .right_width_0_height_0__pin_16_(cby_1__1__90_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__90_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__90_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__90_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__90_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__90_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__90_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__90_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__90_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__90_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__90_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__90_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__90_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__90_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__90_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__90_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__78_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_90_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_90_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_90_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_90_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_90_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_90_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_90_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_90_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_90_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_90_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_90_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_90_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_90_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_90_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_90_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_90_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_90_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_90_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_90_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_90_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_90_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_90_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_90_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_90_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_90_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_90_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_90_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_90_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_90_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_90_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_90_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_90_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[82]),
    .ccff_tail(grid_clb_90_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__8_
  (
    .clk_0_S_in(clk_1_wires[152]),
    .prog_clk_0_S_in(prog_clk_1_wires[152]),
    .prog_clk_0_E_out(prog_clk_0_wires[313]),
    .prog_clk_0_S_out(prog_clk_0_wires[312]),
    .Test_en_E_out(Test_enWires[192]),
    .Test_en_W_in(Test_enWires[191]),
    .SC_OUT_TOP(scff_Wires[202]),
    .SC_IN_BOT(scff_Wires[201]),
    .top_width_0_height_0__pin_0_(cbx_1__1__84_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__84_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__84_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__84_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__84_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__84_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__84_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__84_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__84_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__84_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__84_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__84_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__84_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__84_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__84_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__84_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[84]),
    .right_width_0_height_0__pin_16_(cby_1__1__91_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__91_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__91_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__91_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__91_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__91_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__91_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__91_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__91_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__91_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__91_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__91_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__91_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__91_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__91_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__91_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__79_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_91_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_91_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_91_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_91_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_91_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_91_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_91_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_91_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_91_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_91_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_91_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_91_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_91_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_91_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_91_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_91_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_91_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_91_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_91_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_91_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_91_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_91_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_91_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_91_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_91_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_91_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_91_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_91_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_91_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_91_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_91_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_91_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[83]),
    .ccff_tail(grid_clb_91_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__9_
  (
    .clk_0_N_in(clk_1_wires[160]),
    .prog_clk_0_N_in(prog_clk_1_wires[160]),
    .prog_clk_0_E_out(prog_clk_0_wires[316]),
    .prog_clk_0_S_out(prog_clk_0_wires[315]),
    .Test_en_E_out(Test_enWires[214]),
    .Test_en_W_in(Test_enWires[213]),
    .SC_OUT_TOP(scff_Wires[204]),
    .SC_IN_BOT(scff_Wires[203]),
    .top_width_0_height_0__pin_0_(cbx_1__1__85_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__85_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__85_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__85_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__85_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__85_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__85_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__85_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__85_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__85_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__85_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__85_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__85_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__85_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__85_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__85_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[85]),
    .right_width_0_height_0__pin_16_(cby_1__1__92_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__92_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__92_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__92_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__92_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__92_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__92_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__92_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__92_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__92_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__92_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__92_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__92_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__92_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__92_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__92_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__80_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_92_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_92_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_92_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_92_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_92_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_92_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_92_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_92_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_92_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_92_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_92_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_92_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_92_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_92_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_92_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_92_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_92_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_92_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_92_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_92_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_92_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_92_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_92_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_92_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_92_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_92_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_92_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_92_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_92_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_92_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_92_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_92_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[84]),
    .ccff_tail(grid_clb_92_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__10_
  (
    .clk_0_S_in(clk_1_wires[159]),
    .prog_clk_0_S_in(prog_clk_1_wires[159]),
    .prog_clk_0_E_out(prog_clk_0_wires[319]),
    .prog_clk_0_S_out(prog_clk_0_wires[318]),
    .Test_en_E_out(Test_enWires[236]),
    .Test_en_W_in(Test_enWires[235]),
    .SC_OUT_TOP(scff_Wires[206]),
    .SC_IN_BOT(scff_Wires[205]),
    .top_width_0_height_0__pin_0_(cbx_1__1__86_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__86_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__86_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__86_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__86_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__86_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__86_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__86_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__86_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__86_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__86_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__86_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__86_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__86_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__86_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__86_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[86]),
    .right_width_0_height_0__pin_16_(cby_1__1__93_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__93_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__93_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__93_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__93_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__93_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__93_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__93_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__93_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__93_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__93_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__93_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__93_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__93_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__93_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__93_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__81_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_93_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_93_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_93_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_93_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_93_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_93_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_93_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_93_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_93_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_93_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_93_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_93_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_93_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_93_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_93_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_93_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_93_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_93_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_93_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_93_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_93_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_93_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_93_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_93_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_93_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_93_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_93_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_93_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_93_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_93_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_93_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_93_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[85]),
    .ccff_tail(grid_clb_93_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__11_
  (
    .clk_0_N_in(clk_1_wires[167]),
    .prog_clk_0_N_in(prog_clk_1_wires[167]),
    .prog_clk_0_E_out(prog_clk_0_wires[322]),
    .prog_clk_0_S_out(prog_clk_0_wires[321]),
    .Test_en_E_out(Test_enWires[258]),
    .Test_en_W_in(Test_enWires[257]),
    .SC_OUT_TOP(scff_Wires[208]),
    .SC_IN_BOT(scff_Wires[207]),
    .top_width_0_height_0__pin_0_(cbx_1__1__87_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__87_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__87_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__87_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__87_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__87_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__87_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__87_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__87_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__87_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__87_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__87_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__87_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__87_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__87_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__87_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[87]),
    .right_width_0_height_0__pin_16_(cby_1__1__94_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__94_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__94_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__94_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__94_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__94_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__94_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__94_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__94_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__94_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__94_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__94_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__94_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__94_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__94_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__94_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__82_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_94_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_94_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_94_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_94_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_94_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_94_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_94_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_94_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_94_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_94_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_94_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_94_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_94_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_94_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_94_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_94_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_94_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_94_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_94_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_94_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_94_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_94_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_94_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_94_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_94_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_94_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_94_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_94_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_94_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_94_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_94_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_94_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[86]),
    .ccff_tail(grid_clb_94_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__12_
  (
    .clk_0_S_in(clk_1_wires[166]),
    .prog_clk_0_S_in(prog_clk_1_wires[166]),
    .prog_clk_0_N_out(prog_clk_0_wires[327]),
    .prog_clk_0_E_out(prog_clk_0_wires[325]),
    .prog_clk_0_S_out(prog_clk_0_wires[324]),
    .Test_en_E_out(Test_enWires[280]),
    .Test_en_W_in(Test_enWires[279]),
    .SC_OUT_TOP(scff_Wires[210]),
    .SC_IN_BOT(scff_Wires[209]),
    .top_width_0_height_0__pin_0_(cbx_1__12__7_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__7_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__7_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__7_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__7_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__7_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__7_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__7_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__7_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__7_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__7_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__7_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__7_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__7_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__7_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__7_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_8__12__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__95_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__95_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__95_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__95_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__95_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__95_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__95_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__95_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__95_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__95_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__95_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__95_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__95_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__95_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__95_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__95_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__83_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_95_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_95_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_95_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_95_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_95_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_95_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_95_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_95_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_95_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_95_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_95_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_95_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_95_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_95_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_95_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_95_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_95_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_95_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_95_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_95_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_95_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_95_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_95_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_95_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_95_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_95_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_95_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_95_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_95_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_95_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_95_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_95_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[87]),
    .ccff_tail(grid_clb_95_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__1_
  (
    .clk_0_N_in(clk_1_wires[172]),
    .prog_clk_0_N_in(prog_clk_1_wires[172]),
    .prog_clk_0_E_out(prog_clk_0_wires[330]),
    .prog_clk_0_S_out(prog_clk_0_wires[329]),
    .Test_en_E_out(Test_enWires[40]),
    .Test_en_W_in(Test_enWires[39]),
    .SC_OUT_BOT(scff_Wires[237]),
    .SC_IN_TOP(scff_Wires[235]),
    .top_width_0_height_0__pin_0_(cbx_1__1__88_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__88_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__88_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__88_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__88_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__88_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__88_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__88_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__88_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__88_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__88_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__88_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__88_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__88_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__88_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__88_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[88]),
    .right_width_0_height_0__pin_16_(cby_1__1__96_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__96_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__96_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__96_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__96_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__96_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__96_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__96_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__96_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__96_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__96_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__96_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__96_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__96_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__96_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__96_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__84_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_96_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_96_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_96_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_96_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_96_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_96_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_96_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_96_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_96_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_96_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_96_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_96_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_96_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_96_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_96_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_96_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_96_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_96_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_96_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_96_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_96_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_96_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_96_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_96_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_96_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_96_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_96_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_96_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_96_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_96_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_96_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_96_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_9__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_96_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__2_
  (
    .clk_0_S_in(clk_1_wires[171]),
    .prog_clk_0_S_in(prog_clk_1_wires[171]),
    .prog_clk_0_E_out(prog_clk_0_wires[333]),
    .prog_clk_0_S_out(prog_clk_0_wires[332]),
    .Test_en_E_out(Test_enWires[62]),
    .Test_en_W_in(Test_enWires[61]),
    .SC_OUT_BOT(scff_Wires[234]),
    .SC_IN_TOP(scff_Wires[233]),
    .top_width_0_height_0__pin_0_(cbx_1__1__89_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__89_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__89_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__89_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__89_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__89_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__89_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__89_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__89_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__89_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__89_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__89_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__89_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__89_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__89_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__89_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[89]),
    .right_width_0_height_0__pin_16_(cby_1__1__97_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__97_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__97_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__97_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__97_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__97_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__97_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__97_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__97_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__97_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__97_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__97_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__97_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__97_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__97_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__97_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__85_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_97_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_97_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_97_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_97_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_97_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_97_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_97_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_97_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_97_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_97_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_97_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_97_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_97_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_97_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_97_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_97_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_97_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_97_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_97_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_97_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_97_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_97_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_97_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_97_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_97_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_97_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_97_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_97_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_97_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_97_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_97_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_97_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[88]),
    .ccff_tail(grid_clb_97_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__3_
  (
    .clk_0_N_in(clk_1_wires[179]),
    .prog_clk_0_N_in(prog_clk_1_wires[179]),
    .prog_clk_0_E_out(prog_clk_0_wires[336]),
    .prog_clk_0_S_out(prog_clk_0_wires[335]),
    .Test_en_E_out(Test_enWires[84]),
    .Test_en_W_in(Test_enWires[83]),
    .SC_OUT_BOT(scff_Wires[232]),
    .SC_IN_TOP(scff_Wires[231]),
    .top_width_0_height_0__pin_0_(cbx_1__1__90_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__90_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__90_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__90_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__90_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__90_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__90_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__90_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__90_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__90_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__90_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__90_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__90_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__90_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__90_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__90_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[90]),
    .right_width_0_height_0__pin_16_(cby_1__1__98_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__98_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__98_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__98_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__98_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__98_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__98_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__98_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__98_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__98_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__98_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__98_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__98_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__98_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__98_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__98_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__86_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_98_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_98_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_98_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_98_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_98_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_98_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_98_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_98_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_98_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_98_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_98_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_98_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_98_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_98_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_98_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_98_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_98_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_98_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_98_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_98_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_98_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_98_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_98_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_98_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_98_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_98_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_98_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_98_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_98_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_98_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_98_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_98_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[89]),
    .ccff_tail(grid_clb_98_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__4_
  (
    .clk_0_S_in(clk_1_wires[178]),
    .prog_clk_0_S_in(prog_clk_1_wires[178]),
    .prog_clk_0_E_out(prog_clk_0_wires[339]),
    .prog_clk_0_S_out(prog_clk_0_wires[338]),
    .Test_en_E_out(Test_enWires[106]),
    .Test_en_W_in(Test_enWires[105]),
    .SC_OUT_BOT(scff_Wires[230]),
    .SC_IN_TOP(scff_Wires[229]),
    .top_width_0_height_0__pin_0_(cbx_1__1__91_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__91_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__91_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__91_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__91_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__91_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__91_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__91_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__91_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__91_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__91_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__91_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__91_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__91_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__91_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__91_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[91]),
    .right_width_0_height_0__pin_16_(cby_1__1__99_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__99_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__99_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__99_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__99_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__99_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__99_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__99_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__99_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__99_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__99_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__99_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__99_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__99_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__99_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__99_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__87_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_99_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_99_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_99_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_99_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_99_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_99_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_99_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_99_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_99_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_99_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_99_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_99_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_99_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_99_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_99_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_99_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_99_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_99_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_99_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_99_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_99_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_99_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_99_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_99_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_99_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_99_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_99_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_99_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_99_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_99_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_99_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_99_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[90]),
    .ccff_tail(grid_clb_99_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__5_
  (
    .clk_0_N_in(clk_1_wires[186]),
    .prog_clk_0_N_in(prog_clk_1_wires[186]),
    .prog_clk_0_E_out(prog_clk_0_wires[342]),
    .prog_clk_0_S_out(prog_clk_0_wires[341]),
    .Test_en_E_out(Test_enWires[128]),
    .Test_en_W_in(Test_enWires[127]),
    .SC_OUT_BOT(scff_Wires[228]),
    .SC_IN_TOP(scff_Wires[227]),
    .top_width_0_height_0__pin_0_(cbx_1__1__92_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__92_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__92_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__92_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__92_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__92_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__92_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__92_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__92_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__92_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__92_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__92_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__92_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__92_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__92_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__92_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[92]),
    .right_width_0_height_0__pin_16_(cby_1__1__100_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__100_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__100_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__100_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__100_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__100_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__100_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__100_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__100_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__100_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__100_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__100_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__100_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__100_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__100_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__100_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__88_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_100_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_100_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_100_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_100_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_100_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_100_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_100_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_100_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_100_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_100_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_100_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_100_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_100_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_100_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_100_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_100_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_100_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_100_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_100_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_100_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_100_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_100_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_100_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_100_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_100_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_100_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_100_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_100_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_100_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_100_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_100_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_100_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[91]),
    .ccff_tail(grid_clb_100_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__6_
  (
    .clk_0_S_in(clk_1_wires[185]),
    .prog_clk_0_S_in(prog_clk_1_wires[185]),
    .prog_clk_0_E_out(prog_clk_0_wires[345]),
    .prog_clk_0_S_out(prog_clk_0_wires[344]),
    .Test_en_E_out(Test_enWires[150]),
    .Test_en_W_in(Test_enWires[149]),
    .SC_OUT_BOT(scff_Wires[226]),
    .SC_IN_TOP(scff_Wires[225]),
    .top_width_0_height_0__pin_0_(cbx_1__1__93_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__93_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__93_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__93_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__93_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__93_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__93_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__93_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__93_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__93_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__93_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__93_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__93_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__93_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__93_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__93_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[93]),
    .right_width_0_height_0__pin_16_(cby_1__1__101_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__101_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__101_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__101_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__101_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__101_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__101_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__101_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__101_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__101_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__101_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__101_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__101_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__101_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__101_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__101_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__89_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_101_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_101_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_101_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_101_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_101_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_101_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_101_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_101_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_101_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_101_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_101_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_101_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_101_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_101_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_101_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_101_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_101_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_101_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_101_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_101_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_101_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_101_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_101_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_101_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_101_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_101_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_101_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_101_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_101_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_101_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_101_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_101_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[92]),
    .ccff_tail(grid_clb_101_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__7_
  (
    .clk_0_N_in(clk_1_wires[193]),
    .prog_clk_0_N_in(prog_clk_1_wires[193]),
    .prog_clk_0_E_out(prog_clk_0_wires[348]),
    .prog_clk_0_S_out(prog_clk_0_wires[347]),
    .Test_en_E_out(Test_enWires[172]),
    .Test_en_W_in(Test_enWires[171]),
    .SC_OUT_BOT(scff_Wires[224]),
    .SC_IN_TOP(scff_Wires[223]),
    .top_width_0_height_0__pin_0_(cbx_1__1__94_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__94_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__94_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__94_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__94_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__94_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__94_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__94_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__94_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__94_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__94_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__94_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__94_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__94_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__94_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__94_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[94]),
    .right_width_0_height_0__pin_16_(cby_1__1__102_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__102_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__102_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__102_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__102_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__102_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__102_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__102_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__102_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__102_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__102_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__102_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__102_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__102_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__102_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__102_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__90_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_102_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_102_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_102_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_102_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_102_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_102_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_102_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_102_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_102_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_102_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_102_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_102_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_102_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_102_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_102_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_102_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_102_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_102_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_102_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_102_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_102_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_102_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_102_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_102_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_102_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_102_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_102_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_102_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_102_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_102_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_102_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_102_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[93]),
    .ccff_tail(grid_clb_102_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__8_
  (
    .clk_0_S_in(clk_1_wires[192]),
    .prog_clk_0_S_in(prog_clk_1_wires[192]),
    .prog_clk_0_E_out(prog_clk_0_wires[351]),
    .prog_clk_0_S_out(prog_clk_0_wires[350]),
    .Test_en_E_out(Test_enWires[194]),
    .Test_en_W_in(Test_enWires[193]),
    .SC_OUT_BOT(scff_Wires[222]),
    .SC_IN_TOP(scff_Wires[221]),
    .top_width_0_height_0__pin_0_(cbx_1__1__95_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__95_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__95_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__95_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__95_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__95_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__95_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__95_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__95_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__95_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__95_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__95_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__95_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__95_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__95_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__95_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[95]),
    .right_width_0_height_0__pin_16_(cby_1__1__103_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__103_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__103_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__103_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__103_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__103_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__103_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__103_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__103_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__103_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__103_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__103_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__103_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__103_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__103_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__103_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__91_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_103_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_103_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_103_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_103_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_103_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_103_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_103_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_103_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_103_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_103_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_103_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_103_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_103_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_103_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_103_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_103_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_103_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_103_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_103_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_103_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_103_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_103_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_103_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_103_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_103_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_103_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_103_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_103_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_103_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_103_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_103_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_103_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[94]),
    .ccff_tail(grid_clb_103_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__9_
  (
    .clk_0_N_in(clk_1_wires[200]),
    .prog_clk_0_N_in(prog_clk_1_wires[200]),
    .prog_clk_0_E_out(prog_clk_0_wires[354]),
    .prog_clk_0_S_out(prog_clk_0_wires[353]),
    .Test_en_E_out(Test_enWires[216]),
    .Test_en_W_in(Test_enWires[215]),
    .SC_OUT_BOT(scff_Wires[220]),
    .SC_IN_TOP(scff_Wires[219]),
    .top_width_0_height_0__pin_0_(cbx_1__1__96_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__96_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__96_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__96_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__96_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__96_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__96_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__96_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__96_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__96_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__96_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__96_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__96_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__96_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__96_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__96_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[96]),
    .right_width_0_height_0__pin_16_(cby_1__1__104_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__104_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__104_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__104_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__104_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__104_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__104_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__104_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__104_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__104_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__104_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__104_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__104_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__104_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__104_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__104_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__92_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_104_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_104_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_104_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_104_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_104_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_104_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_104_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_104_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_104_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_104_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_104_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_104_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_104_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_104_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_104_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_104_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_104_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_104_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_104_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_104_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_104_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_104_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_104_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_104_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_104_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_104_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_104_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_104_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_104_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_104_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_104_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_104_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[95]),
    .ccff_tail(grid_clb_104_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__10_
  (
    .clk_0_S_in(clk_1_wires[199]),
    .prog_clk_0_S_in(prog_clk_1_wires[199]),
    .prog_clk_0_E_out(prog_clk_0_wires[357]),
    .prog_clk_0_S_out(prog_clk_0_wires[356]),
    .Test_en_E_out(Test_enWires[238]),
    .Test_en_W_in(Test_enWires[237]),
    .SC_OUT_BOT(scff_Wires[218]),
    .SC_IN_TOP(scff_Wires[217]),
    .top_width_0_height_0__pin_0_(cbx_1__1__97_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__97_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__97_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__97_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__97_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__97_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__97_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__97_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__97_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__97_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__97_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__97_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__97_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__97_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__97_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__97_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[97]),
    .right_width_0_height_0__pin_16_(cby_1__1__105_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__105_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__105_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__105_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__105_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__105_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__105_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__105_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__105_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__105_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__105_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__105_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__105_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__105_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__105_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__105_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__93_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_105_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_105_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_105_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_105_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_105_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_105_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_105_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_105_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_105_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_105_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_105_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_105_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_105_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_105_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_105_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_105_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_105_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_105_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_105_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_105_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_105_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_105_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_105_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_105_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_105_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_105_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_105_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_105_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_105_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_105_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_105_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_105_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[96]),
    .ccff_tail(grid_clb_105_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__11_
  (
    .clk_0_N_in(clk_1_wires[207]),
    .prog_clk_0_N_in(prog_clk_1_wires[207]),
    .prog_clk_0_E_out(prog_clk_0_wires[360]),
    .prog_clk_0_S_out(prog_clk_0_wires[359]),
    .Test_en_E_out(Test_enWires[260]),
    .Test_en_W_in(Test_enWires[259]),
    .SC_OUT_BOT(scff_Wires[216]),
    .SC_IN_TOP(scff_Wires[215]),
    .top_width_0_height_0__pin_0_(cbx_1__1__98_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__98_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__98_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__98_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__98_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__98_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__98_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__98_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__98_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__98_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__98_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__98_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__98_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__98_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__98_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__98_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[98]),
    .right_width_0_height_0__pin_16_(cby_1__1__106_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__106_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__106_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__106_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__106_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__106_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__106_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__106_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__106_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__106_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__106_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__106_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__106_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__106_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__106_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__106_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__94_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_106_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_106_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_106_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_106_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_106_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_106_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_106_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_106_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_106_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_106_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_106_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_106_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_106_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_106_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_106_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_106_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_106_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_106_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_106_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_106_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_106_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_106_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_106_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_106_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_106_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_106_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_106_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_106_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_106_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_106_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_106_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_106_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[97]),
    .ccff_tail(grid_clb_106_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__12_
  (
    .clk_0_S_in(clk_1_wires[206]),
    .prog_clk_0_S_in(prog_clk_1_wires[206]),
    .prog_clk_0_N_out(prog_clk_0_wires[365]),
    .prog_clk_0_E_out(prog_clk_0_wires[363]),
    .prog_clk_0_S_out(prog_clk_0_wires[362]),
    .Test_en_E_out(Test_enWires[282]),
    .Test_en_W_in(Test_enWires[281]),
    .SC_OUT_BOT(scff_Wires[214]),
    .SC_IN_TOP(scff_Wires[213]),
    .top_width_0_height_0__pin_0_(cbx_1__12__8_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__8_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__8_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__8_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__8_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__8_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__8_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__8_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__8_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__8_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__8_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__8_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__8_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__8_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__8_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__8_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_9__12__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__107_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__107_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__107_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__107_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__107_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__107_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__107_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__107_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__107_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__107_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__107_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__107_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__107_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__107_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__107_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__107_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__95_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_107_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_107_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_107_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_107_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_107_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_107_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_107_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_107_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_107_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_107_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_107_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_107_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_107_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_107_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_107_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_107_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_107_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_107_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_107_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_107_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_107_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_107_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_107_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_107_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_107_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_107_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_107_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_107_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_107_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_107_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_107_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_107_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[98]),
    .ccff_tail(grid_clb_107_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__1_
  (
    .clk_0_N_in(clk_1_wires[174]),
    .prog_clk_0_N_in(prog_clk_1_wires[174]),
    .prog_clk_0_E_out(prog_clk_0_wires[368]),
    .prog_clk_0_S_out(prog_clk_0_wires[367]),
    .Test_en_E_out(Test_enWires[42]),
    .Test_en_W_in(Test_enWires[41]),
    .SC_OUT_TOP(scff_Wires[241]),
    .SC_IN_BOT(scff_Wires[240]),
    .top_width_0_height_0__pin_0_(cbx_1__1__99_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__99_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__99_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__99_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__99_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__99_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__99_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__99_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__99_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__99_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__99_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__99_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__99_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__99_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__99_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__99_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[99]),
    .right_width_0_height_0__pin_16_(cby_1__1__108_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__108_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__108_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__108_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__108_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__108_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__108_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__108_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__108_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__108_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__108_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__108_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__108_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__108_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__108_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__108_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__96_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_108_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_108_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_108_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_108_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_108_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_108_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_108_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_108_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_108_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_108_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_108_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_108_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_108_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_108_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_108_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_108_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_108_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_108_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_108_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_108_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_108_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_108_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_108_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_108_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_108_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_108_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_108_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_108_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_108_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_108_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_108_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_108_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_10__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_108_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__2_
  (
    .clk_0_S_in(clk_1_wires[173]),
    .prog_clk_0_S_in(prog_clk_1_wires[173]),
    .prog_clk_0_E_out(prog_clk_0_wires[371]),
    .prog_clk_0_S_out(prog_clk_0_wires[370]),
    .Test_en_E_out(Test_enWires[64]),
    .Test_en_W_in(Test_enWires[63]),
    .SC_OUT_TOP(scff_Wires[243]),
    .SC_IN_BOT(scff_Wires[242]),
    .top_width_0_height_0__pin_0_(cbx_1__1__100_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__100_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__100_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__100_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__100_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__100_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__100_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__100_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__100_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__100_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__100_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__100_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__100_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__100_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__100_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__100_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[100]),
    .right_width_0_height_0__pin_16_(cby_1__1__109_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__109_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__109_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__109_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__109_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__109_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__109_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__109_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__109_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__109_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__109_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__109_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__109_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__109_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__109_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__109_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__97_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_109_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_109_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_109_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_109_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_109_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_109_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_109_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_109_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_109_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_109_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_109_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_109_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_109_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_109_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_109_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_109_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_109_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_109_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_109_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_109_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_109_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_109_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_109_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_109_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_109_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_109_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_109_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_109_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_109_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_109_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_109_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_109_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[99]),
    .ccff_tail(grid_clb_109_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__3_
  (
    .clk_0_N_in(clk_1_wires[181]),
    .prog_clk_0_N_in(prog_clk_1_wires[181]),
    .prog_clk_0_E_out(prog_clk_0_wires[374]),
    .prog_clk_0_S_out(prog_clk_0_wires[373]),
    .Test_en_E_out(Test_enWires[86]),
    .Test_en_W_in(Test_enWires[85]),
    .SC_OUT_TOP(scff_Wires[245]),
    .SC_IN_BOT(scff_Wires[244]),
    .top_width_0_height_0__pin_0_(cbx_1__1__101_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__101_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__101_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__101_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__101_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__101_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__101_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__101_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__101_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__101_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__101_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__101_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__101_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__101_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__101_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__101_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[101]),
    .right_width_0_height_0__pin_16_(cby_1__1__110_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__110_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__110_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__110_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__110_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__110_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__110_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__110_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__110_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__110_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__110_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__110_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__110_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__110_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__110_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__110_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__98_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_110_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_110_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_110_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_110_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_110_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_110_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_110_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_110_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_110_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_110_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_110_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_110_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_110_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_110_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_110_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_110_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_110_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_110_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_110_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_110_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_110_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_110_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_110_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_110_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_110_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_110_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_110_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_110_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_110_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_110_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_110_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_110_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[100]),
    .ccff_tail(grid_clb_110_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__4_
  (
    .clk_0_S_in(clk_1_wires[180]),
    .prog_clk_0_S_in(prog_clk_1_wires[180]),
    .prog_clk_0_E_out(prog_clk_0_wires[377]),
    .prog_clk_0_S_out(prog_clk_0_wires[376]),
    .Test_en_E_out(Test_enWires[108]),
    .Test_en_W_in(Test_enWires[107]),
    .SC_OUT_TOP(scff_Wires[247]),
    .SC_IN_BOT(scff_Wires[246]),
    .top_width_0_height_0__pin_0_(cbx_1__1__102_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__102_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__102_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__102_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__102_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__102_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__102_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__102_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__102_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__102_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__102_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__102_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__102_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__102_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__102_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__102_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[102]),
    .right_width_0_height_0__pin_16_(cby_1__1__111_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__111_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__111_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__111_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__111_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__111_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__111_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__111_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__111_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__111_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__111_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__111_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__111_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__111_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__111_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__111_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__99_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_111_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_111_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_111_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_111_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_111_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_111_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_111_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_111_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_111_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_111_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_111_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_111_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_111_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_111_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_111_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_111_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_111_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_111_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_111_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_111_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_111_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_111_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_111_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_111_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_111_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_111_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_111_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_111_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_111_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_111_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_111_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_111_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[101]),
    .ccff_tail(grid_clb_111_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__5_
  (
    .clk_0_N_in(clk_1_wires[188]),
    .prog_clk_0_N_in(prog_clk_1_wires[188]),
    .prog_clk_0_E_out(prog_clk_0_wires[380]),
    .prog_clk_0_S_out(prog_clk_0_wires[379]),
    .Test_en_E_out(Test_enWires[130]),
    .Test_en_W_in(Test_enWires[129]),
    .SC_OUT_TOP(scff_Wires[249]),
    .SC_IN_BOT(scff_Wires[248]),
    .top_width_0_height_0__pin_0_(cbx_1__1__103_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__103_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__103_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__103_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__103_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__103_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__103_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__103_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__103_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__103_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__103_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__103_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__103_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__103_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__103_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__103_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[103]),
    .right_width_0_height_0__pin_16_(cby_1__1__112_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__112_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__112_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__112_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__112_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__112_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__112_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__112_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__112_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__112_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__112_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__112_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__112_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__112_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__112_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__112_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__100_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_112_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_112_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_112_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_112_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_112_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_112_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_112_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_112_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_112_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_112_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_112_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_112_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_112_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_112_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_112_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_112_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_112_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_112_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_112_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_112_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_112_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_112_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_112_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_112_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_112_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_112_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_112_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_112_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_112_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_112_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_112_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_112_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[102]),
    .ccff_tail(grid_clb_112_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__6_
  (
    .clk_0_S_in(clk_1_wires[187]),
    .prog_clk_0_S_in(prog_clk_1_wires[187]),
    .prog_clk_0_E_out(prog_clk_0_wires[383]),
    .prog_clk_0_S_out(prog_clk_0_wires[382]),
    .Test_en_E_out(Test_enWires[152]),
    .Test_en_W_in(Test_enWires[151]),
    .SC_OUT_TOP(scff_Wires[251]),
    .SC_IN_BOT(scff_Wires[250]),
    .top_width_0_height_0__pin_0_(cbx_1__1__104_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__104_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__104_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__104_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__104_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__104_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__104_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__104_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__104_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__104_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__104_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__104_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__104_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__104_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__104_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__104_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[104]),
    .right_width_0_height_0__pin_16_(cby_1__1__113_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__113_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__113_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__113_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__113_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__113_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__113_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__113_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__113_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__113_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__113_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__113_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__113_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__113_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__113_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__113_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__101_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_113_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_113_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_113_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_113_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_113_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_113_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_113_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_113_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_113_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_113_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_113_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_113_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_113_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_113_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_113_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_113_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_113_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_113_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_113_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_113_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_113_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_113_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_113_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_113_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_113_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_113_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_113_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_113_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_113_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_113_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_113_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_113_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[103]),
    .ccff_tail(grid_clb_113_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__7_
  (
    .clk_0_N_in(clk_1_wires[195]),
    .prog_clk_0_N_in(prog_clk_1_wires[195]),
    .prog_clk_0_E_out(prog_clk_0_wires[386]),
    .prog_clk_0_S_out(prog_clk_0_wires[385]),
    .Test_en_E_out(Test_enWires[174]),
    .Test_en_W_in(Test_enWires[173]),
    .SC_OUT_TOP(scff_Wires[253]),
    .SC_IN_BOT(scff_Wires[252]),
    .top_width_0_height_0__pin_0_(cbx_1__1__105_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__105_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__105_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__105_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__105_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__105_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__105_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__105_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__105_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__105_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__105_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__105_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__105_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__105_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__105_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__105_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[105]),
    .right_width_0_height_0__pin_16_(cby_1__1__114_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__114_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__114_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__114_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__114_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__114_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__114_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__114_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__114_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__114_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__114_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__114_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__114_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__114_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__114_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__114_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__102_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_114_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_114_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_114_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_114_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_114_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_114_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_114_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_114_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_114_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_114_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_114_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_114_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_114_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_114_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_114_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_114_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_114_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_114_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_114_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_114_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_114_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_114_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_114_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_114_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_114_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_114_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_114_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_114_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_114_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_114_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_114_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_114_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[104]),
    .ccff_tail(grid_clb_114_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__8_
  (
    .clk_0_S_in(clk_1_wires[194]),
    .prog_clk_0_S_in(prog_clk_1_wires[194]),
    .prog_clk_0_E_out(prog_clk_0_wires[389]),
    .prog_clk_0_S_out(prog_clk_0_wires[388]),
    .Test_en_E_out(Test_enWires[196]),
    .Test_en_W_in(Test_enWires[195]),
    .SC_OUT_TOP(scff_Wires[255]),
    .SC_IN_BOT(scff_Wires[254]),
    .top_width_0_height_0__pin_0_(cbx_1__1__106_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__106_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__106_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__106_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__106_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__106_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__106_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__106_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__106_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__106_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__106_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__106_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__106_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__106_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__106_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__106_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[106]),
    .right_width_0_height_0__pin_16_(cby_1__1__115_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__115_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__115_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__115_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__115_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__115_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__115_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__115_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__115_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__115_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__115_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__115_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__115_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__115_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__115_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__115_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__103_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_115_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_115_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_115_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_115_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_115_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_115_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_115_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_115_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_115_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_115_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_115_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_115_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_115_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_115_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_115_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_115_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_115_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_115_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_115_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_115_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_115_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_115_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_115_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_115_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_115_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_115_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_115_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_115_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_115_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_115_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_115_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_115_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[105]),
    .ccff_tail(grid_clb_115_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__9_
  (
    .clk_0_N_in(clk_1_wires[202]),
    .prog_clk_0_N_in(prog_clk_1_wires[202]),
    .prog_clk_0_E_out(prog_clk_0_wires[392]),
    .prog_clk_0_S_out(prog_clk_0_wires[391]),
    .Test_en_E_out(Test_enWires[218]),
    .Test_en_W_in(Test_enWires[217]),
    .SC_OUT_TOP(scff_Wires[257]),
    .SC_IN_BOT(scff_Wires[256]),
    .top_width_0_height_0__pin_0_(cbx_1__1__107_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__107_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__107_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__107_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__107_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__107_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__107_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__107_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__107_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__107_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__107_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__107_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__107_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__107_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__107_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__107_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[107]),
    .right_width_0_height_0__pin_16_(cby_1__1__116_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__116_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__116_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__116_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__116_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__116_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__116_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__116_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__116_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__116_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__116_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__116_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__116_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__116_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__116_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__116_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__104_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_116_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_116_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_116_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_116_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_116_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_116_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_116_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_116_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_116_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_116_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_116_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_116_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_116_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_116_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_116_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_116_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_116_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_116_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_116_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_116_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_116_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_116_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_116_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_116_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_116_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_116_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_116_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_116_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_116_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_116_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_116_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_116_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[106]),
    .ccff_tail(grid_clb_116_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__10_
  (
    .clk_0_S_in(clk_1_wires[201]),
    .prog_clk_0_S_in(prog_clk_1_wires[201]),
    .prog_clk_0_E_out(prog_clk_0_wires[395]),
    .prog_clk_0_S_out(prog_clk_0_wires[394]),
    .Test_en_E_out(Test_enWires[240]),
    .Test_en_W_in(Test_enWires[239]),
    .SC_OUT_TOP(scff_Wires[259]),
    .SC_IN_BOT(scff_Wires[258]),
    .top_width_0_height_0__pin_0_(cbx_1__1__108_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__108_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__108_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__108_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__108_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__108_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__108_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__108_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__108_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__108_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__108_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__108_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__108_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__108_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__108_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__108_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[108]),
    .right_width_0_height_0__pin_16_(cby_1__1__117_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__117_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__117_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__117_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__117_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__117_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__117_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__117_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__117_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__117_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__117_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__117_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__117_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__117_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__117_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__117_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__105_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_117_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_117_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_117_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_117_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_117_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_117_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_117_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_117_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_117_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_117_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_117_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_117_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_117_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_117_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_117_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_117_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_117_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_117_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_117_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_117_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_117_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_117_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_117_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_117_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_117_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_117_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_117_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_117_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_117_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_117_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_117_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_117_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[107]),
    .ccff_tail(grid_clb_117_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__11_
  (
    .clk_0_N_in(clk_1_wires[209]),
    .prog_clk_0_N_in(prog_clk_1_wires[209]),
    .prog_clk_0_E_out(prog_clk_0_wires[398]),
    .prog_clk_0_S_out(prog_clk_0_wires[397]),
    .Test_en_E_out(Test_enWires[262]),
    .Test_en_W_in(Test_enWires[261]),
    .SC_OUT_TOP(scff_Wires[261]),
    .SC_IN_BOT(scff_Wires[260]),
    .top_width_0_height_0__pin_0_(cbx_1__1__109_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__109_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__109_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__109_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__109_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__109_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__109_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__109_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__109_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__109_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__109_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__109_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__109_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__109_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__109_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__109_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[109]),
    .right_width_0_height_0__pin_16_(cby_1__1__118_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__118_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__118_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__118_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__118_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__118_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__118_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__118_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__118_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__118_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__118_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__118_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__118_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__118_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__118_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__118_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__106_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_118_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_118_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_118_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_118_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_118_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_118_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_118_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_118_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_118_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_118_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_118_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_118_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_118_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_118_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_118_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_118_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_118_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_118_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_118_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_118_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_118_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_118_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_118_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_118_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_118_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_118_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_118_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_118_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_118_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_118_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_118_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_118_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[108]),
    .ccff_tail(grid_clb_118_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__12_
  (
    .clk_0_S_in(clk_1_wires[208]),
    .prog_clk_0_S_in(prog_clk_1_wires[208]),
    .prog_clk_0_N_out(prog_clk_0_wires[403]),
    .prog_clk_0_E_out(prog_clk_0_wires[401]),
    .prog_clk_0_S_out(prog_clk_0_wires[400]),
    .Test_en_E_out(Test_enWires[284]),
    .Test_en_W_in(Test_enWires[283]),
    .SC_OUT_TOP(scff_Wires[263]),
    .SC_IN_BOT(scff_Wires[262]),
    .top_width_0_height_0__pin_0_(cbx_1__12__9_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__9_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__9_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__9_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__9_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__9_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__9_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__9_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__9_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__9_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__9_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__9_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__9_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__9_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__9_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__9_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_10__12__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__119_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__119_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__119_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__119_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__119_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__119_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__119_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__119_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__119_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__119_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__119_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__119_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__119_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__119_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__119_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__119_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__107_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_119_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_119_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_119_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_119_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_119_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_119_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_119_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_119_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_119_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_119_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_119_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_119_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_119_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_119_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_119_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_119_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_119_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_119_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_119_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_119_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_119_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_119_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_119_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_119_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_119_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_119_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_119_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_119_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_119_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_119_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_119_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_119_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[109]),
    .ccff_tail(grid_clb_119_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__1_
  (
    .clk_0_N_in(clk_1_wires[214]),
    .prog_clk_0_N_in(prog_clk_1_wires[214]),
    .prog_clk_0_E_out(prog_clk_0_wires[406]),
    .prog_clk_0_S_out(prog_clk_0_wires[405]),
    .Test_en_E_out(Test_enWires[44]),
    .Test_en_W_in(Test_enWires[43]),
    .SC_OUT_BOT(scff_Wires[290]),
    .SC_IN_TOP(scff_Wires[288]),
    .top_width_0_height_0__pin_0_(cbx_1__1__110_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__110_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__110_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__110_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__110_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__110_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__110_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__110_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__110_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__110_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__110_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__110_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__110_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__110_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__110_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__110_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[110]),
    .right_width_0_height_0__pin_16_(cby_1__1__120_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__120_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__120_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__120_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__120_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__120_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__120_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__120_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__120_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__120_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__120_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__120_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__120_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__120_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__120_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__120_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__108_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_120_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_120_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_120_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_120_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_120_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_120_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_120_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_120_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_120_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_120_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_120_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_120_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_120_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_120_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_120_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_120_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_120_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_120_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_120_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_120_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_120_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_120_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_120_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_120_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_120_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_120_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_120_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_120_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_120_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_120_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_120_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_120_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_11__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_120_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__2_
  (
    .clk_0_S_in(clk_1_wires[213]),
    .prog_clk_0_S_in(prog_clk_1_wires[213]),
    .prog_clk_0_E_out(prog_clk_0_wires[409]),
    .prog_clk_0_S_out(prog_clk_0_wires[408]),
    .Test_en_E_out(Test_enWires[66]),
    .Test_en_W_in(Test_enWires[65]),
    .SC_OUT_BOT(scff_Wires[287]),
    .SC_IN_TOP(scff_Wires[286]),
    .top_width_0_height_0__pin_0_(cbx_1__1__111_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__111_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__111_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__111_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__111_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__111_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__111_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__111_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__111_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__111_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__111_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__111_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__111_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__111_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__111_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__111_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[111]),
    .right_width_0_height_0__pin_16_(cby_1__1__121_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__121_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__121_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__121_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__121_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__121_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__121_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__121_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__121_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__121_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__121_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__121_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__121_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__121_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__121_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__121_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__109_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_121_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_121_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_121_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_121_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_121_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_121_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_121_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_121_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_121_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_121_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_121_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_121_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_121_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_121_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_121_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_121_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_121_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_121_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_121_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_121_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_121_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_121_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_121_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_121_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_121_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_121_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_121_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_121_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_121_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_121_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_121_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_121_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[110]),
    .ccff_tail(grid_clb_121_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__3_
  (
    .clk_0_N_in(clk_1_wires[221]),
    .prog_clk_0_N_in(prog_clk_1_wires[221]),
    .prog_clk_0_E_out(prog_clk_0_wires[412]),
    .prog_clk_0_S_out(prog_clk_0_wires[411]),
    .Test_en_E_out(Test_enWires[88]),
    .Test_en_W_in(Test_enWires[87]),
    .SC_OUT_BOT(scff_Wires[285]),
    .SC_IN_TOP(scff_Wires[284]),
    .top_width_0_height_0__pin_0_(cbx_1__1__112_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__112_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__112_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__112_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__112_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__112_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__112_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__112_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__112_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__112_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__112_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__112_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__112_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__112_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__112_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__112_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[112]),
    .right_width_0_height_0__pin_16_(cby_1__1__122_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__122_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__122_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__122_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__122_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__122_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__122_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__122_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__122_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__122_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__122_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__122_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__122_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__122_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__122_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__122_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__110_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_122_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_122_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_122_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_122_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_122_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_122_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_122_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_122_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_122_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_122_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_122_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_122_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_122_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_122_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_122_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_122_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_122_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_122_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_122_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_122_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_122_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_122_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_122_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_122_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_122_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_122_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_122_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_122_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_122_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_122_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_122_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_122_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[111]),
    .ccff_tail(grid_clb_122_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__4_
  (
    .clk_0_S_in(clk_1_wires[220]),
    .prog_clk_0_S_in(prog_clk_1_wires[220]),
    .prog_clk_0_E_out(prog_clk_0_wires[415]),
    .prog_clk_0_S_out(prog_clk_0_wires[414]),
    .Test_en_E_out(Test_enWires[110]),
    .Test_en_W_in(Test_enWires[109]),
    .SC_OUT_BOT(scff_Wires[283]),
    .SC_IN_TOP(scff_Wires[282]),
    .top_width_0_height_0__pin_0_(cbx_1__1__113_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__113_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__113_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__113_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__113_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__113_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__113_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__113_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__113_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__113_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__113_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__113_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__113_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__113_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__113_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__113_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[113]),
    .right_width_0_height_0__pin_16_(cby_1__1__123_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__123_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__123_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__123_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__123_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__123_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__123_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__123_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__123_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__123_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__123_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__123_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__123_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__123_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__123_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__123_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__111_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_123_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_123_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_123_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_123_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_123_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_123_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_123_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_123_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_123_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_123_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_123_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_123_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_123_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_123_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_123_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_123_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_123_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_123_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_123_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_123_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_123_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_123_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_123_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_123_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_123_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_123_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_123_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_123_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_123_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_123_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_123_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_123_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[112]),
    .ccff_tail(grid_clb_123_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__5_
  (
    .clk_0_N_in(clk_1_wires[228]),
    .prog_clk_0_N_in(prog_clk_1_wires[228]),
    .prog_clk_0_E_out(prog_clk_0_wires[418]),
    .prog_clk_0_S_out(prog_clk_0_wires[417]),
    .Test_en_E_out(Test_enWires[132]),
    .Test_en_W_in(Test_enWires[131]),
    .SC_OUT_BOT(scff_Wires[281]),
    .SC_IN_TOP(scff_Wires[280]),
    .top_width_0_height_0__pin_0_(cbx_1__1__114_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__114_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__114_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__114_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__114_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__114_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__114_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__114_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__114_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__114_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__114_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__114_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__114_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__114_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__114_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__114_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[114]),
    .right_width_0_height_0__pin_16_(cby_1__1__124_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__124_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__124_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__124_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__124_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__124_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__124_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__124_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__124_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__124_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__124_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__124_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__124_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__124_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__124_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__124_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__112_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_124_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_124_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_124_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_124_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_124_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_124_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_124_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_124_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_124_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_124_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_124_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_124_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_124_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_124_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_124_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_124_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_124_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_124_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_124_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_124_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_124_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_124_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_124_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_124_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_124_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_124_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_124_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_124_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_124_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_124_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_124_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_124_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[113]),
    .ccff_tail(grid_clb_124_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__6_
  (
    .clk_0_S_in(clk_1_wires[227]),
    .prog_clk_0_S_in(prog_clk_1_wires[227]),
    .prog_clk_0_E_out(prog_clk_0_wires[421]),
    .prog_clk_0_S_out(prog_clk_0_wires[420]),
    .Test_en_E_out(Test_enWires[154]),
    .Test_en_W_in(Test_enWires[153]),
    .SC_OUT_BOT(scff_Wires[279]),
    .SC_IN_TOP(scff_Wires[278]),
    .top_width_0_height_0__pin_0_(cbx_1__1__115_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__115_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__115_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__115_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__115_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__115_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__115_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__115_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__115_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__115_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__115_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__115_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__115_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__115_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__115_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__115_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[115]),
    .right_width_0_height_0__pin_16_(cby_1__1__125_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__125_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__125_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__125_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__125_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__125_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__125_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__125_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__125_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__125_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__125_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__125_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__125_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__125_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__125_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__125_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__113_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_125_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_125_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_125_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_125_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_125_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_125_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_125_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_125_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_125_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_125_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_125_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_125_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_125_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_125_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_125_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_125_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_125_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_125_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_125_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_125_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_125_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_125_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_125_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_125_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_125_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_125_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_125_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_125_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_125_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_125_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_125_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_125_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[114]),
    .ccff_tail(grid_clb_125_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__7_
  (
    .clk_0_N_in(clk_1_wires[235]),
    .prog_clk_0_N_in(prog_clk_1_wires[235]),
    .prog_clk_0_E_out(prog_clk_0_wires[424]),
    .prog_clk_0_S_out(prog_clk_0_wires[423]),
    .Test_en_E_out(Test_enWires[176]),
    .Test_en_W_in(Test_enWires[175]),
    .SC_OUT_BOT(scff_Wires[277]),
    .SC_IN_TOP(scff_Wires[276]),
    .top_width_0_height_0__pin_0_(cbx_1__1__116_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__116_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__116_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__116_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__116_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__116_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__116_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__116_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__116_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__116_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__116_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__116_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__116_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__116_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__116_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__116_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[116]),
    .right_width_0_height_0__pin_16_(cby_1__1__126_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__126_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__126_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__126_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__126_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__126_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__126_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__126_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__126_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__126_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__126_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__126_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__126_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__126_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__126_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__126_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__114_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_126_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_126_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_126_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_126_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_126_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_126_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_126_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_126_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_126_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_126_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_126_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_126_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_126_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_126_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_126_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_126_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_126_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_126_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_126_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_126_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_126_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_126_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_126_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_126_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_126_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_126_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_126_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_126_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_126_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_126_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_126_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_126_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[115]),
    .ccff_tail(grid_clb_126_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__8_
  (
    .clk_0_S_in(clk_1_wires[234]),
    .prog_clk_0_S_in(prog_clk_1_wires[234]),
    .prog_clk_0_E_out(prog_clk_0_wires[427]),
    .prog_clk_0_S_out(prog_clk_0_wires[426]),
    .Test_en_E_out(Test_enWires[198]),
    .Test_en_W_in(Test_enWires[197]),
    .SC_OUT_BOT(scff_Wires[275]),
    .SC_IN_TOP(scff_Wires[274]),
    .top_width_0_height_0__pin_0_(cbx_1__1__117_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__117_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__117_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__117_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__117_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__117_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__117_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__117_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__117_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__117_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__117_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__117_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__117_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__117_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__117_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__117_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[117]),
    .right_width_0_height_0__pin_16_(cby_1__1__127_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__127_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__127_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__127_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__127_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__127_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__127_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__127_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__127_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__127_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__127_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__127_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__127_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__127_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__127_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__127_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__115_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_127_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_127_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_127_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_127_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_127_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_127_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_127_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_127_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_127_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_127_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_127_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_127_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_127_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_127_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_127_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_127_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_127_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_127_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_127_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_127_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_127_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_127_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_127_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_127_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_127_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_127_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_127_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_127_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_127_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_127_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_127_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_127_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[116]),
    .ccff_tail(grid_clb_127_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__9_
  (
    .clk_0_N_in(clk_1_wires[242]),
    .prog_clk_0_N_in(prog_clk_1_wires[242]),
    .prog_clk_0_E_out(prog_clk_0_wires[430]),
    .prog_clk_0_S_out(prog_clk_0_wires[429]),
    .Test_en_E_out(Test_enWires[220]),
    .Test_en_W_in(Test_enWires[219]),
    .SC_OUT_BOT(scff_Wires[273]),
    .SC_IN_TOP(scff_Wires[272]),
    .top_width_0_height_0__pin_0_(cbx_1__1__118_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__118_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__118_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__118_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__118_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__118_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__118_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__118_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__118_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__118_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__118_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__118_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__118_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__118_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__118_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__118_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[118]),
    .right_width_0_height_0__pin_16_(cby_1__1__128_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__128_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__128_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__128_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__128_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__128_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__128_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__128_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__128_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__128_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__128_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__128_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__128_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__128_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__128_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__128_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__116_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_128_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_128_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_128_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_128_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_128_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_128_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_128_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_128_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_128_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_128_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_128_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_128_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_128_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_128_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_128_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_128_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_128_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_128_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_128_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_128_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_128_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_128_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_128_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_128_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_128_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_128_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_128_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_128_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_128_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_128_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_128_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_128_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[117]),
    .ccff_tail(grid_clb_128_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__10_
  (
    .clk_0_S_in(clk_1_wires[241]),
    .prog_clk_0_S_in(prog_clk_1_wires[241]),
    .prog_clk_0_E_out(prog_clk_0_wires[433]),
    .prog_clk_0_S_out(prog_clk_0_wires[432]),
    .Test_en_E_out(Test_enWires[242]),
    .Test_en_W_in(Test_enWires[241]),
    .SC_OUT_BOT(scff_Wires[271]),
    .SC_IN_TOP(scff_Wires[270]),
    .top_width_0_height_0__pin_0_(cbx_1__1__119_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__119_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__119_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__119_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__119_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__119_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__119_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__119_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__119_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__119_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__119_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__119_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__119_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__119_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__119_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__119_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[119]),
    .right_width_0_height_0__pin_16_(cby_1__1__129_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__129_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__129_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__129_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__129_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__129_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__129_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__129_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__129_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__129_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__129_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__129_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__129_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__129_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__129_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__129_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__117_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_129_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_129_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_129_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_129_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_129_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_129_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_129_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_129_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_129_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_129_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_129_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_129_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_129_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_129_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_129_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_129_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_129_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_129_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_129_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_129_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_129_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_129_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_129_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_129_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_129_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_129_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_129_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_129_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_129_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_129_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_129_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_129_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[118]),
    .ccff_tail(grid_clb_129_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__11_
  (
    .clk_0_N_in(clk_1_wires[249]),
    .prog_clk_0_N_in(prog_clk_1_wires[249]),
    .prog_clk_0_E_out(prog_clk_0_wires[436]),
    .prog_clk_0_S_out(prog_clk_0_wires[435]),
    .Test_en_E_out(Test_enWires[264]),
    .Test_en_W_in(Test_enWires[263]),
    .SC_OUT_BOT(scff_Wires[269]),
    .SC_IN_TOP(scff_Wires[268]),
    .top_width_0_height_0__pin_0_(cbx_1__1__120_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__120_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__120_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__120_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__120_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__120_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__120_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__120_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__120_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__120_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__120_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__120_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__120_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__120_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__120_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__120_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[120]),
    .right_width_0_height_0__pin_16_(cby_1__1__130_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__130_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__130_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__130_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__130_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__130_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__130_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__130_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__130_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__130_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__130_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__130_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__130_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__130_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__130_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__130_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__118_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_130_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_130_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_130_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_130_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_130_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_130_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_130_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_130_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_130_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_130_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_130_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_130_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_130_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_130_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_130_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_130_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_130_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_130_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_130_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_130_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_130_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_130_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_130_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_130_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_130_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_130_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_130_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_130_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_130_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_130_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_130_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_130_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[119]),
    .ccff_tail(grid_clb_130_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__12_
  (
    .clk_0_S_in(clk_1_wires[248]),
    .prog_clk_0_S_in(prog_clk_1_wires[248]),
    .prog_clk_0_N_out(prog_clk_0_wires[441]),
    .prog_clk_0_E_out(prog_clk_0_wires[439]),
    .prog_clk_0_S_out(prog_clk_0_wires[438]),
    .Test_en_E_out(Test_enWires[286]),
    .Test_en_W_in(Test_enWires[285]),
    .SC_OUT_BOT(scff_Wires[267]),
    .SC_IN_TOP(scff_Wires[266]),
    .top_width_0_height_0__pin_0_(cbx_1__12__10_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__10_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__10_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__10_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__10_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__10_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__10_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__10_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__10_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__10_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__10_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__10_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__10_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__10_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__10_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__10_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_11__12__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__131_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__131_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__131_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__131_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__131_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__131_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__131_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__131_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__131_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__131_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__131_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__131_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__131_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__131_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__131_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__131_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__119_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_131_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_131_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_131_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_131_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_131_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_131_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_131_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_131_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_131_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_131_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_131_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_131_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_131_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_131_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_131_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_131_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_131_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_131_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_131_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_131_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_131_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_131_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_131_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_131_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_131_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_131_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_131_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_131_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_131_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_131_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_131_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_131_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[120]),
    .ccff_tail(grid_clb_131_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__1_
  (
    .clk_0_N_in(clk_1_wires[216]),
    .prog_clk_0_N_in(prog_clk_1_wires[216]),
    .prog_clk_0_E_out(prog_clk_0_wires[444]),
    .prog_clk_0_S_out(prog_clk_0_wires[443]),
    .Test_en_W_in(Test_enWires[45]),
    .SC_OUT_TOP(scff_Wires[294]),
    .SC_IN_BOT(scff_Wires[293]),
    .top_width_0_height_0__pin_0_(cbx_1__1__121_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__121_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__121_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__121_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__121_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__121_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__121_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__121_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__121_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__121_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__121_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__121_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__121_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__121_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__121_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__121_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[121]),
    .right_width_0_height_0__pin_16_(cby_12__1__0_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__0_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__0_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__0_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__0_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__0_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__0_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__0_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__0_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__0_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__0_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__0_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__0_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__0_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__0_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__0_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__120_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_132_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_132_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_132_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_132_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_132_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_132_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_132_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_132_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_132_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_132_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_132_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_132_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_132_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_132_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_132_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_132_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_132_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_132_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_132_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_132_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_132_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_132_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_132_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_132_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_132_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_132_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_132_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_132_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_132_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_132_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_132_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_132_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_12__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_132_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__2_
  (
    .clk_0_S_in(clk_1_wires[215]),
    .prog_clk_0_S_in(prog_clk_1_wires[215]),
    .prog_clk_0_E_out(prog_clk_0_wires[447]),
    .prog_clk_0_S_out(prog_clk_0_wires[446]),
    .Test_en_W_in(Test_enWires[67]),
    .SC_OUT_TOP(scff_Wires[296]),
    .SC_IN_BOT(scff_Wires[295]),
    .top_width_0_height_0__pin_0_(cbx_1__1__122_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__122_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__122_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__122_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__122_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__122_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__122_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__122_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__122_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__122_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__122_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__122_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__122_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__122_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__122_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__122_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[122]),
    .right_width_0_height_0__pin_16_(cby_12__1__1_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__1_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__1_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__1_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__1_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__1_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__1_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__1_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__1_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__1_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__1_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__1_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__1_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__1_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__1_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__1_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__121_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_133_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_133_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_133_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_133_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_133_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_133_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_133_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_133_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_133_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_133_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_133_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_133_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_133_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_133_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_133_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_133_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_133_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_133_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_133_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_133_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_133_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_133_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_133_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_133_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_133_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_133_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_133_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_133_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_133_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_133_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_133_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_133_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[121]),
    .ccff_tail(grid_clb_133_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__3_
  (
    .clk_0_N_in(clk_1_wires[223]),
    .prog_clk_0_N_in(prog_clk_1_wires[223]),
    .prog_clk_0_E_out(prog_clk_0_wires[450]),
    .prog_clk_0_S_out(prog_clk_0_wires[449]),
    .Test_en_W_in(Test_enWires[89]),
    .SC_OUT_TOP(scff_Wires[298]),
    .SC_IN_BOT(scff_Wires[297]),
    .top_width_0_height_0__pin_0_(cbx_1__1__123_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__123_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__123_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__123_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__123_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__123_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__123_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__123_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__123_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__123_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__123_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__123_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__123_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__123_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__123_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__123_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[123]),
    .right_width_0_height_0__pin_16_(cby_12__1__2_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__2_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__2_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__2_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__2_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__2_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__2_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__2_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__2_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__2_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__2_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__2_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__2_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__2_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__2_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__2_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__122_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_134_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_134_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_134_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_134_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_134_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_134_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_134_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_134_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_134_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_134_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_134_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_134_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_134_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_134_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_134_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_134_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_134_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_134_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_134_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_134_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_134_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_134_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_134_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_134_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_134_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_134_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_134_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_134_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_134_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_134_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_134_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_134_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[122]),
    .ccff_tail(grid_clb_134_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__4_
  (
    .clk_0_S_in(clk_1_wires[222]),
    .prog_clk_0_S_in(prog_clk_1_wires[222]),
    .prog_clk_0_E_out(prog_clk_0_wires[453]),
    .prog_clk_0_S_out(prog_clk_0_wires[452]),
    .Test_en_W_in(Test_enWires[111]),
    .SC_OUT_TOP(scff_Wires[300]),
    .SC_IN_BOT(scff_Wires[299]),
    .top_width_0_height_0__pin_0_(cbx_1__1__124_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__124_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__124_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__124_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__124_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__124_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__124_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__124_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__124_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__124_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__124_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__124_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__124_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__124_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__124_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__124_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[124]),
    .right_width_0_height_0__pin_16_(cby_12__1__3_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__3_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__3_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__3_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__3_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__3_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__3_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__3_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__3_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__3_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__3_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__3_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__3_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__3_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__3_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__3_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__123_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_135_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_135_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_135_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_135_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_135_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_135_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_135_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_135_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_135_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_135_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_135_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_135_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_135_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_135_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_135_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_135_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_135_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_135_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_135_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_135_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_135_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_135_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_135_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_135_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_135_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_135_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_135_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_135_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_135_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_135_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_135_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_135_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[123]),
    .ccff_tail(grid_clb_135_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__5_
  (
    .clk_0_N_in(clk_1_wires[230]),
    .prog_clk_0_N_in(prog_clk_1_wires[230]),
    .prog_clk_0_E_out(prog_clk_0_wires[456]),
    .prog_clk_0_S_out(prog_clk_0_wires[455]),
    .Test_en_W_in(Test_enWires[133]),
    .SC_OUT_TOP(scff_Wires[302]),
    .SC_IN_BOT(scff_Wires[301]),
    .top_width_0_height_0__pin_0_(cbx_1__1__125_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__125_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__125_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__125_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__125_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__125_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__125_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__125_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__125_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__125_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__125_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__125_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__125_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__125_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__125_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__125_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[125]),
    .right_width_0_height_0__pin_16_(cby_12__1__4_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__4_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__4_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__4_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__4_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__4_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__4_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__4_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__4_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__4_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__4_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__4_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__4_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__4_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__4_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__4_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__124_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_136_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_136_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_136_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_136_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_136_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_136_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_136_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_136_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_136_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_136_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_136_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_136_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_136_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_136_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_136_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_136_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_136_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_136_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_136_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_136_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_136_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_136_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_136_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_136_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_136_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_136_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_136_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_136_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_136_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_136_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_136_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_136_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[124]),
    .ccff_tail(grid_clb_136_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__6_
  (
    .clk_0_S_in(clk_1_wires[229]),
    .prog_clk_0_S_in(prog_clk_1_wires[229]),
    .prog_clk_0_E_out(prog_clk_0_wires[459]),
    .prog_clk_0_S_out(prog_clk_0_wires[458]),
    .Test_en_W_in(Test_enWires[155]),
    .SC_OUT_TOP(scff_Wires[304]),
    .SC_IN_BOT(scff_Wires[303]),
    .top_width_0_height_0__pin_0_(cbx_1__1__126_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__126_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__126_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__126_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__126_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__126_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__126_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__126_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__126_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__126_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__126_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__126_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__126_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__126_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__126_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__126_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[126]),
    .right_width_0_height_0__pin_16_(cby_12__1__5_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__5_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__5_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__5_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__5_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__5_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__5_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__5_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__5_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__5_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__5_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__5_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__5_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__5_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__5_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__5_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__125_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_137_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_137_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_137_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_137_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_137_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_137_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_137_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_137_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_137_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_137_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_137_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_137_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_137_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_137_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_137_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_137_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_137_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_137_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_137_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_137_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_137_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_137_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_137_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_137_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_137_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_137_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_137_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_137_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_137_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_137_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_137_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_137_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[125]),
    .ccff_tail(grid_clb_137_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__7_
  (
    .clk_0_N_in(clk_1_wires[237]),
    .prog_clk_0_N_in(prog_clk_1_wires[237]),
    .prog_clk_0_E_out(prog_clk_0_wires[462]),
    .prog_clk_0_S_out(prog_clk_0_wires[461]),
    .Test_en_W_in(Test_enWires[177]),
    .SC_OUT_TOP(scff_Wires[306]),
    .SC_IN_BOT(scff_Wires[305]),
    .top_width_0_height_0__pin_0_(cbx_1__1__127_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__127_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__127_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__127_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__127_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__127_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__127_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__127_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__127_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__127_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__127_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__127_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__127_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__127_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__127_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__127_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[127]),
    .right_width_0_height_0__pin_16_(cby_12__1__6_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__6_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__6_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__6_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__6_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__6_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__6_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__6_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__6_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__6_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__6_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__6_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__6_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__6_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__6_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__6_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__126_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_138_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_138_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_138_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_138_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_138_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_138_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_138_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_138_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_138_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_138_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_138_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_138_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_138_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_138_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_138_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_138_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_138_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_138_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_138_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_138_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_138_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_138_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_138_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_138_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_138_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_138_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_138_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_138_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_138_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_138_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_138_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_138_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[126]),
    .ccff_tail(grid_clb_138_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__8_
  (
    .clk_0_S_in(clk_1_wires[236]),
    .prog_clk_0_S_in(prog_clk_1_wires[236]),
    .prog_clk_0_E_out(prog_clk_0_wires[465]),
    .prog_clk_0_S_out(prog_clk_0_wires[464]),
    .Test_en_W_in(Test_enWires[199]),
    .SC_OUT_TOP(scff_Wires[308]),
    .SC_IN_BOT(scff_Wires[307]),
    .top_width_0_height_0__pin_0_(cbx_1__1__128_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__128_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__128_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__128_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__128_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__128_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__128_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__128_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__128_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__128_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__128_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__128_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__128_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__128_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__128_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__128_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[128]),
    .right_width_0_height_0__pin_16_(cby_12__1__7_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__7_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__7_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__7_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__7_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__7_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__7_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__7_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__7_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__7_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__7_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__7_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__7_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__7_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__7_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__7_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__127_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_139_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_139_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_139_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_139_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_139_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_139_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_139_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_139_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_139_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_139_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_139_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_139_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_139_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_139_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_139_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_139_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_139_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_139_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_139_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_139_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_139_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_139_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_139_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_139_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_139_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_139_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_139_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_139_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_139_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_139_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_139_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_139_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[127]),
    .ccff_tail(grid_clb_139_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__9_
  (
    .clk_0_N_in(clk_1_wires[244]),
    .prog_clk_0_N_in(prog_clk_1_wires[244]),
    .prog_clk_0_E_out(prog_clk_0_wires[468]),
    .prog_clk_0_S_out(prog_clk_0_wires[467]),
    .Test_en_W_in(Test_enWires[221]),
    .SC_OUT_TOP(scff_Wires[310]),
    .SC_IN_BOT(scff_Wires[309]),
    .top_width_0_height_0__pin_0_(cbx_1__1__129_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__129_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__129_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__129_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__129_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__129_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__129_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__129_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__129_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__129_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__129_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__129_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__129_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__129_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__129_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__129_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[129]),
    .right_width_0_height_0__pin_16_(cby_12__1__8_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__8_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__8_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__8_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__8_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__8_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__8_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__8_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__8_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__8_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__8_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__8_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__8_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__8_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__8_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__8_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__128_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_140_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_140_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_140_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_140_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_140_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_140_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_140_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_140_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_140_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_140_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_140_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_140_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_140_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_140_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_140_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_140_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_140_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_140_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_140_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_140_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_140_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_140_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_140_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_140_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_140_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_140_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_140_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_140_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_140_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_140_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_140_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_140_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[128]),
    .ccff_tail(grid_clb_140_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__10_
  (
    .clk_0_S_in(clk_1_wires[243]),
    .prog_clk_0_S_in(prog_clk_1_wires[243]),
    .prog_clk_0_E_out(prog_clk_0_wires[471]),
    .prog_clk_0_S_out(prog_clk_0_wires[470]),
    .Test_en_W_in(Test_enWires[243]),
    .SC_OUT_TOP(scff_Wires[312]),
    .SC_IN_BOT(scff_Wires[311]),
    .top_width_0_height_0__pin_0_(cbx_1__1__130_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__130_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__130_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__130_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__130_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__130_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__130_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__130_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__130_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__130_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__130_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__130_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__130_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__130_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__130_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__130_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[130]),
    .right_width_0_height_0__pin_16_(cby_12__1__9_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__9_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__9_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__9_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__9_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__9_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__9_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__9_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__9_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__9_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__9_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__9_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__9_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__9_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__9_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__9_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__129_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_141_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_141_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_141_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_141_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_141_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_141_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_141_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_141_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_141_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_141_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_141_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_141_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_141_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_141_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_141_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_141_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_141_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_141_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_141_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_141_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_141_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_141_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_141_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_141_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_141_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_141_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_141_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_141_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_141_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_141_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_141_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_141_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[129]),
    .ccff_tail(grid_clb_141_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__11_
  (
    .clk_0_N_in(clk_1_wires[251]),
    .prog_clk_0_N_in(prog_clk_1_wires[251]),
    .prog_clk_0_E_out(prog_clk_0_wires[474]),
    .prog_clk_0_S_out(prog_clk_0_wires[473]),
    .Test_en_W_in(Test_enWires[265]),
    .SC_OUT_TOP(scff_Wires[314]),
    .SC_IN_BOT(scff_Wires[313]),
    .top_width_0_height_0__pin_0_(cbx_1__1__131_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__131_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__131_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__131_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__131_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__131_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__131_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__131_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__131_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__131_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__131_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__131_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__131_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__131_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__131_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__131_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[131]),
    .right_width_0_height_0__pin_16_(cby_12__1__10_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__10_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__10_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__10_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__10_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__10_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__10_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__10_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__10_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__10_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__10_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__10_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__10_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__10_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__10_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__10_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__130_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_142_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_142_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_142_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_142_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_142_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_142_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_142_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_142_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_142_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_142_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_142_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_142_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_142_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_142_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_142_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_142_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_142_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_142_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_142_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_142_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_142_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_142_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_142_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_142_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_142_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_142_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_142_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_142_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_142_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_142_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_142_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_142_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[130]),
    .ccff_tail(grid_clb_142_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__12_
  (
    .clk_0_S_in(clk_1_wires[250]),
    .prog_clk_0_S_in(prog_clk_1_wires[250]),
    .prog_clk_0_N_out(prog_clk_0_wires[479]),
    .prog_clk_0_E_out(prog_clk_0_wires[477]),
    .prog_clk_0_S_out(prog_clk_0_wires[476]),
    .Test_en_W_in(Test_enWires[287]),
    .SC_OUT_TOP(scff_Wires[316]),
    .SC_IN_BOT(scff_Wires[315]),
    .top_width_0_height_0__pin_0_(cbx_1__12__11_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__11_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__11_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__11_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__11_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__11_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__11_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__11_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__11_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__11_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__11_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__11_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__11_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__11_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__11_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__11_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_12__12__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_12__1__11_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__11_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__11_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__11_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__11_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__11_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__11_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__11_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__11_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__11_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__11_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__11_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__11_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__11_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__11_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__11_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__131_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_143_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_143_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_143_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_143_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_143_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_143_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_143_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_143_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_143_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_143_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_143_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_143_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_143_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_143_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_143_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_143_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_143_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_143_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_143_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_143_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_143_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_143_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_143_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_143_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_143_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_143_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_143_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_143_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_143_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_143_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_143_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_143_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[131]),
    .ccff_tail(grid_clb_143_ccff_tail[0])
  );


  sb_0__0_
  sb_0__0_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[5]),
    .chany_top_in(cby_0__1__0_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_0_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__0__0_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_11_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_11_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_11_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_11_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_11_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_11_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_11_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_11_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_11_top_width_0_height_0__pin_17_upper[0]),
    .ccff_head(grid_io_bottom_11_ccff_tail[0]),
    .chany_top_out(sb_0__0__0_chany_top_out[0:19]),
    .chanx_right_out(sb_0__0__0_chanx_right_out[0:19]),
    .ccff_tail(ccff_tail[0])
  );


  sb_0__1_
  sb_0__1_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[4]),
    .chany_top_in(cby_0__1__1_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_1_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__0_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_0_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_0_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_0_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_0_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_0_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_0_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_0_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_0_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__0_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_0_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__0_ccff_tail[0]),
    .chany_top_out(sb_0__1__0_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__0_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__0_ccff_tail[0])
  );


  sb_0__1_
  sb_0__2_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[10]),
    .chany_top_in(cby_0__1__2_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_2_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__1_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_1_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_1_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_1_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_1_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_1_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_1_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_1_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_1_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__1_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_1_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__1_ccff_tail[0]),
    .chany_top_out(sb_0__1__1_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__1_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__1_ccff_tail[0])
  );


  sb_0__1_
  sb_0__3_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[15]),
    .chany_top_in(cby_0__1__3_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_3_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__2_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_2_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_2_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_2_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_2_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_2_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_2_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_2_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_2_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__2_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_2_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__2_ccff_tail[0]),
    .chany_top_out(sb_0__1__2_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__2_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__2_ccff_tail[0])
  );


  sb_0__1_
  sb_0__4_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[20]),
    .chany_top_in(cby_0__1__4_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_4_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__3_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_3_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_3_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_3_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_3_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_3_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_3_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_3_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_3_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__3_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_3_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__3_ccff_tail[0]),
    .chany_top_out(sb_0__1__3_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__3_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__3_ccff_tail[0])
  );


  sb_0__1_
  sb_0__5_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[25]),
    .chany_top_in(cby_0__1__5_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_5_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__4_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_4_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_4_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_4_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_4_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_4_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_4_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_4_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_4_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__4_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_4_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__4_ccff_tail[0]),
    .chany_top_out(sb_0__1__4_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__4_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__4_ccff_tail[0])
  );


  sb_0__1_
  sb_0__6_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[30]),
    .chany_top_in(cby_0__1__6_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_6_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__5_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_5_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_5_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_5_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_5_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_5_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_5_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_5_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_5_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__5_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_5_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__5_ccff_tail[0]),
    .chany_top_out(sb_0__1__5_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__5_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__5_ccff_tail[0])
  );


  sb_0__1_
  sb_0__7_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[35]),
    .chany_top_in(cby_0__1__7_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_7_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__6_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_6_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_6_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_6_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_6_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_6_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_6_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_6_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_6_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__6_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_6_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__6_ccff_tail[0]),
    .chany_top_out(sb_0__1__6_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__6_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__6_ccff_tail[0])
  );


  sb_0__1_
  sb_0__8_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[40]),
    .chany_top_in(cby_0__1__8_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_8_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__7_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_7_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_7_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_7_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_7_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_7_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_7_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_7_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_7_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__7_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_7_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__7_ccff_tail[0]),
    .chany_top_out(sb_0__1__7_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__7_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__7_ccff_tail[0])
  );


  sb_0__1_
  sb_0__9_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[45]),
    .chany_top_in(cby_0__1__9_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_9_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__8_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_8_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_8_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_8_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_8_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_8_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_8_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_8_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_8_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__8_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_8_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__8_ccff_tail[0]),
    .chany_top_out(sb_0__1__8_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__8_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__8_ccff_tail[0])
  );


  sb_0__1_
  sb_0__10_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[50]),
    .chany_top_in(cby_0__1__10_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_10_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__9_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_9_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_9_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_9_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_9_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_9_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_9_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_9_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_9_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__9_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_9_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__9_ccff_tail[0]),
    .chany_top_out(sb_0__1__9_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__9_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__9_ccff_tail[0])
  );


  sb_0__1_
  sb_0__11_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[55]),
    .chany_top_in(cby_0__1__11_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_11_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__10_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_10_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_10_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_10_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_10_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_10_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_10_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_10_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_10_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__10_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_10_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__10_ccff_tail[0]),
    .chany_top_out(sb_0__1__10_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__10_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__10_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__10_ccff_tail[0])
  );


  sb_0__2_
  sb_0__12_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[62]),
    .SC_OUT_BOT(scff_Wires[0]),
    .SC_IN_TOP(sc_head),
    .chanx_right_in(cbx_1__12__0_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_0_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_11_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_11_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_11_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_11_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_11_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_11_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_11_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_11_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__11_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_11_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(grid_io_top_0_ccff_tail[0]),
    .chanx_right_out(sb_0__12__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__12__0_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__12__0_ccff_tail[0])
  );


  sb_1__0_
  sb_1__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[2]),
    .SC_OUT_TOP(scff_Wires[27]),
    .SC_IN_TOP(scff_Wires[26]),
    .chany_top_in(cby_1__1__0_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_0_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_0_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_0_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_0_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_0_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_0_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_0_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_0_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__1_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_10_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_10_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_10_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_10_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_10_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_10_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_10_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_10_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_10_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__0_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_11_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_11_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_11_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_11_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_11_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_11_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_11_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_11_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_11_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_10_ccff_tail[0]),
    .chany_top_out(sb_1__0__0_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__0_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__0_ccff_tail[0])
  );


  sb_1__0_
  sb_2__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[65]),
    .chany_top_in(cby_1__1__12_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_12_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_12_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_12_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_12_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_12_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_12_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_12_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_12_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__2_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_9_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_9_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_9_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_9_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_9_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_9_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_9_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_9_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_9_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__1_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_10_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_10_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_10_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_10_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_10_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_10_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_10_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_10_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_10_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_9_ccff_tail[0]),
    .chany_top_out(sb_1__0__1_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__1_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__1_ccff_tail[0])
  );


  sb_1__0_
  sb_3__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[103]),
    .SC_OUT_TOP(scff_Wires[80]),
    .SC_IN_TOP(scff_Wires[79]),
    .chany_top_in(cby_1__1__24_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_24_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_24_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_24_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_24_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_24_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_24_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_24_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_24_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__3_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_8_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_8_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_8_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_8_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_8_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_8_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_8_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_8_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_8_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__2_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_9_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_9_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_9_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_9_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_9_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_9_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_9_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_9_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_9_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_8_ccff_tail[0]),
    .chany_top_out(sb_1__0__2_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__2_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__2_ccff_tail[0])
  );


  sb_1__0_
  sb_4__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[141]),
    .chany_top_in(cby_1__1__36_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_36_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_36_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_36_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_36_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_36_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_36_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_36_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_36_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__4_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_7_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_7_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_7_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_7_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_7_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_7_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_7_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_7_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_7_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__3_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_8_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_8_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_8_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_8_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_8_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_8_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_8_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_8_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_8_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_7_ccff_tail[0]),
    .chany_top_out(sb_1__0__3_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__3_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__3_ccff_tail[0])
  );


  sb_1__0_
  sb_5__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[179]),
    .SC_OUT_TOP(scff_Wires[133]),
    .SC_IN_TOP(scff_Wires[132]),
    .chany_top_in(cby_1__1__48_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_48_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_48_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_48_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_48_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_48_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_48_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_48_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_48_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__5_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_6_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_6_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_6_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_6_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_6_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_6_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_6_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_6_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_6_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__4_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_7_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_7_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_7_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_7_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_7_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_7_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_7_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_7_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_7_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_6_ccff_tail[0]),
    .chany_top_out(sb_1__0__4_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__4_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__4_ccff_tail[0])
  );


  sb_1__0_
  sb_6__0_
  (
    .clk_3_N_out(clk_3_wires[90]),
    .clk_3_S_in(clk),
    .prog_clk_3_N_out(prog_clk_3_wires[90]),
    .prog_clk_3_S_in(prog_clk),
    .prog_clk_0_N_in(prog_clk_0_wires[217]),
    .Test_en_N_out(Test_enWires[1]),
    .Test_en_S_in(Test_en),
    .chany_top_in(cby_1__1__60_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_60_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_60_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_60_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_60_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_60_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_60_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_60_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_60_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__6_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_5_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_5_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_5_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_5_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_5_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_5_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_5_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_5_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_5_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__5_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_6_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_6_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_6_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_6_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_6_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_6_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_6_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_6_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_6_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_5_ccff_tail[0]),
    .chany_top_out(sb_1__0__5_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__5_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__5_ccff_tail[0])
  );


  sb_1__0_
  sb_7__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[255]),
    .SC_OUT_TOP(scff_Wires[186]),
    .SC_IN_TOP(scff_Wires[185]),
    .chany_top_in(cby_1__1__72_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_72_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_72_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_72_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_72_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_72_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_72_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_72_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_72_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__7_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_4_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_4_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_4_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_4_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_4_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_4_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_4_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_4_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_4_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__6_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_5_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_5_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_5_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_5_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_5_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_5_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_5_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_5_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_5_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_4_ccff_tail[0]),
    .chany_top_out(sb_1__0__6_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__6_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__6_ccff_tail[0])
  );


  sb_1__0_
  sb_8__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[293]),
    .chany_top_in(cby_1__1__84_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_84_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_84_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_84_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_84_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_84_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_84_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_84_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_84_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__8_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_3_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_3_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_3_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_3_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_3_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_3_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_3_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_3_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_3_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__7_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_4_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_4_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_4_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_4_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_4_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_4_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_4_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_4_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_4_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_3_ccff_tail[0]),
    .chany_top_out(sb_1__0__7_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__7_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__7_ccff_tail[0])
  );


  sb_1__0_
  sb_9__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[331]),
    .SC_OUT_TOP(scff_Wires[239]),
    .SC_IN_TOP(scff_Wires[238]),
    .chany_top_in(cby_1__1__96_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_96_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_96_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_96_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_96_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_96_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_96_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_96_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_96_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__9_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_2_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_2_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_2_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_2_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_2_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_2_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_2_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_2_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_2_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__8_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_3_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_3_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_3_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_3_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_3_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_3_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_3_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_3_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_3_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_2_ccff_tail[0]),
    .chany_top_out(sb_1__0__8_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__8_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__8_ccff_tail[0])
  );


  sb_1__0_
  sb_10__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[369]),
    .chany_top_in(cby_1__1__108_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_108_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_108_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_108_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_108_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_108_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_108_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_108_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_108_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__10_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_1_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_1_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_1_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_1_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_1_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_1_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_1_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_1_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_1_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__9_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_2_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_2_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_2_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_2_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_2_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_2_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_2_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_2_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_2_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_1_ccff_tail[0]),
    .chany_top_out(sb_1__0__9_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__9_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__9_ccff_tail[0])
  );


  sb_1__0_
  sb_11__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[407]),
    .SC_OUT_TOP(scff_Wires[292]),
    .SC_IN_TOP(scff_Wires[291]),
    .chany_top_in(cby_1__1__120_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_120_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_120_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_120_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_120_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_120_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_120_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_120_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_120_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__11_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_0_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_0_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_0_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_0_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_0_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_0_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_0_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_0_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_0_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__10_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_1_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_1_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_1_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_1_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_1_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_1_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_1_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_1_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_1_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_0_ccff_tail[0]),
    .chany_top_out(sb_1__0__10_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__10_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__10_ccff_tail[0])
  );


  sb_1__1_
  sb_1__1_
  (
    .clk_1_N_in(clk_2_wires[4]),
    .clk_1_W_out(clk_1_wires[2]),
    .clk_1_E_out(clk_1_wires[1]),
    .prog_clk_1_N_in(prog_clk_2_wires[4]),
    .prog_clk_1_W_out(prog_clk_1_wires[2]),
    .prog_clk_1_E_out(prog_clk_1_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[8]),
    .chany_top_in(cby_1__1__1_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_1_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_1_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_1_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_1_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_1_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_1_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_1_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_1_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__11_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_12_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_12_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_12_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_12_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_12_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_12_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_12_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_12_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__0_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_0_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_0_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_0_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_0_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_0_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_0_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_0_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_0_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__0_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_0_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_0_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_0_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_0_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_0_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_0_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_0_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_0_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__11_ccff_tail[0]),
    .chany_top_out(sb_1__1__0_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__0_ccff_tail[0])
  );


  sb_1__1_
  sb_1__2_
  (
    .clk_2_S_out(clk_2_wires[3]),
    .clk_2_E_in(clk_2_wires[1]),
    .prog_clk_2_S_out(prog_clk_2_wires[3]),
    .prog_clk_2_E_in(prog_clk_2_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[13]),
    .chany_top_in(cby_1__1__2_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_2_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_2_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_2_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_2_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_2_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_2_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_2_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_2_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__12_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_13_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_13_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_13_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_13_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_13_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_13_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_13_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_13_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__1_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_1_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_1_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_1_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_1_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_1_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_1_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_1_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_1_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__1_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_1_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_1_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_1_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_1_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_1_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_1_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_1_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_1_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__12_ccff_tail[0]),
    .chany_top_out(sb_1__1__1_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__1_ccff_tail[0])
  );


  sb_1__1_
  sb_1__3_
  (
    .clk_1_N_in(clk_2_wires[11]),
    .clk_1_W_out(clk_1_wires[9]),
    .clk_1_E_out(clk_1_wires[8]),
    .prog_clk_1_N_in(prog_clk_2_wires[11]),
    .prog_clk_1_W_out(prog_clk_1_wires[9]),
    .prog_clk_1_E_out(prog_clk_1_wires[8]),
    .prog_clk_0_N_in(prog_clk_0_wires[18]),
    .chany_top_in(cby_1__1__3_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_3_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_3_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_3_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_3_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_3_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_3_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_3_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_3_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__13_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_14_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_14_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_14_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_14_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_14_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_14_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_14_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_14_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__2_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_2_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_2_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_2_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_2_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_2_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_2_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_2_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_2_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__2_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_2_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_2_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_2_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_2_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_2_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_2_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_2_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_2_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__13_ccff_tail[0]),
    .chany_top_out(sb_1__1__2_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__2_ccff_tail[0])
  );


  sb_1__1_
  sb_1__4_
  (
    .clk_2_S_out(clk_2_wires[10]),
    .clk_2_N_out(clk_2_wires[8]),
    .clk_2_E_in(clk_2_wires[6]),
    .prog_clk_2_S_out(prog_clk_2_wires[10]),
    .prog_clk_2_N_out(prog_clk_2_wires[8]),
    .prog_clk_2_E_in(prog_clk_2_wires[6]),
    .prog_clk_0_N_in(prog_clk_0_wires[23]),
    .chany_top_in(cby_1__1__4_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_4_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_4_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_4_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_4_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_4_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_4_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_4_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_4_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__14_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_15_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_15_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_15_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_15_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_15_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_15_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_15_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_15_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__3_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_3_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_3_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_3_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_3_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_3_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_3_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_3_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_3_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__3_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_3_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_3_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_3_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_3_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_3_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_3_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_3_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_3_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__14_ccff_tail[0]),
    .chany_top_out(sb_1__1__3_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__3_ccff_tail[0])
  );


  sb_1__1_
  sb_1__5_
  (
    .clk_1_S_in(clk_2_wires[9]),
    .clk_1_W_out(clk_1_wires[16]),
    .clk_1_E_out(clk_1_wires[15]),
    .prog_clk_1_S_in(prog_clk_2_wires[9]),
    .prog_clk_1_W_out(prog_clk_1_wires[16]),
    .prog_clk_1_E_out(prog_clk_1_wires[15]),
    .prog_clk_0_N_in(prog_clk_0_wires[28]),
    .chany_top_in(cby_1__1__5_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_5_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_5_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_5_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_5_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_5_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_5_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_5_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_5_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__15_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_16_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_16_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_16_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_16_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_16_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_16_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_16_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_16_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__4_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_4_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_4_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_4_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_4_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_4_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_4_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_4_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_4_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__4_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_4_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_4_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_4_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_4_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_4_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_4_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_4_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_4_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__15_ccff_tail[0]),
    .chany_top_out(sb_1__1__4_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__4_ccff_tail[0])
  );


  sb_1__1_
  sb_1__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[33]),
    .chany_top_in(cby_1__1__6_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_6_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_6_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_6_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_6_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_6_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_6_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_6_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_6_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__16_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_17_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_17_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_17_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_17_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_17_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_17_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_17_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_17_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__5_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_5_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_5_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_5_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_5_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_5_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_5_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_5_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_5_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__5_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_5_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_5_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_5_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_5_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_5_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_5_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_5_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_5_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__16_ccff_tail[0]),
    .chany_top_out(sb_1__1__5_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__5_ccff_tail[0])
  );


  sb_1__1_
  sb_1__7_
  (
    .clk_1_N_in(clk_2_wires[18]),
    .clk_1_W_out(clk_1_wires[23]),
    .clk_1_E_out(clk_1_wires[22]),
    .prog_clk_1_N_in(prog_clk_2_wires[18]),
    .prog_clk_1_W_out(prog_clk_1_wires[23]),
    .prog_clk_1_E_out(prog_clk_1_wires[22]),
    .prog_clk_0_N_in(prog_clk_0_wires[38]),
    .chany_top_in(cby_1__1__7_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_7_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_7_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_7_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_7_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_7_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_7_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_7_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_7_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__17_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_18_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_18_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_18_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_18_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_18_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_18_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_18_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_18_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__6_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_6_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_6_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_6_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_6_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_6_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_6_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_6_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_6_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__6_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_6_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_6_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_6_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_6_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_6_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_6_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_6_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_6_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__17_ccff_tail[0]),
    .chany_top_out(sb_1__1__6_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__6_ccff_tail[0])
  );


  sb_1__1_
  sb_1__8_
  (
    .clk_2_S_out(clk_2_wires[17]),
    .clk_2_N_out(clk_2_wires[15]),
    .clk_2_E_in(clk_2_wires[13]),
    .prog_clk_2_S_out(prog_clk_2_wires[17]),
    .prog_clk_2_N_out(prog_clk_2_wires[15]),
    .prog_clk_2_E_in(prog_clk_2_wires[13]),
    .prog_clk_0_N_in(prog_clk_0_wires[43]),
    .chany_top_in(cby_1__1__8_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_8_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_8_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_8_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_8_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_8_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_8_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_8_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_8_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__18_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_19_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_19_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_19_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_19_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_19_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_19_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_19_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_19_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__7_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_7_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_7_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_7_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_7_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_7_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_7_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_7_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_7_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__7_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_7_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_7_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_7_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_7_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_7_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_7_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_7_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_7_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__18_ccff_tail[0]),
    .chany_top_out(sb_1__1__7_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__7_ccff_tail[0])
  );


  sb_1__1_
  sb_1__9_
  (
    .clk_1_S_in(clk_2_wires[16]),
    .clk_1_W_out(clk_1_wires[30]),
    .clk_1_E_out(clk_1_wires[29]),
    .prog_clk_1_S_in(prog_clk_2_wires[16]),
    .prog_clk_1_W_out(prog_clk_1_wires[30]),
    .prog_clk_1_E_out(prog_clk_1_wires[29]),
    .prog_clk_0_N_in(prog_clk_0_wires[48]),
    .chany_top_in(cby_1__1__9_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_9_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_9_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_9_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_9_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_9_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_9_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_9_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_9_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__19_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_20_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_20_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_20_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_20_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_20_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_20_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_20_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_20_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__8_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_8_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_8_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_8_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_8_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_8_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_8_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_8_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_8_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__8_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_8_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_8_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_8_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_8_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_8_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_8_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_8_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_8_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__19_ccff_tail[0]),
    .chany_top_out(sb_1__1__8_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__8_ccff_tail[0])
  );


  sb_1__1_
  sb_1__10_
  (
    .clk_2_N_out(clk_2_wires[22]),
    .clk_2_E_in(clk_2_wires[20]),
    .prog_clk_2_N_out(prog_clk_2_wires[22]),
    .prog_clk_2_E_in(prog_clk_2_wires[20]),
    .prog_clk_0_N_in(prog_clk_0_wires[53]),
    .chany_top_in(cby_1__1__10_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_10_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_10_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_10_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_10_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_10_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_10_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_10_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_10_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__20_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_21_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_21_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_21_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_21_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_21_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_21_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_21_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_21_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__9_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_9_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_9_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_9_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_9_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_9_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_9_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_9_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_9_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__9_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_9_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_9_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_9_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_9_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_9_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_9_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_9_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_9_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__20_ccff_tail[0]),
    .chany_top_out(sb_1__1__9_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__9_ccff_tail[0])
  );


  sb_1__1_
  sb_1__11_
  (
    .clk_1_S_in(clk_2_wires[23]),
    .clk_1_W_out(clk_1_wires[37]),
    .clk_1_E_out(clk_1_wires[36]),
    .prog_clk_1_S_in(prog_clk_2_wires[23]),
    .prog_clk_1_W_out(prog_clk_1_wires[37]),
    .prog_clk_1_E_out(prog_clk_1_wires[36]),
    .prog_clk_0_N_in(prog_clk_0_wires[58]),
    .chany_top_in(cby_1__1__11_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_11_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_11_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_11_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_11_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_11_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_11_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_11_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_11_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__21_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_22_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_22_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_22_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_22_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_22_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_22_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_22_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_22_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__10_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_10_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_10_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_10_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_10_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_10_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_10_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_10_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_10_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__10_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_10_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_10_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_10_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_10_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_10_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_10_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_10_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_10_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__21_ccff_tail[0]),
    .chany_top_out(sb_1__1__10_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__10_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__10_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__10_ccff_tail[0])
  );


  sb_1__1_
  sb_2__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[68]),
    .chany_top_in(cby_1__1__13_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_13_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_13_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_13_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_13_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_13_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_13_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_13_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_13_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__22_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_24_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_24_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_24_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_24_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_24_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_24_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_24_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_24_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__12_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_12_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_12_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_12_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_12_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_12_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_12_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_12_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_12_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__11_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_12_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_12_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_12_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_12_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_12_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_12_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_12_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_12_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__22_ccff_tail[0]),
    .chany_top_out(sb_1__1__11_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__11_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__11_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__11_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__11_ccff_tail[0])
  );


  sb_1__1_
  sb_2__2_
  (
    .clk_2_N_in(clk_3_wires[69]),
    .clk_2_W_out(clk_2_wires[2]),
    .prog_clk_2_N_in(prog_clk_3_wires[69]),
    .prog_clk_2_W_out(prog_clk_2_wires[2]),
    .prog_clk_0_N_in(prog_clk_0_wires[71]),
    .chany_top_in(cby_1__1__14_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_14_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_14_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_14_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_14_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_14_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_14_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_14_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_14_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__23_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_25_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_25_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_25_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_25_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_25_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_25_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_25_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_25_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__13_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_13_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_13_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_13_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_13_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_13_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_13_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_13_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_13_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__12_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_13_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_13_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_13_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_13_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_13_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_13_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_13_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_13_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__23_ccff_tail[0]),
    .chany_top_out(sb_1__1__12_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__12_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__12_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__12_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__12_ccff_tail[0])
  );


  sb_1__1_
  sb_2__3_
  (
    .clk_3_S_out(clk_3_wires[68]),
    .clk_3_N_in(clk_3_wires[65]),
    .prog_clk_3_S_out(prog_clk_3_wires[68]),
    .prog_clk_3_N_in(prog_clk_3_wires[65]),
    .prog_clk_0_N_in(prog_clk_0_wires[74]),
    .chany_top_in(cby_1__1__15_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_15_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_15_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_15_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_15_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_15_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_15_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_15_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_15_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__24_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_26_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_26_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_26_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_26_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_26_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_26_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_26_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_26_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__14_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_14_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_14_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_14_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_14_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_14_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_14_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_14_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_14_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__13_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_14_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_14_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_14_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_14_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_14_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_14_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_14_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_14_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__24_ccff_tail[0]),
    .chany_top_out(sb_1__1__13_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__13_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__13_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__13_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__13_ccff_tail[0])
  );


  sb_1__1_
  sb_2__4_
  (
    .clk_3_S_out(clk_3_wires[64]),
    .clk_2_N_in(clk_3_wires[59]),
    .clk_3_N_in(clk_3_wires[59]),
    .clk_2_W_out(clk_2_wires[7]),
    .prog_clk_3_S_out(prog_clk_3_wires[64]),
    .prog_clk_2_N_in(prog_clk_3_wires[59]),
    .prog_clk_3_N_in(prog_clk_3_wires[59]),
    .prog_clk_2_W_out(prog_clk_2_wires[7]),
    .prog_clk_0_N_in(prog_clk_0_wires[77]),
    .chany_top_in(cby_1__1__16_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_16_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_16_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_16_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_16_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_16_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_16_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_16_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_16_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__25_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_27_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_27_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_27_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_27_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_27_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_27_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_27_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_27_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__15_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_15_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_15_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_15_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_15_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_15_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_15_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_15_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_15_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__14_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_15_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_15_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_15_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_15_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_15_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_15_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_15_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_15_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__25_ccff_tail[0]),
    .chany_top_out(sb_1__1__14_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__14_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__14_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__14_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__14_ccff_tail[0])
  );


  sb_1__1_
  sb_2__5_
  (
    .clk_3_S_out(clk_3_wires[58]),
    .clk_3_N_in(clk_3_wires[55]),
    .prog_clk_3_S_out(prog_clk_3_wires[58]),
    .prog_clk_3_N_in(prog_clk_3_wires[55]),
    .prog_clk_0_N_in(prog_clk_0_wires[80]),
    .chany_top_in(cby_1__1__17_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_17_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_17_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_17_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_17_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_17_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_17_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_17_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_17_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__26_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_28_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_28_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_28_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_28_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_28_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_28_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_28_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_28_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__16_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_16_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_16_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_16_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_16_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_16_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_16_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_16_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_16_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__15_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_16_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_16_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_16_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_16_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_16_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_16_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_16_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_16_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__26_ccff_tail[0]),
    .chany_top_out(sb_1__1__15_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__15_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__15_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__15_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__15_ccff_tail[0])
  );


  sb_1__1_
  sb_2__6_
  (
    .clk_3_S_out(clk_3_wires[54]),
    .clk_3_N_out(clk_3_wires[52]),
    .clk_3_E_in(clk_3_wires[51]),
    .prog_clk_3_S_out(prog_clk_3_wires[54]),
    .prog_clk_3_N_out(prog_clk_3_wires[52]),
    .prog_clk_3_E_in(prog_clk_3_wires[51]),
    .prog_clk_0_N_in(prog_clk_0_wires[83]),
    .chany_top_in(cby_1__1__18_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_18_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_18_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_18_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_18_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_18_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_18_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_18_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_18_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__27_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_29_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_29_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_29_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_29_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_29_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_29_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_29_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_29_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__17_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_17_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_17_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_17_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_17_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_17_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_17_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_17_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_17_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__16_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_17_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_17_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_17_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_17_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_17_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_17_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_17_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_17_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__27_ccff_tail[0]),
    .chany_top_out(sb_1__1__16_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__16_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__16_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__16_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__16_ccff_tail[0])
  );


  sb_1__1_
  sb_2__7_
  (
    .clk_3_N_out(clk_3_wires[56]),
    .clk_3_S_in(clk_3_wires[53]),
    .prog_clk_3_N_out(prog_clk_3_wires[56]),
    .prog_clk_3_S_in(prog_clk_3_wires[53]),
    .prog_clk_0_N_in(prog_clk_0_wires[86]),
    .chany_top_in(cby_1__1__19_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_19_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_19_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_19_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_19_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_19_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_19_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_19_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_19_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__28_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_30_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_30_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_30_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_30_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_30_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_30_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_30_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_30_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__18_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_18_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_18_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_18_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_18_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_18_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_18_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_18_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_18_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__17_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_18_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_18_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_18_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_18_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_18_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_18_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_18_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_18_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__28_ccff_tail[0]),
    .chany_top_out(sb_1__1__17_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__17_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__17_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__17_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__17_ccff_tail[0])
  );


  sb_1__1_
  sb_2__8_
  (
    .clk_3_N_out(clk_3_wires[62]),
    .clk_2_S_in(clk_3_wires[57]),
    .clk_3_S_in(clk_3_wires[57]),
    .clk_2_W_out(clk_2_wires[14]),
    .prog_clk_3_N_out(prog_clk_3_wires[62]),
    .prog_clk_2_S_in(prog_clk_3_wires[57]),
    .prog_clk_3_S_in(prog_clk_3_wires[57]),
    .prog_clk_2_W_out(prog_clk_2_wires[14]),
    .prog_clk_0_N_in(prog_clk_0_wires[89]),
    .chany_top_in(cby_1__1__20_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_20_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_20_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_20_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_20_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_20_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_20_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_20_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_20_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__29_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_31_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_31_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_31_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_31_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_31_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_31_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_31_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_31_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__19_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_19_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_19_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_19_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_19_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_19_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_19_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_19_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_19_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__18_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_19_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_19_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_19_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_19_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_19_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_19_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_19_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_19_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__29_ccff_tail[0]),
    .chany_top_out(sb_1__1__18_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__18_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__18_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__18_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__18_ccff_tail[0])
  );


  sb_1__1_
  sb_2__9_
  (
    .clk_3_N_out(clk_3_wires[66]),
    .clk_3_S_in(clk_3_wires[63]),
    .prog_clk_3_N_out(prog_clk_3_wires[66]),
    .prog_clk_3_S_in(prog_clk_3_wires[63]),
    .prog_clk_0_N_in(prog_clk_0_wires[92]),
    .chany_top_in(cby_1__1__21_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_21_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_21_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_21_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_21_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_21_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_21_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_21_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_21_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__30_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_32_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_32_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_32_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_32_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_32_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_32_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_32_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_32_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__20_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_20_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_20_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_20_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_20_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_20_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_20_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_20_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_20_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__19_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_20_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_20_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_20_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_20_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_20_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_20_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_20_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_20_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__30_ccff_tail[0]),
    .chany_top_out(sb_1__1__19_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__19_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__19_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__19_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__19_ccff_tail[0])
  );


  sb_1__1_
  sb_2__10_
  (
    .clk_2_S_in(clk_3_wires[67]),
    .clk_2_W_out(clk_2_wires[21]),
    .prog_clk_2_S_in(prog_clk_3_wires[67]),
    .prog_clk_2_W_out(prog_clk_2_wires[21]),
    .prog_clk_0_N_in(prog_clk_0_wires[95]),
    .chany_top_in(cby_1__1__22_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_22_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_22_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_22_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_22_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_22_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_22_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_22_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_22_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__31_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_33_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_33_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_33_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_33_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_33_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_33_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_33_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_33_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__21_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_21_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_21_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_21_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_21_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_21_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_21_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_21_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_21_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__20_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_21_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_21_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_21_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_21_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_21_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_21_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_21_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_21_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__31_ccff_tail[0]),
    .chany_top_out(sb_1__1__20_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__20_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__20_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__20_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__20_ccff_tail[0])
  );


  sb_1__1_
  sb_2__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[98]),
    .chany_top_in(cby_1__1__23_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_23_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_23_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_23_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_23_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_23_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_23_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_23_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_23_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__32_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_34_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_34_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_34_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_34_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_34_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_34_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_34_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_34_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__22_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_22_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_22_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_22_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_22_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_22_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_22_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_22_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_22_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__21_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_22_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_22_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_22_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_22_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_22_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_22_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_22_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_22_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__32_ccff_tail[0]),
    .chany_top_out(sb_1__1__21_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__21_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__21_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__21_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__21_ccff_tail[0])
  );


  sb_1__1_
  sb_3__1_
  (
    .clk_1_N_in(clk_2_wires[30]),
    .clk_1_W_out(clk_1_wires[44]),
    .clk_1_E_out(clk_1_wires[43]),
    .prog_clk_1_N_in(prog_clk_2_wires[30]),
    .prog_clk_1_W_out(prog_clk_1_wires[44]),
    .prog_clk_1_E_out(prog_clk_1_wires[43]),
    .prog_clk_0_N_in(prog_clk_0_wires[106]),
    .chany_top_in(cby_1__1__25_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_25_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_25_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_25_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_25_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_25_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_25_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_25_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_25_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__33_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_36_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_36_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_36_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_36_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_36_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_36_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_36_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_36_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__24_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_24_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_24_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_24_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_24_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_24_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_24_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_24_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_24_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__22_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_24_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_24_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_24_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_24_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_24_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_24_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_24_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_24_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__33_ccff_tail[0]),
    .chany_top_out(sb_1__1__22_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__22_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__22_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__22_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__22_ccff_tail[0])
  );


  sb_1__1_
  sb_3__2_
  (
    .clk_2_S_out(clk_2_wires[29]),
    .clk_2_E_in(clk_2_wires[28]),
    .prog_clk_2_S_out(prog_clk_2_wires[29]),
    .prog_clk_2_E_in(prog_clk_2_wires[28]),
    .prog_clk_0_N_in(prog_clk_0_wires[109]),
    .chany_top_in(cby_1__1__26_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_26_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_26_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_26_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_26_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_26_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_26_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_26_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_26_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__34_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_37_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_37_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_37_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_37_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_37_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_37_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_37_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_37_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__25_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_25_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_25_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_25_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_25_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_25_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_25_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_25_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_25_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__23_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_25_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_25_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_25_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_25_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_25_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_25_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_25_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_25_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__34_ccff_tail[0]),
    .chany_top_out(sb_1__1__23_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__23_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__23_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__23_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__23_ccff_tail[0])
  );


  sb_1__1_
  sb_3__3_
  (
    .clk_1_N_in(clk_2_wires[41]),
    .clk_1_W_out(clk_1_wires[51]),
    .clk_1_E_out(clk_1_wires[50]),
    .prog_clk_1_N_in(prog_clk_2_wires[41]),
    .prog_clk_1_W_out(prog_clk_1_wires[51]),
    .prog_clk_1_E_out(prog_clk_1_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[112]),
    .chany_top_in(cby_1__1__27_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_27_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_27_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_27_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_27_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_27_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_27_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_27_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_27_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__35_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_38_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_38_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_38_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_38_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_38_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_38_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_38_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_38_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__26_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_26_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_26_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_26_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_26_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_26_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_26_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_26_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_26_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__24_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_26_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_26_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_26_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_26_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_26_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_26_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_26_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_26_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__35_ccff_tail[0]),
    .chany_top_out(sb_1__1__24_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__24_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__24_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__24_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__24_ccff_tail[0])
  );


  sb_1__1_
  sb_3__4_
  (
    .clk_2_S_out(clk_2_wires[40]),
    .clk_2_N_out(clk_2_wires[38]),
    .clk_2_E_in(clk_2_wires[37]),
    .prog_clk_2_S_out(prog_clk_2_wires[40]),
    .prog_clk_2_N_out(prog_clk_2_wires[38]),
    .prog_clk_2_E_in(prog_clk_2_wires[37]),
    .prog_clk_0_N_in(prog_clk_0_wires[115]),
    .chany_top_in(cby_1__1__28_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_28_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_28_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_28_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_28_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_28_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_28_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_28_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_28_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__36_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_39_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_39_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_39_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_39_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_39_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_39_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_39_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_39_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__27_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_27_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_27_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_27_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_27_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_27_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_27_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_27_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_27_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__25_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_27_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_27_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_27_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_27_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_27_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_27_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_27_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_27_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__36_ccff_tail[0]),
    .chany_top_out(sb_1__1__25_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__25_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__25_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__25_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__25_ccff_tail[0])
  );


  sb_1__1_
  sb_3__5_
  (
    .clk_1_S_in(clk_2_wires[39]),
    .clk_1_W_out(clk_1_wires[58]),
    .clk_1_E_out(clk_1_wires[57]),
    .prog_clk_1_S_in(prog_clk_2_wires[39]),
    .prog_clk_1_W_out(prog_clk_1_wires[58]),
    .prog_clk_1_E_out(prog_clk_1_wires[57]),
    .prog_clk_0_N_in(prog_clk_0_wires[118]),
    .chany_top_in(cby_1__1__29_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_29_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_29_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_29_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_29_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_29_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_29_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_29_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_29_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__37_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_40_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_40_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_40_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_40_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_40_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_40_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_40_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_40_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__28_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_28_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_28_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_28_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_28_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_28_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_28_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_28_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_28_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__26_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_28_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_28_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_28_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_28_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_28_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_28_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_28_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_28_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__37_ccff_tail[0]),
    .chany_top_out(sb_1__1__26_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__26_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__26_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__26_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__26_ccff_tail[0])
  );


  sb_1__1_
  sb_3__6_
  (
    .clk_3_W_out(clk_3_wires[50]),
    .clk_3_E_in(clk_3_wires[47]),
    .prog_clk_3_W_out(prog_clk_3_wires[50]),
    .prog_clk_3_E_in(prog_clk_3_wires[47]),
    .prog_clk_0_N_in(prog_clk_0_wires[121]),
    .chany_top_in(cby_1__1__30_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_30_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_30_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_30_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_30_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_30_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_30_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_30_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_30_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__38_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_41_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_41_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_41_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_41_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_41_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_41_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_41_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_41_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__29_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_29_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_29_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_29_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_29_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_29_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_29_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_29_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_29_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__27_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_29_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_29_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_29_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_29_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_29_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_29_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_29_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_29_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__38_ccff_tail[0]),
    .chany_top_out(sb_1__1__27_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__27_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__27_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__27_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__27_ccff_tail[0])
  );


  sb_1__1_
  sb_3__7_
  (
    .clk_1_N_in(clk_2_wires[54]),
    .clk_1_W_out(clk_1_wires[65]),
    .clk_1_E_out(clk_1_wires[64]),
    .prog_clk_1_N_in(prog_clk_2_wires[54]),
    .prog_clk_1_W_out(prog_clk_1_wires[65]),
    .prog_clk_1_E_out(prog_clk_1_wires[64]),
    .prog_clk_0_N_in(prog_clk_0_wires[124]),
    .chany_top_in(cby_1__1__31_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_31_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_31_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_31_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_31_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_31_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_31_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_31_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_31_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__39_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_42_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_42_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_42_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_42_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_42_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_42_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_42_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_42_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__30_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_30_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_30_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_30_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_30_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_30_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_30_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_30_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_30_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__28_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_30_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_30_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_30_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_30_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_30_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_30_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_30_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_30_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__39_ccff_tail[0]),
    .chany_top_out(sb_1__1__28_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__28_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__28_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__28_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__28_ccff_tail[0])
  );


  sb_1__1_
  sb_3__8_
  (
    .clk_2_S_out(clk_2_wires[53]),
    .clk_2_N_out(clk_2_wires[51]),
    .clk_2_E_in(clk_2_wires[50]),
    .prog_clk_2_S_out(prog_clk_2_wires[53]),
    .prog_clk_2_N_out(prog_clk_2_wires[51]),
    .prog_clk_2_E_in(prog_clk_2_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[127]),
    .chany_top_in(cby_1__1__32_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_32_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_32_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_32_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_32_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_32_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_32_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_32_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_32_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__40_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_43_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_43_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_43_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_43_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_43_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_43_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_43_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_43_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__31_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_31_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_31_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_31_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_31_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_31_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_31_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_31_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_31_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__29_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_31_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_31_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_31_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_31_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_31_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_31_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_31_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_31_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__40_ccff_tail[0]),
    .chany_top_out(sb_1__1__29_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__29_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__29_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__29_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__29_ccff_tail[0])
  );


  sb_1__1_
  sb_3__9_
  (
    .clk_1_S_in(clk_2_wires[52]),
    .clk_1_W_out(clk_1_wires[72]),
    .clk_1_E_out(clk_1_wires[71]),
    .prog_clk_1_S_in(prog_clk_2_wires[52]),
    .prog_clk_1_W_out(prog_clk_1_wires[72]),
    .prog_clk_1_E_out(prog_clk_1_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[130]),
    .chany_top_in(cby_1__1__33_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_33_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_33_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_33_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_33_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_33_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_33_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_33_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_33_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__41_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_44_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_44_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_44_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_44_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_44_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_44_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_44_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_44_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__32_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_32_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_32_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_32_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_32_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_32_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_32_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_32_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_32_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__30_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_32_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_32_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_32_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_32_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_32_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_32_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_32_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_32_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__41_ccff_tail[0]),
    .chany_top_out(sb_1__1__30_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__30_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__30_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__30_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__30_ccff_tail[0])
  );


  sb_1__1_
  sb_3__10_
  (
    .clk_2_N_out(clk_2_wires[64]),
    .clk_2_E_in(clk_2_wires[63]),
    .prog_clk_2_N_out(prog_clk_2_wires[64]),
    .prog_clk_2_E_in(prog_clk_2_wires[63]),
    .prog_clk_0_N_in(prog_clk_0_wires[133]),
    .chany_top_in(cby_1__1__34_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_34_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_34_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_34_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_34_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_34_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_34_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_34_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_34_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__42_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_45_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_45_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_45_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_45_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_45_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_45_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_45_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_45_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__33_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_33_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_33_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_33_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_33_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_33_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_33_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_33_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_33_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__31_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_33_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_33_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_33_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_33_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_33_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_33_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_33_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_33_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__42_ccff_tail[0]),
    .chany_top_out(sb_1__1__31_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__31_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__31_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__31_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__31_ccff_tail[0])
  );


  sb_1__1_
  sb_3__11_
  (
    .clk_1_S_in(clk_2_wires[65]),
    .clk_1_W_out(clk_1_wires[79]),
    .clk_1_E_out(clk_1_wires[78]),
    .prog_clk_1_S_in(prog_clk_2_wires[65]),
    .prog_clk_1_W_out(prog_clk_1_wires[79]),
    .prog_clk_1_E_out(prog_clk_1_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[136]),
    .chany_top_in(cby_1__1__35_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_35_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_35_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_35_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_35_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_35_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_35_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_35_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_35_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__43_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_46_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_46_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_46_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_46_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_46_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_46_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_46_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_46_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__34_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_34_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_34_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_34_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_34_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_34_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_34_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_34_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_34_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__32_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_34_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_34_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_34_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_34_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_34_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_34_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_34_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_34_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__43_ccff_tail[0]),
    .chany_top_out(sb_1__1__32_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__32_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__32_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__32_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__32_ccff_tail[0])
  );


  sb_1__1_
  sb_4__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[144]),
    .chany_top_in(cby_1__1__37_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_37_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_37_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_37_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_37_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_37_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_37_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_37_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_37_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__44_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_48_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_48_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_48_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_48_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_48_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_48_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_48_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_48_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__36_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_36_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_36_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_36_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_36_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_36_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_36_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_36_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_36_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__33_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_36_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_36_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_36_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_36_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_36_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_36_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_36_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_36_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__44_ccff_tail[0]),
    .chany_top_out(sb_1__1__33_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__33_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__33_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__33_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__33_ccff_tail[0])
  );


  sb_1__1_
  sb_4__2_
  (
    .clk_2_N_in(clk_3_wires[25]),
    .clk_2_W_out(clk_2_wires[27]),
    .clk_2_E_out(clk_2_wires[25]),
    .prog_clk_2_N_in(prog_clk_3_wires[25]),
    .prog_clk_2_W_out(prog_clk_2_wires[27]),
    .prog_clk_2_E_out(prog_clk_2_wires[25]),
    .prog_clk_0_N_in(prog_clk_0_wires[147]),
    .chany_top_in(cby_1__1__38_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_38_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_38_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_38_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_38_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_38_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_38_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_38_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_38_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__45_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_49_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_49_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_49_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_49_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_49_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_49_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_49_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_49_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__37_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_37_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_37_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_37_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_37_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_37_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_37_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_37_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_37_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__34_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_37_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_37_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_37_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_37_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_37_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_37_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_37_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_37_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__45_ccff_tail[0]),
    .chany_top_out(sb_1__1__34_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__34_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__34_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__34_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__34_ccff_tail[0])
  );


  sb_1__1_
  sb_4__3_
  (
    .clk_3_S_out(clk_3_wires[24]),
    .clk_3_N_in(clk_3_wires[21]),
    .prog_clk_3_S_out(prog_clk_3_wires[24]),
    .prog_clk_3_N_in(prog_clk_3_wires[21]),
    .prog_clk_0_N_in(prog_clk_0_wires[150]),
    .chany_top_in(cby_1__1__39_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_39_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_39_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_39_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_39_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_39_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_39_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_39_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_39_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__46_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_50_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_50_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_50_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_50_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_50_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_50_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_50_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_50_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__38_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_38_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_38_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_38_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_38_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_38_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_38_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_38_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_38_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__35_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_38_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_38_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_38_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_38_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_38_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_38_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_38_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_38_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__46_ccff_tail[0]),
    .chany_top_out(sb_1__1__35_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__35_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__35_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__35_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__35_ccff_tail[0])
  );


  sb_1__1_
  sb_4__4_
  (
    .clk_3_S_out(clk_3_wires[20]),
    .clk_2_N_in(clk_3_wires[15]),
    .clk_3_N_in(clk_3_wires[15]),
    .clk_2_W_out(clk_2_wires[36]),
    .clk_2_E_out(clk_2_wires[34]),
    .prog_clk_3_S_out(prog_clk_3_wires[20]),
    .prog_clk_2_N_in(prog_clk_3_wires[15]),
    .prog_clk_3_N_in(prog_clk_3_wires[15]),
    .prog_clk_2_W_out(prog_clk_2_wires[36]),
    .prog_clk_2_E_out(prog_clk_2_wires[34]),
    .prog_clk_0_N_in(prog_clk_0_wires[153]),
    .chany_top_in(cby_1__1__40_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_40_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_40_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_40_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_40_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_40_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_40_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_40_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_40_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__47_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_51_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_51_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_51_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_51_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_51_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_51_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_51_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_51_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__39_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_39_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_39_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_39_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_39_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_39_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_39_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_39_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_39_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__36_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_39_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_39_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_39_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_39_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_39_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_39_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_39_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_39_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__47_ccff_tail[0]),
    .chany_top_out(sb_1__1__36_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__36_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__36_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__36_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__36_ccff_tail[0])
  );


  sb_1__1_
  sb_4__5_
  (
    .clk_3_S_out(clk_3_wires[14]),
    .clk_3_N_in(clk_3_wires[11]),
    .prog_clk_3_S_out(prog_clk_3_wires[14]),
    .prog_clk_3_N_in(prog_clk_3_wires[11]),
    .prog_clk_0_N_in(prog_clk_0_wires[156]),
    .chany_top_in(cby_1__1__41_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_41_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_41_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_41_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_41_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_41_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_41_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_41_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_41_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__48_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_52_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_52_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_52_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_52_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_52_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_52_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_52_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_52_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__40_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_40_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_40_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_40_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_40_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_40_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_40_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_40_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_40_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__37_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_40_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_40_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_40_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_40_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_40_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_40_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_40_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_40_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__48_ccff_tail[0]),
    .chany_top_out(sb_1__1__37_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__37_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__37_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__37_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__37_ccff_tail[0])
  );


  sb_1__1_
  sb_4__6_
  (
    .clk_3_W_out(clk_3_wires[46]),
    .clk_3_S_out(clk_3_wires[10]),
    .clk_3_N_out(clk_3_wires[8]),
    .clk_3_E_in(clk_3_wires[7]),
    .prog_clk_3_W_out(prog_clk_3_wires[46]),
    .prog_clk_3_S_out(prog_clk_3_wires[10]),
    .prog_clk_3_N_out(prog_clk_3_wires[8]),
    .prog_clk_3_E_in(prog_clk_3_wires[7]),
    .prog_clk_0_N_in(prog_clk_0_wires[159]),
    .chany_top_in(cby_1__1__42_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_42_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_42_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_42_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_42_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_42_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_42_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_42_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_42_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__49_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_53_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_53_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_53_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_53_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_53_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_53_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_53_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_53_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__41_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_41_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_41_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_41_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_41_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_41_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_41_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_41_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_41_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__38_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_41_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_41_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_41_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_41_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_41_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_41_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_41_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_41_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__49_ccff_tail[0]),
    .chany_top_out(sb_1__1__38_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__38_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__38_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__38_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__38_ccff_tail[0])
  );


  sb_1__1_
  sb_4__7_
  (
    .clk_3_N_out(clk_3_wires[12]),
    .clk_3_S_in(clk_3_wires[9]),
    .prog_clk_3_N_out(prog_clk_3_wires[12]),
    .prog_clk_3_S_in(prog_clk_3_wires[9]),
    .prog_clk_0_N_in(prog_clk_0_wires[162]),
    .chany_top_in(cby_1__1__43_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_43_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_43_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_43_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_43_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_43_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_43_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_43_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_43_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__50_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_54_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_54_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_54_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_54_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_54_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_54_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_54_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_54_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__42_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_42_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_42_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_42_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_42_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_42_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_42_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_42_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_42_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__39_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_42_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_42_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_42_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_42_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_42_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_42_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_42_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_42_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__50_ccff_tail[0]),
    .chany_top_out(sb_1__1__39_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__39_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__39_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__39_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__39_ccff_tail[0])
  );


  sb_1__1_
  sb_4__8_
  (
    .clk_3_N_out(clk_3_wires[18]),
    .clk_2_S_in(clk_3_wires[13]),
    .clk_3_S_in(clk_3_wires[13]),
    .clk_2_W_out(clk_2_wires[49]),
    .clk_2_E_out(clk_2_wires[47]),
    .prog_clk_3_N_out(prog_clk_3_wires[18]),
    .prog_clk_2_S_in(prog_clk_3_wires[13]),
    .prog_clk_3_S_in(prog_clk_3_wires[13]),
    .prog_clk_2_W_out(prog_clk_2_wires[49]),
    .prog_clk_2_E_out(prog_clk_2_wires[47]),
    .prog_clk_0_N_in(prog_clk_0_wires[165]),
    .chany_top_in(cby_1__1__44_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_44_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_44_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_44_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_44_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_44_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_44_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_44_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_44_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__51_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_55_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_55_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_55_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_55_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_55_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_55_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_55_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_55_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__43_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_43_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_43_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_43_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_43_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_43_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_43_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_43_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_43_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__40_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_43_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_43_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_43_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_43_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_43_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_43_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_43_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_43_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__51_ccff_tail[0]),
    .chany_top_out(sb_1__1__40_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__40_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__40_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__40_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__40_ccff_tail[0])
  );


  sb_1__1_
  sb_4__9_
  (
    .clk_3_N_out(clk_3_wires[22]),
    .clk_3_S_in(clk_3_wires[19]),
    .prog_clk_3_N_out(prog_clk_3_wires[22]),
    .prog_clk_3_S_in(prog_clk_3_wires[19]),
    .prog_clk_0_N_in(prog_clk_0_wires[168]),
    .chany_top_in(cby_1__1__45_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_45_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_45_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_45_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_45_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_45_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_45_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_45_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_45_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__52_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_56_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_56_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_56_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_56_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_56_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_56_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_56_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_56_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__44_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_44_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_44_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_44_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_44_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_44_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_44_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_44_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_44_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__41_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_44_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_44_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_44_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_44_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_44_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_44_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_44_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_44_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__52_ccff_tail[0]),
    .chany_top_out(sb_1__1__41_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__41_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__41_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__41_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__41_ccff_tail[0])
  );


  sb_1__1_
  sb_4__10_
  (
    .clk_2_S_in(clk_3_wires[23]),
    .clk_2_W_out(clk_2_wires[62]),
    .clk_2_E_out(clk_2_wires[60]),
    .prog_clk_2_S_in(prog_clk_3_wires[23]),
    .prog_clk_2_W_out(prog_clk_2_wires[62]),
    .prog_clk_2_E_out(prog_clk_2_wires[60]),
    .prog_clk_0_N_in(prog_clk_0_wires[171]),
    .chany_top_in(cby_1__1__46_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_46_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_46_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_46_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_46_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_46_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_46_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_46_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_46_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__53_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_57_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_57_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_57_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_57_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_57_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_57_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_57_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_57_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__45_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_45_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_45_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_45_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_45_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_45_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_45_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_45_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_45_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__42_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_45_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_45_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_45_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_45_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_45_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_45_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_45_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_45_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__53_ccff_tail[0]),
    .chany_top_out(sb_1__1__42_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__42_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__42_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__42_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__42_ccff_tail[0])
  );


  sb_1__1_
  sb_4__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[174]),
    .chany_top_in(cby_1__1__47_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_47_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_47_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_47_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_47_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_47_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_47_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_47_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_47_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__54_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_58_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_58_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_58_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_58_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_58_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_58_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_58_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_58_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__46_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_46_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_46_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_46_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_46_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_46_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_46_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_46_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_46_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__43_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_46_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_46_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_46_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_46_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_46_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_46_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_46_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_46_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__54_ccff_tail[0]),
    .chany_top_out(sb_1__1__43_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__43_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__43_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__43_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__43_ccff_tail[0])
  );


  sb_1__1_
  sb_5__1_
  (
    .clk_1_N_in(clk_2_wires[32]),
    .clk_1_W_out(clk_1_wires[86]),
    .clk_1_E_out(clk_1_wires[85]),
    .prog_clk_1_N_in(prog_clk_2_wires[32]),
    .prog_clk_1_W_out(prog_clk_1_wires[86]),
    .prog_clk_1_E_out(prog_clk_1_wires[85]),
    .prog_clk_0_N_in(prog_clk_0_wires[182]),
    .chany_top_in(cby_1__1__49_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_49_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_49_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_49_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_49_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_49_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_49_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_49_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_49_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__55_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_60_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_60_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_60_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_60_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_60_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_60_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_60_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_60_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__48_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_48_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_48_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_48_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_48_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_48_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_48_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_48_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_48_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__44_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_48_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_48_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_48_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_48_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_48_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_48_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_48_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_48_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__55_ccff_tail[0]),
    .chany_top_out(sb_1__1__44_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__44_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__44_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__44_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__44_ccff_tail[0])
  );


  sb_1__1_
  sb_5__2_
  (
    .clk_2_S_out(clk_2_wires[31]),
    .clk_2_W_in(clk_2_wires[26]),
    .prog_clk_2_S_out(prog_clk_2_wires[31]),
    .prog_clk_2_W_in(prog_clk_2_wires[26]),
    .prog_clk_0_N_in(prog_clk_0_wires[185]),
    .chany_top_in(cby_1__1__50_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_50_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_50_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_50_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_50_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_50_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_50_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_50_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_50_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__56_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_61_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_61_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_61_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_61_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_61_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_61_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_61_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_61_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__49_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_49_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_49_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_49_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_49_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_49_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_49_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_49_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_49_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__45_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_49_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_49_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_49_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_49_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_49_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_49_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_49_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_49_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__56_ccff_tail[0]),
    .chany_top_out(sb_1__1__45_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__45_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__45_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__45_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__45_ccff_tail[0])
  );


  sb_1__1_
  sb_5__3_
  (
    .clk_1_N_in(clk_2_wires[45]),
    .clk_1_W_out(clk_1_wires[93]),
    .clk_1_E_out(clk_1_wires[92]),
    .prog_clk_1_N_in(prog_clk_2_wires[45]),
    .prog_clk_1_W_out(prog_clk_1_wires[93]),
    .prog_clk_1_E_out(prog_clk_1_wires[92]),
    .prog_clk_0_N_in(prog_clk_0_wires[188]),
    .chany_top_in(cby_1__1__51_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_51_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_51_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_51_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_51_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_51_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_51_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_51_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_51_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__57_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_62_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_62_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_62_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_62_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_62_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_62_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_62_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_62_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__50_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_50_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_50_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_50_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_50_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_50_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_50_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_50_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_50_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__46_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_50_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_50_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_50_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_50_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_50_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_50_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_50_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_50_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__57_ccff_tail[0]),
    .chany_top_out(sb_1__1__46_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__46_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__46_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__46_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__46_ccff_tail[0])
  );


  sb_1__1_
  sb_5__4_
  (
    .clk_2_S_out(clk_2_wires[44]),
    .clk_2_N_out(clk_2_wires[42]),
    .clk_2_W_in(clk_2_wires[35]),
    .prog_clk_2_S_out(prog_clk_2_wires[44]),
    .prog_clk_2_N_out(prog_clk_2_wires[42]),
    .prog_clk_2_W_in(prog_clk_2_wires[35]),
    .prog_clk_0_N_in(prog_clk_0_wires[191]),
    .chany_top_in(cby_1__1__52_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_52_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_52_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_52_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_52_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_52_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_52_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_52_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_52_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__58_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_63_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_63_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_63_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_63_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_63_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_63_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_63_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_63_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__51_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_51_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_51_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_51_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_51_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_51_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_51_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_51_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_51_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__47_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_51_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_51_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_51_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_51_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_51_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_51_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_51_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_51_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__58_ccff_tail[0]),
    .chany_top_out(sb_1__1__47_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__47_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__47_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__47_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__47_ccff_tail[0])
  );


  sb_1__1_
  sb_5__5_
  (
    .clk_1_S_in(clk_2_wires[43]),
    .clk_1_W_out(clk_1_wires[100]),
    .clk_1_E_out(clk_1_wires[99]),
    .prog_clk_1_S_in(prog_clk_2_wires[43]),
    .prog_clk_1_W_out(prog_clk_1_wires[100]),
    .prog_clk_1_E_out(prog_clk_1_wires[99]),
    .prog_clk_0_N_in(prog_clk_0_wires[194]),
    .chany_top_in(cby_1__1__53_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_53_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_53_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_53_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_53_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_53_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_53_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_53_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_53_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__59_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_64_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_64_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_64_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_64_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_64_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_64_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_64_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_64_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__52_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_52_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_52_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_52_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_52_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_52_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_52_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_52_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_52_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__48_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_52_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_52_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_52_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_52_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_52_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_52_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_52_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_52_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__59_ccff_tail[0]),
    .chany_top_out(sb_1__1__48_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__48_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__48_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__48_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__48_ccff_tail[0])
  );


  sb_1__1_
  sb_5__6_
  (
    .clk_3_W_out(clk_3_wires[6]),
    .clk_3_E_in(clk_3_wires[3]),
    .prog_clk_3_W_out(prog_clk_3_wires[6]),
    .prog_clk_3_E_in(prog_clk_3_wires[3]),
    .prog_clk_0_N_in(prog_clk_0_wires[197]),
    .chany_top_in(cby_1__1__54_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_54_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_54_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_54_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_54_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_54_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_54_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_54_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_54_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__60_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_65_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_65_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_65_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_65_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_65_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_65_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_65_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_65_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__53_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_53_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_53_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_53_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_53_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_53_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_53_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_53_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_53_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__49_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_53_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_53_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_53_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_53_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_53_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_53_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_53_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_53_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__60_ccff_tail[0]),
    .chany_top_out(sb_1__1__49_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__49_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__49_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__49_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__49_ccff_tail[0])
  );


  sb_1__1_
  sb_5__7_
  (
    .clk_1_N_in(clk_2_wires[58]),
    .clk_1_W_out(clk_1_wires[107]),
    .clk_1_E_out(clk_1_wires[106]),
    .prog_clk_1_N_in(prog_clk_2_wires[58]),
    .prog_clk_1_W_out(prog_clk_1_wires[107]),
    .prog_clk_1_E_out(prog_clk_1_wires[106]),
    .prog_clk_0_N_in(prog_clk_0_wires[200]),
    .chany_top_in(cby_1__1__55_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_55_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_55_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_55_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_55_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_55_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_55_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_55_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_55_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__61_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_66_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_66_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_66_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_66_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_66_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_66_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_66_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_66_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__54_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_54_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_54_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_54_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_54_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_54_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_54_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_54_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_54_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__50_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_54_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_54_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_54_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_54_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_54_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_54_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_54_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_54_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__61_ccff_tail[0]),
    .chany_top_out(sb_1__1__50_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__50_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__50_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__50_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__50_ccff_tail[0])
  );


  sb_1__1_
  sb_5__8_
  (
    .clk_2_S_out(clk_2_wires[57]),
    .clk_2_N_out(clk_2_wires[55]),
    .clk_2_W_in(clk_2_wires[48]),
    .prog_clk_2_S_out(prog_clk_2_wires[57]),
    .prog_clk_2_N_out(prog_clk_2_wires[55]),
    .prog_clk_2_W_in(prog_clk_2_wires[48]),
    .prog_clk_0_N_in(prog_clk_0_wires[203]),
    .chany_top_in(cby_1__1__56_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_56_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_56_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_56_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_56_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_56_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_56_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_56_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_56_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__62_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_67_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_67_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_67_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_67_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_67_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_67_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_67_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_67_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__55_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_55_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_55_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_55_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_55_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_55_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_55_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_55_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_55_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__51_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_55_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_55_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_55_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_55_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_55_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_55_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_55_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_55_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__62_ccff_tail[0]),
    .chany_top_out(sb_1__1__51_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__51_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__51_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__51_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__51_ccff_tail[0])
  );


  sb_1__1_
  sb_5__9_
  (
    .clk_1_S_in(clk_2_wires[56]),
    .clk_1_W_out(clk_1_wires[114]),
    .clk_1_E_out(clk_1_wires[113]),
    .prog_clk_1_S_in(prog_clk_2_wires[56]),
    .prog_clk_1_W_out(prog_clk_1_wires[114]),
    .prog_clk_1_E_out(prog_clk_1_wires[113]),
    .prog_clk_0_N_in(prog_clk_0_wires[206]),
    .chany_top_in(cby_1__1__57_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_57_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_57_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_57_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_57_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_57_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_57_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_57_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_57_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__63_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_68_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_68_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_68_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_68_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_68_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_68_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_68_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_68_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__56_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_56_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_56_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_56_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_56_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_56_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_56_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_56_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_56_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__52_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_56_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_56_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_56_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_56_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_56_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_56_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_56_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_56_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__63_ccff_tail[0]),
    .chany_top_out(sb_1__1__52_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__52_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__52_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__52_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__52_ccff_tail[0])
  );


  sb_1__1_
  sb_5__10_
  (
    .clk_2_N_out(clk_2_wires[66]),
    .clk_2_W_in(clk_2_wires[61]),
    .prog_clk_2_N_out(prog_clk_2_wires[66]),
    .prog_clk_2_W_in(prog_clk_2_wires[61]),
    .prog_clk_0_N_in(prog_clk_0_wires[209]),
    .chany_top_in(cby_1__1__58_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_58_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_58_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_58_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_58_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_58_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_58_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_58_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_58_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__64_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_69_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_69_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_69_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_69_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_69_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_69_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_69_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_69_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__57_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_57_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_57_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_57_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_57_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_57_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_57_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_57_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_57_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__53_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_57_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_57_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_57_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_57_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_57_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_57_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_57_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_57_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__64_ccff_tail[0]),
    .chany_top_out(sb_1__1__53_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__53_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__53_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__53_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__53_ccff_tail[0])
  );


  sb_1__1_
  sb_5__11_
  (
    .clk_1_S_in(clk_2_wires[67]),
    .clk_1_W_out(clk_1_wires[121]),
    .clk_1_E_out(clk_1_wires[120]),
    .prog_clk_1_S_in(prog_clk_2_wires[67]),
    .prog_clk_1_W_out(prog_clk_1_wires[121]),
    .prog_clk_1_E_out(prog_clk_1_wires[120]),
    .prog_clk_0_N_in(prog_clk_0_wires[212]),
    .chany_top_in(cby_1__1__59_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_59_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_59_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_59_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_59_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_59_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_59_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_59_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_59_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__65_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_70_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_70_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_70_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_70_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_70_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_70_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_70_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_70_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__58_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_58_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_58_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_58_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_58_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_58_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_58_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_58_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_58_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__54_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_58_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_58_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_58_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_58_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_58_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_58_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_58_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_58_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__65_ccff_tail[0]),
    .chany_top_out(sb_1__1__54_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__54_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__54_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__54_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__54_ccff_tail[0])
  );


  sb_1__1_
  sb_6__1_
  (
    .clk_3_N_out(clk_3_wires[92]),
    .clk_3_S_in(clk_3_wires[89]),
    .prog_clk_3_N_out(prog_clk_3_wires[92]),
    .prog_clk_3_S_in(prog_clk_3_wires[89]),
    .prog_clk_0_N_in(prog_clk_0_wires[220]),
    .Test_en_N_out(Test_enWires[3]),
    .Test_en_S_in(Test_enWires[2]),
    .chany_top_in(cby_1__1__61_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_61_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_61_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_61_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_61_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_61_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_61_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_61_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_61_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__66_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_72_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_72_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_72_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_72_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_72_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_72_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_72_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_72_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__60_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_60_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_60_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_60_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_60_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_60_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_60_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_60_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_60_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__55_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_60_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_60_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_60_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_60_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_60_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_60_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_60_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_60_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__66_ccff_tail[0]),
    .chany_top_out(sb_1__1__55_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__55_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__55_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__55_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__55_ccff_tail[0])
  );


  sb_1__1_
  sb_6__2_
  (
    .clk_3_N_out(clk_3_wires[94]),
    .clk_3_S_in(clk_3_wires[91]),
    .prog_clk_3_N_out(prog_clk_3_wires[94]),
    .prog_clk_3_S_in(prog_clk_3_wires[91]),
    .prog_clk_0_N_in(prog_clk_0_wires[223]),
    .Test_en_N_out(Test_enWires[5]),
    .Test_en_S_in(Test_enWires[4]),
    .chany_top_in(cby_1__1__62_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_62_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_62_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_62_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_62_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_62_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_62_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_62_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_62_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__67_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_73_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_73_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_73_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_73_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_73_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_73_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_73_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_73_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__61_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_61_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_61_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_61_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_61_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_61_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_61_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_61_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_61_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__56_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_61_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_61_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_61_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_61_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_61_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_61_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_61_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_61_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__67_ccff_tail[0]),
    .chany_top_out(sb_1__1__56_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__56_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__56_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__56_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__56_ccff_tail[0])
  );


  sb_1__1_
  sb_6__3_
  (
    .clk_3_N_out(clk_3_wires[96]),
    .clk_3_S_in(clk_3_wires[93]),
    .prog_clk_3_N_out(prog_clk_3_wires[96]),
    .prog_clk_3_S_in(prog_clk_3_wires[93]),
    .prog_clk_0_N_in(prog_clk_0_wires[226]),
    .Test_en_N_out(Test_enWires[7]),
    .Test_en_S_in(Test_enWires[6]),
    .chany_top_in(cby_1__1__63_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_63_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_63_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_63_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_63_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_63_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_63_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_63_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_63_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__68_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_74_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_74_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_74_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_74_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_74_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_74_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_74_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_74_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__62_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_62_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_62_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_62_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_62_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_62_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_62_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_62_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_62_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__57_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_62_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_62_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_62_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_62_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_62_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_62_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_62_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_62_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__68_ccff_tail[0]),
    .chany_top_out(sb_1__1__57_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__57_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__57_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__57_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__57_ccff_tail[0])
  );


  sb_1__1_
  sb_6__4_
  (
    .clk_3_N_out(clk_3_wires[98]),
    .clk_3_S_in(clk_3_wires[95]),
    .prog_clk_3_N_out(prog_clk_3_wires[98]),
    .prog_clk_3_S_in(prog_clk_3_wires[95]),
    .prog_clk_0_N_in(prog_clk_0_wires[229]),
    .Test_en_N_out(Test_enWires[9]),
    .Test_en_S_in(Test_enWires[8]),
    .chany_top_in(cby_1__1__64_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_64_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_64_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_64_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_64_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_64_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_64_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_64_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_64_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__69_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_75_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_75_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_75_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_75_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_75_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_75_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_75_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_75_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__63_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_63_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_63_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_63_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_63_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_63_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_63_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_63_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_63_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__58_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_63_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_63_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_63_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_63_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_63_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_63_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_63_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_63_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__69_ccff_tail[0]),
    .chany_top_out(sb_1__1__58_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__58_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__58_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__58_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__58_ccff_tail[0])
  );


  sb_1__1_
  sb_6__5_
  (
    .clk_3_N_out(clk_3_wires[100]),
    .clk_3_S_in(clk_3_wires[97]),
    .prog_clk_3_N_out(prog_clk_3_wires[100]),
    .prog_clk_3_S_in(prog_clk_3_wires[97]),
    .prog_clk_0_N_in(prog_clk_0_wires[232]),
    .Test_en_N_out(Test_enWires[11]),
    .Test_en_S_in(Test_enWires[10]),
    .chany_top_in(cby_1__1__65_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_65_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_65_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_65_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_65_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_65_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_65_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_65_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_65_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__70_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_76_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_76_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_76_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_76_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_76_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_76_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_76_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_76_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__64_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_64_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_64_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_64_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_64_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_64_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_64_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_64_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_64_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__59_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_64_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_64_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_64_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_64_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_64_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_64_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_64_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_64_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__70_ccff_tail[0]),
    .chany_top_out(sb_1__1__59_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__59_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__59_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__59_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__59_ccff_tail[0])
  );


  sb_1__1_
  sb_6__6_
  (
    .clk_3_S_in(clk_3_wires[99]),
    .clk_3_W_out(clk_3_wires[2]),
    .clk_3_E_out(clk_3_wires[0]),
    .prog_clk_3_S_in(prog_clk_3_wires[99]),
    .prog_clk_3_W_out(prog_clk_3_wires[2]),
    .prog_clk_3_E_out(prog_clk_3_wires[0]),
    .prog_clk_0_N_in(prog_clk_0_wires[235]),
    .Test_en_N_out(Test_enWires[13]),
    .Test_en_S_in(Test_enWires[12]),
    .chany_top_in(cby_1__1__66_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_66_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_66_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_66_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_66_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_66_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_66_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_66_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_66_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__71_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_77_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_77_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_77_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_77_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_77_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_77_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_77_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_77_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__65_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_65_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_65_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_65_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_65_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_65_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_65_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_65_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_65_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__60_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_65_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_65_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_65_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_65_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_65_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_65_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_65_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_65_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__71_ccff_tail[0]),
    .chany_top_out(sb_1__1__60_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__60_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__60_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__60_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__60_ccff_tail[0])
  );


  sb_1__1_
  sb_6__7_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[238]),
    .Test_en_N_out(Test_enWires[15]),
    .Test_en_S_in(Test_enWires[14]),
    .chany_top_in(cby_1__1__67_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_67_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_67_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_67_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_67_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_67_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_67_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_67_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_67_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__72_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_78_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_78_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_78_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_78_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_78_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_78_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_78_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_78_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__66_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_66_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_66_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_66_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_66_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_66_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_66_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_66_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_66_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__61_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_66_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_66_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_66_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_66_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_66_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_66_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_66_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_66_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__72_ccff_tail[0]),
    .chany_top_out(sb_1__1__61_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__61_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__61_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__61_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__61_ccff_tail[0])
  );


  sb_1__1_
  sb_6__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[241]),
    .Test_en_N_out(Test_enWires[17]),
    .Test_en_S_in(Test_enWires[16]),
    .chany_top_in(cby_1__1__68_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_68_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_68_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_68_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_68_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_68_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_68_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_68_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_68_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__73_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_79_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_79_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_79_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_79_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_79_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_79_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_79_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_79_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__67_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_67_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_67_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_67_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_67_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_67_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_67_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_67_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_67_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__62_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_67_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_67_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_67_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_67_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_67_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_67_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_67_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_67_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__73_ccff_tail[0]),
    .chany_top_out(sb_1__1__62_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__62_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__62_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__62_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__62_ccff_tail[0])
  );


  sb_1__1_
  sb_6__9_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[244]),
    .Test_en_N_out(Test_enWires[19]),
    .Test_en_S_in(Test_enWires[18]),
    .chany_top_in(cby_1__1__69_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_69_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_69_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_69_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_69_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_69_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_69_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_69_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_69_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__74_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_80_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_80_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_80_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_80_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_80_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_80_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_80_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_80_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__68_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_68_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_68_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_68_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_68_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_68_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_68_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_68_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_68_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__63_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_68_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_68_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_68_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_68_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_68_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_68_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_68_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_68_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__74_ccff_tail[0]),
    .chany_top_out(sb_1__1__63_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__63_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__63_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__63_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__63_ccff_tail[0])
  );


  sb_1__1_
  sb_6__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[247]),
    .Test_en_N_out(Test_enWires[21]),
    .Test_en_S_in(Test_enWires[20]),
    .chany_top_in(cby_1__1__70_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_70_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_70_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_70_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_70_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_70_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_70_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_70_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_70_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__75_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_81_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_81_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_81_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_81_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_81_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_81_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_81_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_81_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__69_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_69_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_69_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_69_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_69_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_69_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_69_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_69_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_69_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__64_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_69_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_69_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_69_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_69_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_69_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_69_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_69_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_69_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__75_ccff_tail[0]),
    .chany_top_out(sb_1__1__64_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__64_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__64_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__64_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__64_ccff_tail[0])
  );


  sb_1__1_
  sb_6__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[250]),
    .Test_en_N_out(Test_enWires[23]),
    .Test_en_S_in(Test_enWires[22]),
    .chany_top_in(cby_1__1__71_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_71_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_71_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_71_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_71_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_71_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_71_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_71_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_71_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__76_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_82_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_82_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_82_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_82_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_82_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_82_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_82_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_82_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__70_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_70_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_70_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_70_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_70_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_70_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_70_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_70_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_70_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__65_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_70_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_70_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_70_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_70_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_70_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_70_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_70_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_70_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__76_ccff_tail[0]),
    .chany_top_out(sb_1__1__65_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__65_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__65_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__65_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__65_ccff_tail[0])
  );


  sb_1__1_
  sb_7__1_
  (
    .clk_1_N_in(clk_2_wires[74]),
    .clk_1_W_out(clk_1_wires[128]),
    .clk_1_E_out(clk_1_wires[127]),
    .prog_clk_1_N_in(prog_clk_2_wires[74]),
    .prog_clk_1_W_out(prog_clk_1_wires[128]),
    .prog_clk_1_E_out(prog_clk_1_wires[127]),
    .prog_clk_0_N_in(prog_clk_0_wires[258]),
    .chany_top_in(cby_1__1__73_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_73_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_73_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_73_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_73_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_73_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_73_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_73_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_73_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__77_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_84_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_84_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_84_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_84_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_84_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_84_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_84_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_84_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__72_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_72_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_72_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_72_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_72_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_72_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_72_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_72_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_72_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__66_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_72_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_72_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_72_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_72_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_72_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_72_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_72_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_72_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__77_ccff_tail[0]),
    .chany_top_out(sb_1__1__66_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__66_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__66_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__66_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__66_ccff_tail[0])
  );


  sb_1__1_
  sb_7__2_
  (
    .clk_2_S_out(clk_2_wires[73]),
    .clk_2_E_in(clk_2_wires[72]),
    .prog_clk_2_S_out(prog_clk_2_wires[73]),
    .prog_clk_2_E_in(prog_clk_2_wires[72]),
    .prog_clk_0_N_in(prog_clk_0_wires[261]),
    .chany_top_in(cby_1__1__74_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_74_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_74_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_74_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_74_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_74_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_74_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_74_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_74_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__78_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_85_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_85_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_85_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_85_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_85_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_85_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_85_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_85_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__73_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_73_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_73_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_73_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_73_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_73_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_73_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_73_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_73_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__67_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_73_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_73_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_73_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_73_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_73_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_73_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_73_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_73_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__78_ccff_tail[0]),
    .chany_top_out(sb_1__1__67_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__67_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__67_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__67_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__67_ccff_tail[0])
  );


  sb_1__1_
  sb_7__3_
  (
    .clk_1_N_in(clk_2_wires[85]),
    .clk_1_W_out(clk_1_wires[135]),
    .clk_1_E_out(clk_1_wires[134]),
    .prog_clk_1_N_in(prog_clk_2_wires[85]),
    .prog_clk_1_W_out(prog_clk_1_wires[135]),
    .prog_clk_1_E_out(prog_clk_1_wires[134]),
    .prog_clk_0_N_in(prog_clk_0_wires[264]),
    .chany_top_in(cby_1__1__75_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_75_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_75_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_75_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_75_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_75_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_75_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_75_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_75_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__79_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_86_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_86_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_86_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_86_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_86_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_86_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_86_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_86_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__74_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_74_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_74_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_74_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_74_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_74_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_74_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_74_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_74_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__68_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_74_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_74_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_74_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_74_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_74_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_74_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_74_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_74_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__79_ccff_tail[0]),
    .chany_top_out(sb_1__1__68_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__68_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__68_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__68_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__68_ccff_tail[0])
  );


  sb_1__1_
  sb_7__4_
  (
    .clk_2_S_out(clk_2_wires[84]),
    .clk_2_N_out(clk_2_wires[82]),
    .clk_2_E_in(clk_2_wires[81]),
    .prog_clk_2_S_out(prog_clk_2_wires[84]),
    .prog_clk_2_N_out(prog_clk_2_wires[82]),
    .prog_clk_2_E_in(prog_clk_2_wires[81]),
    .prog_clk_0_N_in(prog_clk_0_wires[267]),
    .chany_top_in(cby_1__1__76_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_76_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_76_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_76_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_76_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_76_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_76_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_76_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_76_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__80_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_87_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_87_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_87_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_87_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_87_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_87_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_87_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_87_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__75_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_75_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_75_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_75_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_75_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_75_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_75_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_75_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_75_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__69_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_75_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_75_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_75_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_75_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_75_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_75_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_75_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_75_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__80_ccff_tail[0]),
    .chany_top_out(sb_1__1__69_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__69_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__69_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__69_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__69_ccff_tail[0])
  );


  sb_1__1_
  sb_7__5_
  (
    .clk_1_S_in(clk_2_wires[83]),
    .clk_1_W_out(clk_1_wires[142]),
    .clk_1_E_out(clk_1_wires[141]),
    .prog_clk_1_S_in(prog_clk_2_wires[83]),
    .prog_clk_1_W_out(prog_clk_1_wires[142]),
    .prog_clk_1_E_out(prog_clk_1_wires[141]),
    .prog_clk_0_N_in(prog_clk_0_wires[270]),
    .chany_top_in(cby_1__1__77_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_77_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_77_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_77_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_77_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_77_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_77_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_77_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_77_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__81_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_88_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_88_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_88_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_88_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_88_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_88_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_88_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_88_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__76_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_76_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_76_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_76_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_76_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_76_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_76_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_76_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_76_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__70_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_76_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_76_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_76_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_76_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_76_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_76_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_76_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_76_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__81_ccff_tail[0]),
    .chany_top_out(sb_1__1__70_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__70_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__70_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__70_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__70_ccff_tail[0])
  );


  sb_1__1_
  sb_7__6_
  (
    .clk_3_E_out(clk_3_wires[4]),
    .clk_3_W_in(clk_3_wires[1]),
    .prog_clk_3_E_out(prog_clk_3_wires[4]),
    .prog_clk_3_W_in(prog_clk_3_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[273]),
    .chany_top_in(cby_1__1__78_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_78_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_78_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_78_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_78_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_78_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_78_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_78_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_78_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__82_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_89_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_89_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_89_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_89_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_89_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_89_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_89_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_89_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__77_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_77_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_77_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_77_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_77_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_77_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_77_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_77_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_77_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__71_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_77_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_77_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_77_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_77_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_77_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_77_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_77_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_77_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__82_ccff_tail[0]),
    .chany_top_out(sb_1__1__71_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__71_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__71_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__71_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__71_ccff_tail[0])
  );


  sb_1__1_
  sb_7__7_
  (
    .clk_1_N_in(clk_2_wires[98]),
    .clk_1_W_out(clk_1_wires[149]),
    .clk_1_E_out(clk_1_wires[148]),
    .prog_clk_1_N_in(prog_clk_2_wires[98]),
    .prog_clk_1_W_out(prog_clk_1_wires[149]),
    .prog_clk_1_E_out(prog_clk_1_wires[148]),
    .prog_clk_0_N_in(prog_clk_0_wires[276]),
    .chany_top_in(cby_1__1__79_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_79_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_79_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_79_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_79_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_79_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_79_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_79_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_79_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__83_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_90_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_90_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_90_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_90_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_90_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_90_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_90_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_90_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__78_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_78_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_78_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_78_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_78_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_78_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_78_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_78_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_78_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__72_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_78_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_78_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_78_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_78_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_78_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_78_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_78_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_78_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__83_ccff_tail[0]),
    .chany_top_out(sb_1__1__72_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__72_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__72_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__72_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__72_ccff_tail[0])
  );


  sb_1__1_
  sb_7__8_
  (
    .clk_2_S_out(clk_2_wires[97]),
    .clk_2_N_out(clk_2_wires[95]),
    .clk_2_E_in(clk_2_wires[94]),
    .prog_clk_2_S_out(prog_clk_2_wires[97]),
    .prog_clk_2_N_out(prog_clk_2_wires[95]),
    .prog_clk_2_E_in(prog_clk_2_wires[94]),
    .prog_clk_0_N_in(prog_clk_0_wires[279]),
    .chany_top_in(cby_1__1__80_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_80_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_80_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_80_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_80_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_80_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_80_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_80_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_80_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__84_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_91_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_91_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_91_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_91_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_91_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_91_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_91_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_91_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__79_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_79_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_79_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_79_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_79_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_79_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_79_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_79_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_79_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__73_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_79_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_79_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_79_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_79_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_79_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_79_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_79_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_79_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__84_ccff_tail[0]),
    .chany_top_out(sb_1__1__73_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__73_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__73_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__73_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__73_ccff_tail[0])
  );


  sb_1__1_
  sb_7__9_
  (
    .clk_1_S_in(clk_2_wires[96]),
    .clk_1_W_out(clk_1_wires[156]),
    .clk_1_E_out(clk_1_wires[155]),
    .prog_clk_1_S_in(prog_clk_2_wires[96]),
    .prog_clk_1_W_out(prog_clk_1_wires[156]),
    .prog_clk_1_E_out(prog_clk_1_wires[155]),
    .prog_clk_0_N_in(prog_clk_0_wires[282]),
    .chany_top_in(cby_1__1__81_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_81_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_81_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_81_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_81_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_81_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_81_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_81_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_81_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__85_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_92_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_92_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_92_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_92_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_92_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_92_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_92_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_92_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__80_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_80_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_80_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_80_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_80_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_80_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_80_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_80_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_80_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__74_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_80_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_80_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_80_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_80_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_80_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_80_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_80_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_80_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__85_ccff_tail[0]),
    .chany_top_out(sb_1__1__74_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__74_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__74_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__74_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__74_ccff_tail[0])
  );


  sb_1__1_
  sb_7__10_
  (
    .clk_2_N_out(clk_2_wires[108]),
    .clk_2_E_in(clk_2_wires[107]),
    .prog_clk_2_N_out(prog_clk_2_wires[108]),
    .prog_clk_2_E_in(prog_clk_2_wires[107]),
    .prog_clk_0_N_in(prog_clk_0_wires[285]),
    .chany_top_in(cby_1__1__82_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_82_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_82_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_82_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_82_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_82_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_82_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_82_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_82_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__86_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_93_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_93_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_93_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_93_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_93_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_93_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_93_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_93_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__81_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_81_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_81_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_81_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_81_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_81_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_81_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_81_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_81_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__75_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_81_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_81_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_81_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_81_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_81_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_81_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_81_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_81_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__86_ccff_tail[0]),
    .chany_top_out(sb_1__1__75_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__75_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__75_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__75_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__75_ccff_tail[0])
  );


  sb_1__1_
  sb_7__11_
  (
    .clk_1_S_in(clk_2_wires[109]),
    .clk_1_W_out(clk_1_wires[163]),
    .clk_1_E_out(clk_1_wires[162]),
    .prog_clk_1_S_in(prog_clk_2_wires[109]),
    .prog_clk_1_W_out(prog_clk_1_wires[163]),
    .prog_clk_1_E_out(prog_clk_1_wires[162]),
    .prog_clk_0_N_in(prog_clk_0_wires[288]),
    .chany_top_in(cby_1__1__83_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_83_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_83_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_83_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_83_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_83_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_83_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_83_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_83_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__87_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_94_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_94_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_94_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_94_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_94_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_94_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_94_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_94_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__82_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_82_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_82_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_82_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_82_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_82_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_82_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_82_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_82_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__76_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_82_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_82_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_82_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_82_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_82_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_82_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_82_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_82_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__87_ccff_tail[0]),
    .chany_top_out(sb_1__1__76_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__76_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__76_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__76_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__76_ccff_tail[0])
  );


  sb_1__1_
  sb_8__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[296]),
    .chany_top_in(cby_1__1__85_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_85_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_85_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_85_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_85_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_85_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_85_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_85_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_85_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__88_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_96_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_96_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_96_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_96_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_96_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_96_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_96_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_96_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__84_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_84_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_84_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_84_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_84_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_84_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_84_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_84_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_84_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__77_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_84_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_84_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_84_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_84_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_84_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_84_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_84_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_84_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__88_ccff_tail[0]),
    .chany_top_out(sb_1__1__77_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__77_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__77_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__77_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__77_ccff_tail[0])
  );


  sb_1__1_
  sb_8__2_
  (
    .clk_2_N_in(clk_3_wires[43]),
    .clk_2_W_out(clk_2_wires[71]),
    .clk_2_E_out(clk_2_wires[69]),
    .prog_clk_2_N_in(prog_clk_3_wires[43]),
    .prog_clk_2_W_out(prog_clk_2_wires[71]),
    .prog_clk_2_E_out(prog_clk_2_wires[69]),
    .prog_clk_0_N_in(prog_clk_0_wires[299]),
    .chany_top_in(cby_1__1__86_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_86_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_86_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_86_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_86_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_86_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_86_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_86_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_86_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__89_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_97_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_97_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_97_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_97_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_97_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_97_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_97_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_97_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__85_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_85_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_85_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_85_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_85_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_85_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_85_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_85_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_85_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__78_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_85_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_85_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_85_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_85_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_85_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_85_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_85_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_85_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__89_ccff_tail[0]),
    .chany_top_out(sb_1__1__78_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__78_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__78_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__78_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__78_ccff_tail[0])
  );


  sb_1__1_
  sb_8__3_
  (
    .clk_3_S_out(clk_3_wires[42]),
    .clk_3_N_in(clk_3_wires[39]),
    .prog_clk_3_S_out(prog_clk_3_wires[42]),
    .prog_clk_3_N_in(prog_clk_3_wires[39]),
    .prog_clk_0_N_in(prog_clk_0_wires[302]),
    .chany_top_in(cby_1__1__87_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_87_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_87_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_87_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_87_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_87_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_87_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_87_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_87_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__90_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_98_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_98_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_98_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_98_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_98_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_98_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_98_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_98_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__86_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_86_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_86_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_86_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_86_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_86_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_86_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_86_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_86_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__79_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_86_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_86_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_86_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_86_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_86_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_86_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_86_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_86_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__90_ccff_tail[0]),
    .chany_top_out(sb_1__1__79_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__79_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__79_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__79_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__79_ccff_tail[0])
  );


  sb_1__1_
  sb_8__4_
  (
    .clk_3_S_out(clk_3_wires[38]),
    .clk_2_N_in(clk_3_wires[33]),
    .clk_3_N_in(clk_3_wires[33]),
    .clk_2_W_out(clk_2_wires[80]),
    .clk_2_E_out(clk_2_wires[78]),
    .prog_clk_3_S_out(prog_clk_3_wires[38]),
    .prog_clk_2_N_in(prog_clk_3_wires[33]),
    .prog_clk_3_N_in(prog_clk_3_wires[33]),
    .prog_clk_2_W_out(prog_clk_2_wires[80]),
    .prog_clk_2_E_out(prog_clk_2_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[305]),
    .chany_top_in(cby_1__1__88_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_88_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_88_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_88_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_88_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_88_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_88_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_88_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_88_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__91_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_99_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_99_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_99_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_99_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_99_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_99_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_99_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_99_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__87_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_87_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_87_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_87_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_87_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_87_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_87_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_87_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_87_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__80_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_87_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_87_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_87_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_87_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_87_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_87_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_87_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_87_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__91_ccff_tail[0]),
    .chany_top_out(sb_1__1__80_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__80_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__80_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__80_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__80_ccff_tail[0])
  );


  sb_1__1_
  sb_8__5_
  (
    .clk_3_S_out(clk_3_wires[32]),
    .clk_3_N_in(clk_3_wires[29]),
    .prog_clk_3_S_out(prog_clk_3_wires[32]),
    .prog_clk_3_N_in(prog_clk_3_wires[29]),
    .prog_clk_0_N_in(prog_clk_0_wires[308]),
    .chany_top_in(cby_1__1__89_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_89_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_89_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_89_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_89_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_89_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_89_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_89_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_89_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__92_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_100_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_100_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_100_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_100_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_100_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_100_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_100_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_100_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__88_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_88_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_88_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_88_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_88_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_88_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_88_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_88_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_88_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__81_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_88_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_88_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_88_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_88_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_88_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_88_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_88_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_88_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__92_ccff_tail[0]),
    .chany_top_out(sb_1__1__81_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__81_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__81_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__81_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__81_ccff_tail[0])
  );


  sb_1__1_
  sb_8__6_
  (
    .clk_3_E_out(clk_3_wires[44]),
    .clk_3_S_out(clk_3_wires[28]),
    .clk_3_N_out(clk_3_wires[26]),
    .clk_3_W_in(clk_3_wires[5]),
    .prog_clk_3_E_out(prog_clk_3_wires[44]),
    .prog_clk_3_S_out(prog_clk_3_wires[28]),
    .prog_clk_3_N_out(prog_clk_3_wires[26]),
    .prog_clk_3_W_in(prog_clk_3_wires[5]),
    .prog_clk_0_N_in(prog_clk_0_wires[311]),
    .chany_top_in(cby_1__1__90_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_90_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_90_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_90_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_90_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_90_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_90_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_90_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_90_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__93_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_101_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_101_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_101_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_101_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_101_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_101_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_101_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_101_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__89_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_89_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_89_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_89_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_89_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_89_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_89_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_89_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_89_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__82_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_89_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_89_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_89_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_89_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_89_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_89_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_89_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_89_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__93_ccff_tail[0]),
    .chany_top_out(sb_1__1__82_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__82_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__82_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__82_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__82_ccff_tail[0])
  );


  sb_1__1_
  sb_8__7_
  (
    .clk_3_N_out(clk_3_wires[30]),
    .clk_3_S_in(clk_3_wires[27]),
    .prog_clk_3_N_out(prog_clk_3_wires[30]),
    .prog_clk_3_S_in(prog_clk_3_wires[27]),
    .prog_clk_0_N_in(prog_clk_0_wires[314]),
    .chany_top_in(cby_1__1__91_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_91_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_91_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_91_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_91_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_91_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_91_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_91_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_91_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__94_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_102_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_102_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_102_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_102_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_102_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_102_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_102_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_102_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__90_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_90_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_90_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_90_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_90_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_90_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_90_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_90_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_90_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__83_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_90_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_90_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_90_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_90_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_90_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_90_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_90_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_90_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__94_ccff_tail[0]),
    .chany_top_out(sb_1__1__83_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__83_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__83_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__83_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__83_ccff_tail[0])
  );


  sb_1__1_
  sb_8__8_
  (
    .clk_3_N_out(clk_3_wires[36]),
    .clk_2_S_in(clk_3_wires[31]),
    .clk_3_S_in(clk_3_wires[31]),
    .clk_2_W_out(clk_2_wires[93]),
    .clk_2_E_out(clk_2_wires[91]),
    .prog_clk_3_N_out(prog_clk_3_wires[36]),
    .prog_clk_2_S_in(prog_clk_3_wires[31]),
    .prog_clk_3_S_in(prog_clk_3_wires[31]),
    .prog_clk_2_W_out(prog_clk_2_wires[93]),
    .prog_clk_2_E_out(prog_clk_2_wires[91]),
    .prog_clk_0_N_in(prog_clk_0_wires[317]),
    .chany_top_in(cby_1__1__92_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_92_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_92_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_92_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_92_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_92_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_92_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_92_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_92_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__95_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_103_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_103_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_103_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_103_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_103_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_103_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_103_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_103_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__91_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_91_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_91_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_91_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_91_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_91_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_91_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_91_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_91_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__84_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_91_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_91_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_91_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_91_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_91_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_91_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_91_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_91_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__95_ccff_tail[0]),
    .chany_top_out(sb_1__1__84_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__84_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__84_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__84_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__84_ccff_tail[0])
  );


  sb_1__1_
  sb_8__9_
  (
    .clk_3_N_out(clk_3_wires[40]),
    .clk_3_S_in(clk_3_wires[37]),
    .prog_clk_3_N_out(prog_clk_3_wires[40]),
    .prog_clk_3_S_in(prog_clk_3_wires[37]),
    .prog_clk_0_N_in(prog_clk_0_wires[320]),
    .chany_top_in(cby_1__1__93_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_93_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_93_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_93_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_93_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_93_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_93_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_93_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_93_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__96_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_104_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_104_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_104_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_104_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_104_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_104_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_104_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_104_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__92_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_92_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_92_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_92_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_92_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_92_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_92_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_92_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_92_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__85_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_92_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_92_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_92_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_92_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_92_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_92_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_92_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_92_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__96_ccff_tail[0]),
    .chany_top_out(sb_1__1__85_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__85_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__85_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__85_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__85_ccff_tail[0])
  );


  sb_1__1_
  sb_8__10_
  (
    .clk_2_S_in(clk_3_wires[41]),
    .clk_2_W_out(clk_2_wires[106]),
    .clk_2_E_out(clk_2_wires[104]),
    .prog_clk_2_S_in(prog_clk_3_wires[41]),
    .prog_clk_2_W_out(prog_clk_2_wires[106]),
    .prog_clk_2_E_out(prog_clk_2_wires[104]),
    .prog_clk_0_N_in(prog_clk_0_wires[323]),
    .chany_top_in(cby_1__1__94_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_94_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_94_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_94_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_94_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_94_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_94_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_94_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_94_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__97_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_105_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_105_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_105_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_105_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_105_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_105_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_105_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_105_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__93_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_93_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_93_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_93_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_93_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_93_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_93_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_93_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_93_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__86_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_93_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_93_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_93_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_93_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_93_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_93_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_93_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_93_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__97_ccff_tail[0]),
    .chany_top_out(sb_1__1__86_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__86_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__86_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__86_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__86_ccff_tail[0])
  );


  sb_1__1_
  sb_8__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[326]),
    .chany_top_in(cby_1__1__95_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_95_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_95_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_95_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_95_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_95_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_95_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_95_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_95_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__98_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_106_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_106_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_106_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_106_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_106_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_106_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_106_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_106_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__94_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_94_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_94_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_94_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_94_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_94_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_94_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_94_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_94_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__87_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_94_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_94_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_94_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_94_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_94_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_94_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_94_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_94_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__98_ccff_tail[0]),
    .chany_top_out(sb_1__1__87_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__87_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__87_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__87_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__87_ccff_tail[0])
  );


  sb_1__1_
  sb_9__1_
  (
    .clk_1_N_in(clk_2_wires[76]),
    .clk_1_W_out(clk_1_wires[170]),
    .clk_1_E_out(clk_1_wires[169]),
    .prog_clk_1_N_in(prog_clk_2_wires[76]),
    .prog_clk_1_W_out(prog_clk_1_wires[170]),
    .prog_clk_1_E_out(prog_clk_1_wires[169]),
    .prog_clk_0_N_in(prog_clk_0_wires[334]),
    .chany_top_in(cby_1__1__97_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_97_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_97_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_97_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_97_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_97_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_97_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_97_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_97_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__99_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_108_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_108_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_108_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_108_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_108_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_108_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_108_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_108_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__96_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_96_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_96_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_96_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_96_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_96_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_96_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_96_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_96_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__88_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_96_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_96_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_96_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_96_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_96_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_96_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_96_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_96_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__99_ccff_tail[0]),
    .chany_top_out(sb_1__1__88_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__88_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__88_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__88_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__88_ccff_tail[0])
  );


  sb_1__1_
  sb_9__2_
  (
    .clk_2_S_out(clk_2_wires[75]),
    .clk_2_W_in(clk_2_wires[70]),
    .prog_clk_2_S_out(prog_clk_2_wires[75]),
    .prog_clk_2_W_in(prog_clk_2_wires[70]),
    .prog_clk_0_N_in(prog_clk_0_wires[337]),
    .chany_top_in(cby_1__1__98_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_98_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_98_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_98_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_98_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_98_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_98_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_98_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_98_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__100_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_109_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_109_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_109_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_109_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_109_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_109_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_109_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_109_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__97_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_97_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_97_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_97_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_97_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_97_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_97_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_97_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_97_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__89_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_97_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_97_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_97_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_97_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_97_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_97_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_97_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_97_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__100_ccff_tail[0]),
    .chany_top_out(sb_1__1__89_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__89_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__89_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__89_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__89_ccff_tail[0])
  );


  sb_1__1_
  sb_9__3_
  (
    .clk_1_N_in(clk_2_wires[89]),
    .clk_1_W_out(clk_1_wires[177]),
    .clk_1_E_out(clk_1_wires[176]),
    .prog_clk_1_N_in(prog_clk_2_wires[89]),
    .prog_clk_1_W_out(prog_clk_1_wires[177]),
    .prog_clk_1_E_out(prog_clk_1_wires[176]),
    .prog_clk_0_N_in(prog_clk_0_wires[340]),
    .chany_top_in(cby_1__1__99_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_99_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_99_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_99_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_99_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_99_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_99_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_99_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_99_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__101_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_110_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_110_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_110_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_110_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_110_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_110_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_110_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_110_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__98_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_98_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_98_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_98_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_98_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_98_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_98_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_98_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_98_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__90_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_98_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_98_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_98_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_98_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_98_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_98_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_98_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_98_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__101_ccff_tail[0]),
    .chany_top_out(sb_1__1__90_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__90_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__90_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__90_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__90_ccff_tail[0])
  );


  sb_1__1_
  sb_9__4_
  (
    .clk_2_S_out(clk_2_wires[88]),
    .clk_2_N_out(clk_2_wires[86]),
    .clk_2_W_in(clk_2_wires[79]),
    .prog_clk_2_S_out(prog_clk_2_wires[88]),
    .prog_clk_2_N_out(prog_clk_2_wires[86]),
    .prog_clk_2_W_in(prog_clk_2_wires[79]),
    .prog_clk_0_N_in(prog_clk_0_wires[343]),
    .chany_top_in(cby_1__1__100_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_100_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_100_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_100_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_100_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_100_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_100_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_100_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_100_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__102_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_111_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_111_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_111_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_111_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_111_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_111_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_111_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_111_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__99_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_99_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_99_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_99_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_99_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_99_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_99_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_99_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_99_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__91_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_99_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_99_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_99_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_99_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_99_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_99_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_99_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_99_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__102_ccff_tail[0]),
    .chany_top_out(sb_1__1__91_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__91_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__91_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__91_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__91_ccff_tail[0])
  );


  sb_1__1_
  sb_9__5_
  (
    .clk_1_S_in(clk_2_wires[87]),
    .clk_1_W_out(clk_1_wires[184]),
    .clk_1_E_out(clk_1_wires[183]),
    .prog_clk_1_S_in(prog_clk_2_wires[87]),
    .prog_clk_1_W_out(prog_clk_1_wires[184]),
    .prog_clk_1_E_out(prog_clk_1_wires[183]),
    .prog_clk_0_N_in(prog_clk_0_wires[346]),
    .chany_top_in(cby_1__1__101_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_101_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_101_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_101_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_101_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_101_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_101_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_101_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_101_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__103_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_112_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_112_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_112_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_112_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_112_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_112_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_112_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_112_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__100_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_100_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_100_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_100_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_100_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_100_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_100_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_100_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_100_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__92_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_100_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_100_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_100_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_100_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_100_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_100_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_100_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_100_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__103_ccff_tail[0]),
    .chany_top_out(sb_1__1__92_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__92_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__92_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__92_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__92_ccff_tail[0])
  );


  sb_1__1_
  sb_9__6_
  (
    .clk_3_E_out(clk_3_wires[48]),
    .clk_3_W_in(clk_3_wires[45]),
    .prog_clk_3_E_out(prog_clk_3_wires[48]),
    .prog_clk_3_W_in(prog_clk_3_wires[45]),
    .prog_clk_0_N_in(prog_clk_0_wires[349]),
    .chany_top_in(cby_1__1__102_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_102_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_102_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_102_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_102_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_102_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_102_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_102_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_102_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__104_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_113_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_113_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_113_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_113_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_113_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_113_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_113_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_113_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__101_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_101_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_101_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_101_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_101_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_101_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_101_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_101_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_101_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__93_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_101_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_101_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_101_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_101_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_101_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_101_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_101_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_101_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__104_ccff_tail[0]),
    .chany_top_out(sb_1__1__93_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__93_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__93_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__93_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__93_ccff_tail[0])
  );


  sb_1__1_
  sb_9__7_
  (
    .clk_1_N_in(clk_2_wires[102]),
    .clk_1_W_out(clk_1_wires[191]),
    .clk_1_E_out(clk_1_wires[190]),
    .prog_clk_1_N_in(prog_clk_2_wires[102]),
    .prog_clk_1_W_out(prog_clk_1_wires[191]),
    .prog_clk_1_E_out(prog_clk_1_wires[190]),
    .prog_clk_0_N_in(prog_clk_0_wires[352]),
    .chany_top_in(cby_1__1__103_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_103_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_103_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_103_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_103_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_103_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_103_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_103_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_103_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__105_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_114_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_114_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_114_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_114_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_114_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_114_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_114_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_114_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__102_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_102_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_102_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_102_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_102_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_102_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_102_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_102_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_102_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__94_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_102_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_102_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_102_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_102_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_102_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_102_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_102_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_102_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__105_ccff_tail[0]),
    .chany_top_out(sb_1__1__94_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__94_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__94_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__94_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__94_ccff_tail[0])
  );


  sb_1__1_
  sb_9__8_
  (
    .clk_2_S_out(clk_2_wires[101]),
    .clk_2_N_out(clk_2_wires[99]),
    .clk_2_W_in(clk_2_wires[92]),
    .prog_clk_2_S_out(prog_clk_2_wires[101]),
    .prog_clk_2_N_out(prog_clk_2_wires[99]),
    .prog_clk_2_W_in(prog_clk_2_wires[92]),
    .prog_clk_0_N_in(prog_clk_0_wires[355]),
    .chany_top_in(cby_1__1__104_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_104_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_104_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_104_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_104_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_104_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_104_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_104_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_104_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__106_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_115_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_115_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_115_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_115_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_115_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_115_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_115_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_115_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__103_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_103_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_103_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_103_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_103_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_103_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_103_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_103_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_103_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__95_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_103_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_103_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_103_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_103_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_103_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_103_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_103_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_103_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__106_ccff_tail[0]),
    .chany_top_out(sb_1__1__95_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__95_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__95_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__95_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__95_ccff_tail[0])
  );


  sb_1__1_
  sb_9__9_
  (
    .clk_1_S_in(clk_2_wires[100]),
    .clk_1_W_out(clk_1_wires[198]),
    .clk_1_E_out(clk_1_wires[197]),
    .prog_clk_1_S_in(prog_clk_2_wires[100]),
    .prog_clk_1_W_out(prog_clk_1_wires[198]),
    .prog_clk_1_E_out(prog_clk_1_wires[197]),
    .prog_clk_0_N_in(prog_clk_0_wires[358]),
    .chany_top_in(cby_1__1__105_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_105_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_105_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_105_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_105_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_105_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_105_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_105_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_105_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__107_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_116_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_116_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_116_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_116_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_116_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_116_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_116_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_116_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__104_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_104_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_104_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_104_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_104_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_104_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_104_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_104_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_104_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__96_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_104_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_104_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_104_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_104_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_104_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_104_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_104_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_104_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__107_ccff_tail[0]),
    .chany_top_out(sb_1__1__96_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__96_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__96_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__96_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__96_ccff_tail[0])
  );


  sb_1__1_
  sb_9__10_
  (
    .clk_2_N_out(clk_2_wires[110]),
    .clk_2_W_in(clk_2_wires[105]),
    .prog_clk_2_N_out(prog_clk_2_wires[110]),
    .prog_clk_2_W_in(prog_clk_2_wires[105]),
    .prog_clk_0_N_in(prog_clk_0_wires[361]),
    .chany_top_in(cby_1__1__106_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_106_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_106_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_106_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_106_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_106_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_106_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_106_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_106_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__108_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_117_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_117_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_117_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_117_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_117_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_117_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_117_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_117_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__105_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_105_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_105_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_105_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_105_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_105_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_105_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_105_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_105_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__97_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_105_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_105_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_105_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_105_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_105_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_105_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_105_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_105_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__108_ccff_tail[0]),
    .chany_top_out(sb_1__1__97_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__97_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__97_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__97_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__97_ccff_tail[0])
  );


  sb_1__1_
  sb_9__11_
  (
    .clk_1_S_in(clk_2_wires[111]),
    .clk_1_W_out(clk_1_wires[205]),
    .clk_1_E_out(clk_1_wires[204]),
    .prog_clk_1_S_in(prog_clk_2_wires[111]),
    .prog_clk_1_W_out(prog_clk_1_wires[205]),
    .prog_clk_1_E_out(prog_clk_1_wires[204]),
    .prog_clk_0_N_in(prog_clk_0_wires[364]),
    .chany_top_in(cby_1__1__107_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_107_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_107_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_107_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_107_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_107_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_107_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_107_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_107_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__109_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_118_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_118_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_118_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_118_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_118_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_118_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_118_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_118_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__106_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_106_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_106_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_106_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_106_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_106_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_106_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_106_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_106_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__98_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_106_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_106_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_106_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_106_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_106_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_106_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_106_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_106_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__109_ccff_tail[0]),
    .chany_top_out(sb_1__1__98_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__98_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__98_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__98_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__98_ccff_tail[0])
  );


  sb_1__1_
  sb_10__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[372]),
    .chany_top_in(cby_1__1__109_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_109_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_109_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_109_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_109_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_109_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_109_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_109_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_109_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__110_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_120_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_120_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_120_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_120_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_120_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_120_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_120_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_120_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__108_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_108_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_108_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_108_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_108_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_108_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_108_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_108_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_108_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__99_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_108_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_108_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_108_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_108_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_108_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_108_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_108_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_108_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__110_ccff_tail[0]),
    .chany_top_out(sb_1__1__99_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__99_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__99_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__99_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__99_ccff_tail[0])
  );


  sb_1__1_
  sb_10__2_
  (
    .clk_2_N_in(clk_3_wires[87]),
    .clk_2_E_out(clk_2_wires[114]),
    .prog_clk_2_N_in(prog_clk_3_wires[87]),
    .prog_clk_2_E_out(prog_clk_2_wires[114]),
    .prog_clk_0_N_in(prog_clk_0_wires[375]),
    .chany_top_in(cby_1__1__110_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_110_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_110_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_110_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_110_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_110_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_110_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_110_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_110_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__111_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_121_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_121_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_121_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_121_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_121_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_121_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_121_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_121_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__109_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_109_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_109_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_109_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_109_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_109_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_109_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_109_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_109_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__100_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_109_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_109_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_109_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_109_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_109_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_109_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_109_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_109_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__111_ccff_tail[0]),
    .chany_top_out(sb_1__1__100_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__100_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__100_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__100_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__100_ccff_tail[0])
  );


  sb_1__1_
  sb_10__3_
  (
    .clk_3_S_out(clk_3_wires[86]),
    .clk_3_N_in(clk_3_wires[83]),
    .prog_clk_3_S_out(prog_clk_3_wires[86]),
    .prog_clk_3_N_in(prog_clk_3_wires[83]),
    .prog_clk_0_N_in(prog_clk_0_wires[378]),
    .chany_top_in(cby_1__1__111_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_111_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_111_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_111_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_111_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_111_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_111_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_111_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_111_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__112_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_122_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_122_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_122_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_122_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_122_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_122_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_122_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_122_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__110_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_110_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_110_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_110_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_110_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_110_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_110_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_110_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_110_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__101_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_110_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_110_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_110_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_110_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_110_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_110_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_110_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_110_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__112_ccff_tail[0]),
    .chany_top_out(sb_1__1__101_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__101_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__101_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__101_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__101_ccff_tail[0])
  );


  sb_1__1_
  sb_10__4_
  (
    .clk_3_S_out(clk_3_wires[82]),
    .clk_2_N_in(clk_3_wires[77]),
    .clk_3_N_in(clk_3_wires[77]),
    .clk_2_E_out(clk_2_wires[119]),
    .prog_clk_3_S_out(prog_clk_3_wires[82]),
    .prog_clk_2_N_in(prog_clk_3_wires[77]),
    .prog_clk_3_N_in(prog_clk_3_wires[77]),
    .prog_clk_2_E_out(prog_clk_2_wires[119]),
    .prog_clk_0_N_in(prog_clk_0_wires[381]),
    .chany_top_in(cby_1__1__112_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_112_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_112_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_112_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_112_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_112_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_112_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_112_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_112_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__113_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_123_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_123_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_123_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_123_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_123_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_123_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_123_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_123_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__111_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_111_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_111_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_111_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_111_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_111_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_111_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_111_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_111_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__102_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_111_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_111_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_111_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_111_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_111_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_111_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_111_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_111_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__113_ccff_tail[0]),
    .chany_top_out(sb_1__1__102_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__102_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__102_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__102_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__102_ccff_tail[0])
  );


  sb_1__1_
  sb_10__5_
  (
    .clk_3_S_out(clk_3_wires[76]),
    .clk_3_N_in(clk_3_wires[73]),
    .prog_clk_3_S_out(prog_clk_3_wires[76]),
    .prog_clk_3_N_in(prog_clk_3_wires[73]),
    .prog_clk_0_N_in(prog_clk_0_wires[384]),
    .chany_top_in(cby_1__1__113_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_113_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_113_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_113_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_113_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_113_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_113_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_113_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_113_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__114_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_124_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_124_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_124_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_124_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_124_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_124_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_124_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_124_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__112_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_112_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_112_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_112_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_112_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_112_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_112_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_112_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_112_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__103_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_112_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_112_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_112_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_112_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_112_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_112_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_112_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_112_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__114_ccff_tail[0]),
    .chany_top_out(sb_1__1__103_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__103_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__103_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__103_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__103_ccff_tail[0])
  );


  sb_1__1_
  sb_10__6_
  (
    .clk_3_S_out(clk_3_wires[72]),
    .clk_3_N_out(clk_3_wires[70]),
    .clk_3_W_in(clk_3_wires[49]),
    .prog_clk_3_S_out(prog_clk_3_wires[72]),
    .prog_clk_3_N_out(prog_clk_3_wires[70]),
    .prog_clk_3_W_in(prog_clk_3_wires[49]),
    .prog_clk_0_N_in(prog_clk_0_wires[387]),
    .chany_top_in(cby_1__1__114_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_114_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_114_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_114_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_114_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_114_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_114_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_114_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_114_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__115_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_125_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_125_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_125_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_125_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_125_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_125_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_125_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_125_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__113_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_113_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_113_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_113_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_113_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_113_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_113_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_113_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_113_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__104_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_113_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_113_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_113_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_113_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_113_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_113_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_113_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_113_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__115_ccff_tail[0]),
    .chany_top_out(sb_1__1__104_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__104_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__104_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__104_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__104_ccff_tail[0])
  );


  sb_1__1_
  sb_10__7_
  (
    .clk_3_N_out(clk_3_wires[74]),
    .clk_3_S_in(clk_3_wires[71]),
    .prog_clk_3_N_out(prog_clk_3_wires[74]),
    .prog_clk_3_S_in(prog_clk_3_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[390]),
    .chany_top_in(cby_1__1__115_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_115_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_115_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_115_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_115_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_115_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_115_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_115_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_115_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__116_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_126_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_126_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_126_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_126_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_126_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_126_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_126_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_126_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__114_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_114_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_114_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_114_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_114_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_114_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_114_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_114_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_114_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__105_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_114_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_114_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_114_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_114_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_114_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_114_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_114_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_114_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__116_ccff_tail[0]),
    .chany_top_out(sb_1__1__105_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__105_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__105_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__105_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__105_ccff_tail[0])
  );


  sb_1__1_
  sb_10__8_
  (
    .clk_3_N_out(clk_3_wires[80]),
    .clk_2_S_in(clk_3_wires[75]),
    .clk_3_S_in(clk_3_wires[75]),
    .clk_2_E_out(clk_2_wires[126]),
    .prog_clk_3_N_out(prog_clk_3_wires[80]),
    .prog_clk_2_S_in(prog_clk_3_wires[75]),
    .prog_clk_3_S_in(prog_clk_3_wires[75]),
    .prog_clk_2_E_out(prog_clk_2_wires[126]),
    .prog_clk_0_N_in(prog_clk_0_wires[393]),
    .chany_top_in(cby_1__1__116_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_116_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_116_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_116_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_116_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_116_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_116_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_116_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_116_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__117_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_127_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_127_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_127_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_127_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_127_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_127_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_127_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_127_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__115_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_115_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_115_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_115_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_115_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_115_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_115_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_115_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_115_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__106_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_115_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_115_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_115_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_115_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_115_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_115_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_115_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_115_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__117_ccff_tail[0]),
    .chany_top_out(sb_1__1__106_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__106_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__106_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__106_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__106_ccff_tail[0])
  );


  sb_1__1_
  sb_10__9_
  (
    .clk_3_N_out(clk_3_wires[84]),
    .clk_3_S_in(clk_3_wires[81]),
    .prog_clk_3_N_out(prog_clk_3_wires[84]),
    .prog_clk_3_S_in(prog_clk_3_wires[81]),
    .prog_clk_0_N_in(prog_clk_0_wires[396]),
    .chany_top_in(cby_1__1__117_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_117_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_117_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_117_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_117_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_117_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_117_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_117_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_117_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__118_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_128_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_128_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_128_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_128_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_128_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_128_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_128_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_128_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__116_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_116_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_116_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_116_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_116_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_116_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_116_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_116_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_116_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__107_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_116_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_116_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_116_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_116_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_116_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_116_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_116_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_116_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__118_ccff_tail[0]),
    .chany_top_out(sb_1__1__107_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__107_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__107_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__107_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__107_ccff_tail[0])
  );


  sb_1__1_
  sb_10__10_
  (
    .clk_2_S_in(clk_3_wires[85]),
    .clk_2_E_out(clk_2_wires[133]),
    .prog_clk_2_S_in(prog_clk_3_wires[85]),
    .prog_clk_2_E_out(prog_clk_2_wires[133]),
    .prog_clk_0_N_in(prog_clk_0_wires[399]),
    .chany_top_in(cby_1__1__118_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_118_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_118_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_118_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_118_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_118_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_118_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_118_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_118_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__119_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_129_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_129_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_129_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_129_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_129_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_129_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_129_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_129_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__117_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_117_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_117_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_117_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_117_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_117_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_117_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_117_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_117_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__108_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_117_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_117_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_117_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_117_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_117_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_117_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_117_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_117_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__119_ccff_tail[0]),
    .chany_top_out(sb_1__1__108_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__108_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__108_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__108_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__108_ccff_tail[0])
  );


  sb_1__1_
  sb_10__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[402]),
    .chany_top_in(cby_1__1__119_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_119_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_119_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_119_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_119_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_119_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_119_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_119_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_119_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__120_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_130_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_130_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_130_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_130_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_130_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_130_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_130_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_130_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__118_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_118_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_118_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_118_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_118_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_118_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_118_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_118_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_118_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__109_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_118_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_118_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_118_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_118_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_118_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_118_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_118_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_118_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__120_ccff_tail[0]),
    .chany_top_out(sb_1__1__109_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__109_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__109_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__109_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__109_ccff_tail[0])
  );


  sb_1__1_
  sb_11__1_
  (
    .clk_1_N_in(clk_2_wires[116]),
    .clk_1_W_out(clk_1_wires[212]),
    .clk_1_E_out(clk_1_wires[211]),
    .prog_clk_1_N_in(prog_clk_2_wires[116]),
    .prog_clk_1_W_out(prog_clk_1_wires[212]),
    .prog_clk_1_E_out(prog_clk_1_wires[211]),
    .prog_clk_0_N_in(prog_clk_0_wires[410]),
    .chany_top_in(cby_1__1__121_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_121_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_121_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_121_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_121_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_121_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_121_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_121_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_121_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__121_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_132_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_132_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_132_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_132_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_132_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_132_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_132_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_132_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__120_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_120_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_120_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_120_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_120_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_120_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_120_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_120_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_120_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__110_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_120_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_120_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_120_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_120_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_120_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_120_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_120_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_120_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__121_ccff_tail[0]),
    .chany_top_out(sb_1__1__110_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__110_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__110_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__110_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__110_ccff_tail[0])
  );


  sb_1__1_
  sb_11__2_
  (
    .clk_2_S_out(clk_2_wires[115]),
    .clk_2_W_in(clk_2_wires[113]),
    .prog_clk_2_S_out(prog_clk_2_wires[115]),
    .prog_clk_2_W_in(prog_clk_2_wires[113]),
    .prog_clk_0_N_in(prog_clk_0_wires[413]),
    .chany_top_in(cby_1__1__122_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_122_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_122_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_122_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_122_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_122_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_122_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_122_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_122_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__122_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_133_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_133_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_133_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_133_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_133_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_133_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_133_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_133_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__121_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_121_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_121_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_121_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_121_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_121_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_121_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_121_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_121_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__111_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_121_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_121_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_121_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_121_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_121_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_121_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_121_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_121_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__122_ccff_tail[0]),
    .chany_top_out(sb_1__1__111_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__111_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__111_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__111_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__111_ccff_tail[0])
  );


  sb_1__1_
  sb_11__3_
  (
    .clk_1_N_in(clk_2_wires[123]),
    .clk_1_W_out(clk_1_wires[219]),
    .clk_1_E_out(clk_1_wires[218]),
    .prog_clk_1_N_in(prog_clk_2_wires[123]),
    .prog_clk_1_W_out(prog_clk_1_wires[219]),
    .prog_clk_1_E_out(prog_clk_1_wires[218]),
    .prog_clk_0_N_in(prog_clk_0_wires[416]),
    .chany_top_in(cby_1__1__123_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_123_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_123_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_123_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_123_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_123_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_123_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_123_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_123_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__123_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_134_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_134_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_134_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_134_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_134_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_134_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_134_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_134_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__122_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_122_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_122_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_122_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_122_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_122_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_122_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_122_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_122_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__112_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_122_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_122_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_122_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_122_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_122_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_122_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_122_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_122_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__123_ccff_tail[0]),
    .chany_top_out(sb_1__1__112_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__112_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__112_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__112_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__112_ccff_tail[0])
  );


  sb_1__1_
  sb_11__4_
  (
    .clk_2_S_out(clk_2_wires[122]),
    .clk_2_N_out(clk_2_wires[120]),
    .clk_2_W_in(clk_2_wires[118]),
    .prog_clk_2_S_out(prog_clk_2_wires[122]),
    .prog_clk_2_N_out(prog_clk_2_wires[120]),
    .prog_clk_2_W_in(prog_clk_2_wires[118]),
    .prog_clk_0_N_in(prog_clk_0_wires[419]),
    .chany_top_in(cby_1__1__124_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_124_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_124_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_124_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_124_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_124_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_124_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_124_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_124_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__124_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_135_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_135_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_135_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_135_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_135_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_135_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_135_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_135_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__123_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_123_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_123_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_123_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_123_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_123_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_123_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_123_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_123_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__113_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_123_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_123_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_123_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_123_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_123_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_123_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_123_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_123_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__124_ccff_tail[0]),
    .chany_top_out(sb_1__1__113_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__113_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__113_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__113_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__113_ccff_tail[0])
  );


  sb_1__1_
  sb_11__5_
  (
    .clk_1_S_in(clk_2_wires[121]),
    .clk_1_W_out(clk_1_wires[226]),
    .clk_1_E_out(clk_1_wires[225]),
    .prog_clk_1_S_in(prog_clk_2_wires[121]),
    .prog_clk_1_W_out(prog_clk_1_wires[226]),
    .prog_clk_1_E_out(prog_clk_1_wires[225]),
    .prog_clk_0_N_in(prog_clk_0_wires[422]),
    .chany_top_in(cby_1__1__125_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_125_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_125_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_125_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_125_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_125_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_125_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_125_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_125_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__125_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_136_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_136_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_136_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_136_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_136_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_136_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_136_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_136_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__124_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_124_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_124_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_124_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_124_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_124_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_124_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_124_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_124_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__114_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_124_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_124_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_124_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_124_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_124_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_124_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_124_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_124_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__125_ccff_tail[0]),
    .chany_top_out(sb_1__1__114_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__114_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__114_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__114_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__114_ccff_tail[0])
  );


  sb_1__1_
  sb_11__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[425]),
    .chany_top_in(cby_1__1__126_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_126_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_126_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_126_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_126_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_126_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_126_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_126_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_126_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__126_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_137_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_137_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_137_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_137_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_137_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_137_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_137_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_137_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__125_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_125_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_125_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_125_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_125_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_125_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_125_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_125_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_125_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__115_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_125_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_125_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_125_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_125_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_125_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_125_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_125_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_125_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__126_ccff_tail[0]),
    .chany_top_out(sb_1__1__115_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__115_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__115_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__115_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__115_ccff_tail[0])
  );


  sb_1__1_
  sb_11__7_
  (
    .clk_1_N_in(clk_2_wires[130]),
    .clk_1_W_out(clk_1_wires[233]),
    .clk_1_E_out(clk_1_wires[232]),
    .prog_clk_1_N_in(prog_clk_2_wires[130]),
    .prog_clk_1_W_out(prog_clk_1_wires[233]),
    .prog_clk_1_E_out(prog_clk_1_wires[232]),
    .prog_clk_0_N_in(prog_clk_0_wires[428]),
    .chany_top_in(cby_1__1__127_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_127_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_127_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_127_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_127_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_127_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_127_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_127_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_127_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__127_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_138_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_138_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_138_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_138_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_138_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_138_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_138_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_138_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__126_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_126_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_126_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_126_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_126_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_126_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_126_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_126_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_126_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__116_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_126_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_126_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_126_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_126_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_126_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_126_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_126_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_126_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__127_ccff_tail[0]),
    .chany_top_out(sb_1__1__116_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__116_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__116_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__116_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__116_ccff_tail[0])
  );


  sb_1__1_
  sb_11__8_
  (
    .clk_2_S_out(clk_2_wires[129]),
    .clk_2_N_out(clk_2_wires[127]),
    .clk_2_W_in(clk_2_wires[125]),
    .prog_clk_2_S_out(prog_clk_2_wires[129]),
    .prog_clk_2_N_out(prog_clk_2_wires[127]),
    .prog_clk_2_W_in(prog_clk_2_wires[125]),
    .prog_clk_0_N_in(prog_clk_0_wires[431]),
    .chany_top_in(cby_1__1__128_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_128_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_128_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_128_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_128_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_128_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_128_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_128_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_128_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__128_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_139_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_139_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_139_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_139_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_139_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_139_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_139_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_139_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__127_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_127_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_127_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_127_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_127_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_127_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_127_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_127_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_127_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__117_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_127_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_127_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_127_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_127_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_127_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_127_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_127_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_127_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__128_ccff_tail[0]),
    .chany_top_out(sb_1__1__117_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__117_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__117_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__117_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__117_ccff_tail[0])
  );


  sb_1__1_
  sb_11__9_
  (
    .clk_1_S_in(clk_2_wires[128]),
    .clk_1_W_out(clk_1_wires[240]),
    .clk_1_E_out(clk_1_wires[239]),
    .prog_clk_1_S_in(prog_clk_2_wires[128]),
    .prog_clk_1_W_out(prog_clk_1_wires[240]),
    .prog_clk_1_E_out(prog_clk_1_wires[239]),
    .prog_clk_0_N_in(prog_clk_0_wires[434]),
    .chany_top_in(cby_1__1__129_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_129_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_129_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_129_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_129_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_129_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_129_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_129_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_129_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__129_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_140_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_140_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_140_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_140_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_140_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_140_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_140_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_140_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__128_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_128_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_128_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_128_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_128_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_128_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_128_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_128_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_128_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__118_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_128_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_128_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_128_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_128_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_128_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_128_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_128_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_128_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__129_ccff_tail[0]),
    .chany_top_out(sb_1__1__118_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__118_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__118_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__118_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__118_ccff_tail[0])
  );


  sb_1__1_
  sb_11__10_
  (
    .clk_2_N_out(clk_2_wires[134]),
    .clk_2_W_in(clk_2_wires[132]),
    .prog_clk_2_N_out(prog_clk_2_wires[134]),
    .prog_clk_2_W_in(prog_clk_2_wires[132]),
    .prog_clk_0_N_in(prog_clk_0_wires[437]),
    .chany_top_in(cby_1__1__130_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_130_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_130_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_130_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_130_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_130_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_130_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_130_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_130_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__130_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_141_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_141_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_141_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_141_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_141_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_141_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_141_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_141_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__129_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_129_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_129_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_129_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_129_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_129_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_129_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_129_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_129_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__119_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_129_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_129_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_129_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_129_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_129_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_129_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_129_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_129_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__130_ccff_tail[0]),
    .chany_top_out(sb_1__1__119_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__119_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__119_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__119_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__119_ccff_tail[0])
  );


  sb_1__1_
  sb_11__11_
  (
    .clk_1_S_in(clk_2_wires[135]),
    .clk_1_W_out(clk_1_wires[247]),
    .clk_1_E_out(clk_1_wires[246]),
    .prog_clk_1_S_in(prog_clk_2_wires[135]),
    .prog_clk_1_W_out(prog_clk_1_wires[247]),
    .prog_clk_1_E_out(prog_clk_1_wires[246]),
    .prog_clk_0_N_in(prog_clk_0_wires[440]),
    .chany_top_in(cby_1__1__131_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_131_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_131_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_131_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_131_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_131_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_131_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_131_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_131_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__131_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_142_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_142_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_142_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_142_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_142_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_142_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_142_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_142_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__130_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_130_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_130_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_130_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_130_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_130_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_130_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_130_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_130_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__120_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_130_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_130_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_130_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_130_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_130_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_130_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_130_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_130_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__131_ccff_tail[0]),
    .chany_top_out(sb_1__1__120_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__120_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__120_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__120_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__120_ccff_tail[0])
  );


  sb_1__2_
  sb_1__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[60]),
    .chanx_right_in(cbx_1__12__1_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_1_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_23_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_23_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_23_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_23_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_23_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_23_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_23_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_23_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__11_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_11_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_11_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_11_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_11_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_11_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_11_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_11_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_11_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__12__0_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_0_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_11_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_11_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_11_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_11_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_11_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_11_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_11_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_11_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_1_ccff_tail[0]),
    .chanx_right_out(sb_1__12__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__0_ccff_tail[0])
  );


  sb_1__2_
  sb_2__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[100]),
    .SC_OUT_BOT(scff_Wires[53]),
    .SC_IN_BOT(scff_Wires[52]),
    .chanx_right_in(cbx_1__12__2_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_2_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_35_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_35_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_35_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_35_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_35_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_35_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_35_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_35_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__23_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_23_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_23_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_23_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_23_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_23_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_23_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_23_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_23_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__12__1_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_1_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_23_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_23_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_23_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_23_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_23_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_23_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_23_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_23_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_2_ccff_tail[0]),
    .chanx_right_out(sb_1__12__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__1_ccff_tail[0])
  );


  sb_1__2_
  sb_3__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[138]),
    .chanx_right_in(cbx_1__12__3_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_3_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_47_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_47_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_47_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_47_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_47_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_47_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_47_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_47_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__35_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_35_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_35_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_35_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_35_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_35_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_35_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_35_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_35_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__12__2_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_2_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_35_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_35_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_35_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_35_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_35_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_35_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_35_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_35_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_3_ccff_tail[0]),
    .chanx_right_out(sb_1__12__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__2_ccff_tail[0])
  );


  sb_1__2_
  sb_4__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[176]),
    .SC_OUT_BOT(scff_Wires[106]),
    .SC_IN_BOT(scff_Wires[105]),
    .chanx_right_in(cbx_1__12__4_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_4_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_59_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_59_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_59_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_59_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_59_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_59_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_59_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_59_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__47_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_47_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_47_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_47_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_47_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_47_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_47_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_47_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_47_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__12__3_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_3_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_47_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_47_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_47_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_47_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_47_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_47_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_47_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_47_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_4_ccff_tail[0]),
    .chanx_right_out(sb_1__12__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__3_ccff_tail[0])
  );


  sb_1__2_
  sb_5__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[214]),
    .chanx_right_in(cbx_1__12__5_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_5_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_71_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_71_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_71_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_71_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_71_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_71_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_71_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_71_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__59_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_59_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_59_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_59_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_59_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_59_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_59_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_59_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_59_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__12__4_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_4_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_59_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_59_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_59_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_59_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_59_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_59_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_59_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_59_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_5_ccff_tail[0]),
    .chanx_right_out(sb_1__12__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__4_ccff_tail[0])
  );


  sb_1__2_
  sb_6__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[252]),
    .SC_OUT_BOT(scff_Wires[159]),
    .SC_IN_BOT(scff_Wires[158]),
    .chanx_right_in(cbx_1__12__6_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_6_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_83_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_83_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_83_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_83_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_83_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_83_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_83_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_83_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__71_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_71_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_71_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_71_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_71_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_71_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_71_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_71_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_71_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__12__5_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_5_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_71_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_71_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_71_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_71_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_71_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_71_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_71_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_71_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_6_ccff_tail[0]),
    .chanx_right_out(sb_1__12__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__5_ccff_tail[0])
  );


  sb_1__2_
  sb_7__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[290]),
    .chanx_right_in(cbx_1__12__7_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_7_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_95_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_95_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_95_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_95_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_95_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_95_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_95_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_95_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__83_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_83_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_83_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_83_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_83_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_83_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_83_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_83_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_83_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__12__6_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_6_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_83_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_83_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_83_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_83_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_83_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_83_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_83_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_83_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_7_ccff_tail[0]),
    .chanx_right_out(sb_1__12__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__6_ccff_tail[0])
  );


  sb_1__2_
  sb_8__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[328]),
    .SC_OUT_BOT(scff_Wires[212]),
    .SC_IN_BOT(scff_Wires[211]),
    .chanx_right_in(cbx_1__12__8_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_8_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_107_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_107_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_107_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_107_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_107_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_107_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_107_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_107_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__95_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_95_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_95_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_95_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_95_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_95_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_95_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_95_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_95_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__12__7_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_7_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_95_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_95_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_95_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_95_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_95_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_95_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_95_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_95_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_8_ccff_tail[0]),
    .chanx_right_out(sb_1__12__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__7_ccff_tail[0])
  );


  sb_1__2_
  sb_9__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[366]),
    .chanx_right_in(cbx_1__12__9_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_9_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_119_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_119_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_119_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_119_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_119_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_119_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_119_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_119_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__107_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_107_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_107_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_107_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_107_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_107_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_107_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_107_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_107_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__12__8_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_8_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_107_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_107_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_107_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_107_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_107_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_107_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_107_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_107_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_9_ccff_tail[0]),
    .chanx_right_out(sb_1__12__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__8_ccff_tail[0])
  );


  sb_1__2_
  sb_10__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[404]),
    .SC_OUT_BOT(scff_Wires[265]),
    .SC_IN_BOT(scff_Wires[264]),
    .chanx_right_in(cbx_1__12__10_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_10_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_131_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_131_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_131_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_131_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_131_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_131_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_131_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_131_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__119_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_119_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_119_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_119_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_119_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_119_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_119_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_119_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_119_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__12__9_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_9_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_119_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_119_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_119_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_119_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_119_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_119_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_119_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_119_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_10_ccff_tail[0]),
    .chanx_right_out(sb_1__12__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__9_ccff_tail[0])
  );


  sb_1__2_
  sb_11__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[442]),
    .chanx_right_in(cbx_1__12__11_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_11_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_143_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_143_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_143_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_143_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_143_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_143_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_143_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_143_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__131_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_131_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_131_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_131_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_131_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_131_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_131_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_131_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_131_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__12__10_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_10_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_131_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_131_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_131_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_131_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_131_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_131_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_131_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_131_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_11_ccff_tail[0]),
    .chanx_right_out(sb_1__12__10_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__12__10_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__12__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__12__10_ccff_tail[0])
  );


  sb_2__0_
  sb_12__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[445]),
    .chany_top_in(cby_12__1__0_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_132_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_132_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_132_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_132_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_132_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_132_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_132_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_132_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_11_left_width_0_height_0__pin_1_lower[0]),
    .chanx_left_in(cbx_1__0__11_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_0_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_0_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_0_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_0_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_0_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_0_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_0_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_0_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_0_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_right_11_ccff_tail[0]),
    .chany_top_out(sb_12__0__0_chany_top_out[0:19]),
    .chanx_left_out(sb_12__0__0_chanx_left_out[0:19]),
    .ccff_tail(sb_12__0__0_ccff_tail[0])
  );


  sb_2__1_
  sb_12__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[448]),
    .chany_top_in(cby_12__1__1_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_133_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_133_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_133_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_133_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_133_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_133_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_133_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_133_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_10_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__0_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_11_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_132_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_132_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_132_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_132_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_132_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_132_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_132_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_132_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__121_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_132_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_132_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_132_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_132_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_132_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_132_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_132_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_132_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_10_ccff_tail[0]),
    .chany_top_out(sb_12__1__0_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__0_chanx_left_out[0:19]),
    .ccff_tail(sb_12__1__0_ccff_tail[0])
  );


  sb_2__1_
  sb_12__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[451]),
    .chany_top_in(cby_12__1__2_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_134_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_134_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_134_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_134_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_134_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_134_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_134_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_134_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_9_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__1_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_10_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_133_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_133_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_133_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_133_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_133_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_133_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_133_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_133_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__122_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_133_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_133_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_133_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_133_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_133_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_133_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_133_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_133_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_9_ccff_tail[0]),
    .chany_top_out(sb_12__1__1_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__1_chanx_left_out[0:19]),
    .ccff_tail(sb_12__1__1_ccff_tail[0])
  );


  sb_2__1_
  sb_12__3_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[454]),
    .chany_top_in(cby_12__1__3_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_135_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_135_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_135_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_135_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_135_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_135_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_135_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_135_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_8_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__2_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_9_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_134_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_134_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_134_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_134_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_134_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_134_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_134_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_134_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__123_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_134_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_134_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_134_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_134_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_134_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_134_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_134_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_134_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_8_ccff_tail[0]),
    .chany_top_out(sb_12__1__2_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__2_chanx_left_out[0:19]),
    .ccff_tail(sb_12__1__2_ccff_tail[0])
  );


  sb_2__1_
  sb_12__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[457]),
    .chany_top_in(cby_12__1__4_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_136_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_136_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_136_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_136_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_136_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_136_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_136_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_136_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_7_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__3_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_8_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_135_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_135_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_135_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_135_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_135_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_135_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_135_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_135_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__124_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_135_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_135_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_135_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_135_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_135_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_135_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_135_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_135_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_7_ccff_tail[0]),
    .chany_top_out(sb_12__1__3_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__3_chanx_left_out[0:19]),
    .ccff_tail(sb_12__1__3_ccff_tail[0])
  );


  sb_2__1_
  sb_12__5_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[460]),
    .chany_top_in(cby_12__1__5_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_137_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_137_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_137_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_137_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_137_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_137_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_137_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_137_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_6_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__4_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_7_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_136_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_136_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_136_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_136_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_136_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_136_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_136_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_136_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__125_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_136_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_136_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_136_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_136_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_136_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_136_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_136_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_136_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_6_ccff_tail[0]),
    .chany_top_out(sb_12__1__4_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__4_chanx_left_out[0:19]),
    .ccff_tail(sb_12__1__4_ccff_tail[0])
  );


  sb_2__1_
  sb_12__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[463]),
    .chany_top_in(cby_12__1__6_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_138_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_138_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_138_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_138_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_138_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_138_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_138_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_138_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_5_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__5_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_6_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_137_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_137_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_137_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_137_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_137_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_137_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_137_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_137_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__126_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_137_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_137_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_137_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_137_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_137_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_137_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_137_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_137_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_5_ccff_tail[0]),
    .chany_top_out(sb_12__1__5_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__5_chanx_left_out[0:19]),
    .ccff_tail(sb_12__1__5_ccff_tail[0])
  );


  sb_2__1_
  sb_12__7_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[466]),
    .chany_top_in(cby_12__1__7_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_139_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_139_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_139_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_139_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_139_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_139_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_139_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_139_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_4_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__6_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_5_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_138_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_138_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_138_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_138_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_138_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_138_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_138_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_138_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__127_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_138_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_138_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_138_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_138_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_138_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_138_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_138_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_138_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_4_ccff_tail[0]),
    .chany_top_out(sb_12__1__6_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__6_chanx_left_out[0:19]),
    .ccff_tail(sb_12__1__6_ccff_tail[0])
  );


  sb_2__1_
  sb_12__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[469]),
    .chany_top_in(cby_12__1__8_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_140_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_140_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_140_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_140_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_140_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_140_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_140_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_140_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_3_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__7_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_4_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_139_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_139_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_139_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_139_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_139_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_139_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_139_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_139_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__128_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_139_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_139_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_139_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_139_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_139_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_139_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_139_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_139_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_3_ccff_tail[0]),
    .chany_top_out(sb_12__1__7_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__7_chanx_left_out[0:19]),
    .ccff_tail(sb_12__1__7_ccff_tail[0])
  );


  sb_2__1_
  sb_12__9_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[472]),
    .chany_top_in(cby_12__1__9_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_141_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_141_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_141_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_141_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_141_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_141_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_141_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_141_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_2_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__8_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_3_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_140_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_140_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_140_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_140_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_140_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_140_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_140_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_140_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__129_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_140_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_140_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_140_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_140_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_140_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_140_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_140_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_140_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_2_ccff_tail[0]),
    .chany_top_out(sb_12__1__8_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__8_chanx_left_out[0:19]),
    .ccff_tail(sb_12__1__8_ccff_tail[0])
  );


  sb_2__1_
  sb_12__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[475]),
    .chany_top_in(cby_12__1__10_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_142_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_142_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_142_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_142_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_142_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_142_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_142_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_142_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_1_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__9_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_2_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_141_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_141_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_141_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_141_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_141_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_141_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_141_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_141_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__130_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_141_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_141_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_141_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_141_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_141_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_141_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_141_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_141_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_1_ccff_tail[0]),
    .chany_top_out(sb_12__1__9_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__9_chanx_left_out[0:19]),
    .ccff_tail(sb_12__1__9_ccff_tail[0])
  );


  sb_2__1_
  sb_12__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[478]),
    .chany_top_in(cby_12__1__11_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_143_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_143_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_143_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_143_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_143_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_143_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_143_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_143_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_0_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__10_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_1_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_142_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_142_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_142_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_142_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_142_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_142_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_142_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_142_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__131_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_142_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_142_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_142_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_142_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_142_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_142_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_142_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_142_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_0_ccff_tail[0]),
    .chany_top_out(sb_12__1__10_chany_top_out[0:19]),
    .chany_bottom_out(sb_12__1__10_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__1__10_chanx_left_out[0:19]),
    .ccff_tail(sb_12__1__10_ccff_tail[0])
  );


  sb_2__2_
  sb_12__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[480]),
    .SC_OUT_BOT(sc_tail),
    .SC_IN_BOT(scff_Wires[317]),
    .chany_bottom_in(cby_12__1__11_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_0_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_143_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_143_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_143_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_143_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_143_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_143_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_143_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_143_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__12__11_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_11_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_143_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_143_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_143_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_143_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_143_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_143_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_143_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_143_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(ccff_head[0]),
    .chany_bottom_out(sb_12__12__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_12__12__0_chanx_left_out[0:19]),
    .ccff_tail(sb_12__12__0_ccff_tail[0])
  );


  cbx_1__0_
  cbx_1__0_
  (
    .prog_clk_0_W_out(prog_clk_0_wires[5]),
    .prog_clk_0_N_in(prog_clk_0_wires[0]),
    .SC_OUT_BOT(scff_Wires[26]),
    .SC_IN_TOP(scff_Wires[25]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_11_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_11_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_11_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_11_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_11_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_11_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_11_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_11_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_11_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_11_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_11_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_11_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_11_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_11_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_11_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_11_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_11_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_11_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__0_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__0_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__0_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__0_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__0_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__0_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__0_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__0_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__0_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[123:131]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[123:131]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[123:131]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_0__0__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__0_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__0_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__0_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__0_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__0_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__0_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__0_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__0_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__0_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__0_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_11_ccff_tail[0])
  );


  cbx_1__0_
  cbx_2__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[63]),
    .SC_OUT_TOP(scff_Wires[28]),
    .SC_IN_BOT(scff_Wires[27]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_10_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_10_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_10_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_10_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_10_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_10_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_10_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_10_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_10_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_10_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_10_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_10_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_10_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_10_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_10_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_10_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_10_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_10_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__1_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__1_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__1_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__1_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__1_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__1_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__1_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__1_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__1_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[114:122]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[114:122]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[114:122]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__1_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__1_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__1_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__1_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__1_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__1_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__1_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__1_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__1_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__1_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__1_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_10_ccff_tail[0])
  );


  cbx_1__0_
  cbx_3__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[101]),
    .SC_OUT_BOT(scff_Wires[79]),
    .SC_IN_TOP(scff_Wires[78]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_9_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_9_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_9_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_9_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_9_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_9_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_9_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_9_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_9_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_9_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_9_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_9_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_9_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_9_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_9_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_9_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_9_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_9_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__2_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__2_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__2_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__2_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__2_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__2_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__2_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__2_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__2_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[105:113]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[105:113]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[105:113]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__2_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__2_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__2_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__2_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__2_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__2_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__2_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__2_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__2_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__2_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__2_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_9_ccff_tail[0])
  );


  cbx_1__0_
  cbx_4__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[139]),
    .SC_OUT_TOP(scff_Wires[81]),
    .SC_IN_BOT(scff_Wires[80]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_8_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_8_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_8_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_8_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_8_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_8_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_8_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_8_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_8_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_8_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_8_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_8_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_8_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_8_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_8_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_8_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_8_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_8_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__3_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__3_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__3_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__3_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__3_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__3_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__3_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__3_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__3_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[96:104]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[96:104]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[96:104]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__3_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__3_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__3_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__3_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__3_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__3_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__3_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__3_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__3_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__3_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__3_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_8_ccff_tail[0])
  );


  cbx_1__0_
  cbx_5__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[177]),
    .SC_OUT_BOT(scff_Wires[132]),
    .SC_IN_TOP(scff_Wires[131]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_7_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_7_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_7_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_7_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_7_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_7_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_7_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_7_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_7_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_7_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_7_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_7_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_7_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_7_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_7_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_7_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_7_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_7_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__4_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__4_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__4_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__4_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__4_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__4_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__4_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__4_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__4_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87:95]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87:95]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87:95]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__4_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__4_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__4_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__4_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__4_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__4_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__4_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__4_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__4_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__4_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__4_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_7_ccff_tail[0])
  );


  cbx_1__0_
  cbx_6__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[215]),
    .SC_OUT_TOP(scff_Wires[134]),
    .SC_IN_BOT(scff_Wires[133]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_6_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_6_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_6_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_6_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_6_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_6_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_6_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_6_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_6_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_6_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_6_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_6_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_6_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_6_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_6_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_6_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_6_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_6_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__5_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__5_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__5_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__5_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__5_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__5_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__5_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__5_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__5_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78:86]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78:86]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78:86]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__5_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__5_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__5_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__5_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__5_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__5_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__5_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__5_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__5_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__5_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__5_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_6_ccff_tail[0])
  );


  cbx_1__0_
  cbx_7__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[253]),
    .SC_OUT_BOT(scff_Wires[185]),
    .SC_IN_TOP(scff_Wires[184]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_5_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_5_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_5_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_5_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_5_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_5_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_5_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_5_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_5_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_5_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_5_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_5_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_5_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_5_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_5_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_5_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_5_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_5_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__6_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__6_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__6_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__6_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__6_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__6_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__6_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__6_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__6_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69:77]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69:77]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69:77]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__6_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__6_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__6_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__6_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__6_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__6_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__6_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__6_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__6_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__6_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__6_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_5_ccff_tail[0])
  );


  cbx_1__0_
  cbx_8__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[291]),
    .SC_OUT_TOP(scff_Wires[187]),
    .SC_IN_BOT(scff_Wires[186]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_4_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_4_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_4_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_4_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_4_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_4_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_4_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_4_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_4_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_4_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_4_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_4_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_4_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_4_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_4_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_4_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_4_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_4_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__7_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__7_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__7_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__7_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__7_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__7_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__7_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__7_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__7_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60:68]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60:68]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60:68]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__7_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__7_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__7_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__7_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__7_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__7_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__7_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__7_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__7_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__7_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__7_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__7_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_4_ccff_tail[0])
  );


  cbx_1__0_
  cbx_9__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[329]),
    .SC_OUT_BOT(scff_Wires[238]),
    .SC_IN_TOP(scff_Wires[237]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_3_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_3_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_3_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_3_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_3_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_3_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_3_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_3_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_3_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_3_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_3_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_3_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_3_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_3_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_3_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_3_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_3_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_3_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__8_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__8_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__8_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__8_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__8_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__8_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__8_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__8_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__8_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51:59]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51:59]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51:59]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__8_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__8_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__8_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__8_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__8_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__8_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__8_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__8_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__8_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__8_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__8_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__8_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_3_ccff_tail[0])
  );


  cbx_1__0_
  cbx_10__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[367]),
    .SC_OUT_TOP(scff_Wires[240]),
    .SC_IN_BOT(scff_Wires[239]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_2_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_2_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_2_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_2_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_2_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_2_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_2_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_2_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_2_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_2_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_2_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_2_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_2_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_2_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_2_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_2_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_2_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_2_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__9_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__9_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__9_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__9_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__9_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__9_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__9_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__9_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__9_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42:50]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42:50]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42:50]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__9_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__9_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__9_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__9_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__9_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__9_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__9_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__9_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__9_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__9_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__9_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__9_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_2_ccff_tail[0])
  );


  cbx_1__0_
  cbx_11__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[405]),
    .SC_OUT_BOT(scff_Wires[291]),
    .SC_IN_TOP(scff_Wires[290]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_1_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_1_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_1_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_1_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_1_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_1_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_1_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_1_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_1_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_1_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_1_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_1_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_1_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_1_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_1_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_1_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_1_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_1_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__10_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__10_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__10_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__10_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__10_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__10_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__10_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__10_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__10_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33:41]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33:41]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33:41]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__10_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__10_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__10_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__10_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__10_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__10_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__10_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__10_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__10_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__10_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__10_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__10_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_1_ccff_tail[0])
  );


  cbx_1__0_
  cbx_12__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[443]),
    .SC_OUT_TOP(scff_Wires[293]),
    .SC_IN_BOT(scff_Wires[292]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_0_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_0_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_0_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_0_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_0_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_0_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_0_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_0_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_0_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_0_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_0_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_0_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_0_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_0_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_0_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_0_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_0_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_0_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__11_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__11_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__11_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__11_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__11_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__11_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__11_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__11_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__11_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24:32]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24:32]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24:32]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__0__0_chanx_left_out[0:19]),
    .ccff_head(sb_12__0__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__11_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__11_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__11_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__11_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__11_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__11_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__11_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__11_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__11_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__11_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_0_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__1_
  (
    .clk_1_S_out(clk_1_wires[4]),
    .clk_1_N_out(clk_1_wires[3]),
    .clk_1_E_in(clk_1_wires[2]),
    .prog_clk_1_S_out(prog_clk_1_wires[4]),
    .prog_clk_1_N_out(prog_clk_1_wires[3]),
    .prog_clk_1_E_in(prog_clk_1_wires[2]),
    .prog_clk_0_N_in(prog_clk_0_wires[6]),
    .prog_clk_0_W_out(prog_clk_0_wires[4]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[0]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[0]),
    .SC_OUT_BOT(scff_Wires[23]),
    .SC_IN_TOP(scff_Wires[22]),
    .chanx_left_in(sb_0__1__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__0_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__0_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__0_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__0_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__0_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__0_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__0_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__0_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__0_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__0_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__0_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__0_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__0_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__0_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__0_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__0_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__0_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__0_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[11]),
    .prog_clk_0_W_out(prog_clk_0_wires[10]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[1]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[1]),
    .SC_OUT_BOT(scff_Wires[21]),
    .SC_IN_TOP(scff_Wires[20]),
    .chanx_left_in(sb_0__1__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__1_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__1_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__1_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__1_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__1_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__1_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__1_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__1_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__1_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__1_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__1_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__1_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__1_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__1_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__1_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__1_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__1_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__1_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__1_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__3_
  (
    .clk_1_S_out(clk_1_wires[11]),
    .clk_1_N_out(clk_1_wires[10]),
    .clk_1_E_in(clk_1_wires[9]),
    .prog_clk_1_S_out(prog_clk_1_wires[11]),
    .prog_clk_1_N_out(prog_clk_1_wires[10]),
    .prog_clk_1_E_in(prog_clk_1_wires[9]),
    .prog_clk_0_N_in(prog_clk_0_wires[16]),
    .prog_clk_0_W_out(prog_clk_0_wires[15]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[2]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[2]),
    .SC_OUT_BOT(scff_Wires[19]),
    .SC_IN_TOP(scff_Wires[18]),
    .chanx_left_in(sb_0__1__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__2_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__2_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__2_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__2_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__2_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__2_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__2_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__2_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__2_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__2_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__2_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__2_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__2_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__2_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__2_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__2_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__2_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__2_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__2_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[21]),
    .prog_clk_0_W_out(prog_clk_0_wires[20]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[3]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[3]),
    .SC_OUT_BOT(scff_Wires[17]),
    .SC_IN_TOP(scff_Wires[16]),
    .chanx_left_in(sb_0__1__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__3_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__3_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__3_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__3_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__3_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__3_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__3_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__3_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__3_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__3_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__3_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__3_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__3_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__3_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__3_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__3_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__3_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__3_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__3_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__5_
  (
    .clk_1_S_out(clk_1_wires[18]),
    .clk_1_N_out(clk_1_wires[17]),
    .clk_1_E_in(clk_1_wires[16]),
    .prog_clk_1_S_out(prog_clk_1_wires[18]),
    .prog_clk_1_N_out(prog_clk_1_wires[17]),
    .prog_clk_1_E_in(prog_clk_1_wires[16]),
    .prog_clk_0_N_in(prog_clk_0_wires[26]),
    .prog_clk_0_W_out(prog_clk_0_wires[25]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[4]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[4]),
    .SC_OUT_BOT(scff_Wires[15]),
    .SC_IN_TOP(scff_Wires[14]),
    .chanx_left_in(sb_0__1__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__4_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__4_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__4_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__4_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__4_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__4_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__4_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__4_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__4_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__4_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__4_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__4_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__4_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__4_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__4_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__4_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__4_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__4_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__4_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[31]),
    .prog_clk_0_W_out(prog_clk_0_wires[30]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[5]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[5]),
    .SC_OUT_BOT(scff_Wires[13]),
    .SC_IN_TOP(scff_Wires[12]),
    .chanx_left_in(sb_0__1__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__5_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__5_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__5_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__5_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__5_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__5_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__5_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__5_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__5_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__5_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__5_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__5_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__5_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__5_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__5_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__5_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__5_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__5_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__5_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__7_
  (
    .clk_1_S_out(clk_1_wires[25]),
    .clk_1_N_out(clk_1_wires[24]),
    .clk_1_E_in(clk_1_wires[23]),
    .prog_clk_1_S_out(prog_clk_1_wires[25]),
    .prog_clk_1_N_out(prog_clk_1_wires[24]),
    .prog_clk_1_E_in(prog_clk_1_wires[23]),
    .prog_clk_0_N_in(prog_clk_0_wires[36]),
    .prog_clk_0_W_out(prog_clk_0_wires[35]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[6]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[6]),
    .SC_OUT_BOT(scff_Wires[11]),
    .SC_IN_TOP(scff_Wires[10]),
    .chanx_left_in(sb_0__1__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__6_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__6_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__6_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__6_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__6_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__6_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__6_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__6_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__6_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__6_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__6_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__6_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__6_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__6_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__6_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__6_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__6_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__6_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__6_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[41]),
    .prog_clk_0_W_out(prog_clk_0_wires[40]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[7]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[7]),
    .SC_OUT_BOT(scff_Wires[9]),
    .SC_IN_TOP(scff_Wires[8]),
    .chanx_left_in(sb_0__1__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__7_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__7_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__7_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__7_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__7_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__7_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__7_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__7_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__7_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__7_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__7_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__7_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__7_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__7_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__7_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__7_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__7_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__7_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__7_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__7_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__9_
  (
    .clk_1_S_out(clk_1_wires[32]),
    .clk_1_N_out(clk_1_wires[31]),
    .clk_1_E_in(clk_1_wires[30]),
    .prog_clk_1_S_out(prog_clk_1_wires[32]),
    .prog_clk_1_N_out(prog_clk_1_wires[31]),
    .prog_clk_1_E_in(prog_clk_1_wires[30]),
    .prog_clk_0_N_in(prog_clk_0_wires[46]),
    .prog_clk_0_W_out(prog_clk_0_wires[45]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[8]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[8]),
    .SC_OUT_BOT(scff_Wires[7]),
    .SC_IN_TOP(scff_Wires[6]),
    .chanx_left_in(sb_0__1__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__8_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__8_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__8_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__8_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__8_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__8_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__8_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__8_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__8_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__8_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__8_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__8_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__8_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__8_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__8_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__8_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__8_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__8_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__8_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__8_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[51]),
    .prog_clk_0_W_out(prog_clk_0_wires[50]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[9]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[9]),
    .SC_OUT_BOT(scff_Wires[5]),
    .SC_IN_TOP(scff_Wires[4]),
    .chanx_left_in(sb_0__1__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__9_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__9_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__9_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__9_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__9_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__9_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__9_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__9_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__9_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__9_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__9_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__9_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__9_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__9_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__9_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__9_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__9_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__9_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__9_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__9_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__11_
  (
    .clk_1_S_out(clk_1_wires[39]),
    .clk_1_N_out(clk_1_wires[38]),
    .clk_1_E_in(clk_1_wires[37]),
    .prog_clk_1_S_out(prog_clk_1_wires[39]),
    .prog_clk_1_N_out(prog_clk_1_wires[38]),
    .prog_clk_1_E_in(prog_clk_1_wires[37]),
    .prog_clk_0_N_in(prog_clk_0_wires[56]),
    .prog_clk_0_W_out(prog_clk_0_wires[55]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[10]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[10]),
    .SC_OUT_BOT(scff_Wires[3]),
    .SC_IN_TOP(scff_Wires[2]),
    .chanx_left_in(sb_0__1__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__10_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__10_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__10_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__10_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__10_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__10_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__10_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__10_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__10_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__10_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__10_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__10_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__10_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__10_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__10_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__10_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__10_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__10_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__10_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__10_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__1_
  (
    .clk_1_S_out(clk_1_wires[6]),
    .clk_1_N_out(clk_1_wires[5]),
    .clk_1_W_in(clk_1_wires[1]),
    .prog_clk_1_S_out(prog_clk_1_wires[6]),
    .prog_clk_1_N_out(prog_clk_1_wires[5]),
    .prog_clk_1_W_in(prog_clk_1_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[66]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[11]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[11]),
    .SC_OUT_TOP(scff_Wires[30]),
    .SC_IN_BOT(scff_Wires[29]),
    .chanx_left_in(sb_1__1__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__11_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__11_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__11_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__11_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__11_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__11_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__11_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__11_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__11_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__11_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__11_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__11_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__11_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__11_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__11_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__11_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__11_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__11_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__11_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__11_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__2_
  (
    .clk_2_E_in(clk_2_wires[2]),
    .clk_2_W_out(clk_2_wires[1]),
    .prog_clk_2_E_in(prog_clk_2_wires[2]),
    .prog_clk_2_W_out(prog_clk_2_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[69]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[12]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[12]),
    .SC_OUT_TOP(scff_Wires[32]),
    .SC_IN_BOT(scff_Wires[31]),
    .chanx_left_in(sb_1__1__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__12_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__12_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__12_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__12_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__12_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__12_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__12_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__12_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__12_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__12_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__12_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__12_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__12_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__12_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__12_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__12_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__12_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__12_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__12_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__12_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__12_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__3_
  (
    .clk_1_S_out(clk_1_wires[13]),
    .clk_1_N_out(clk_1_wires[12]),
    .clk_1_W_in(clk_1_wires[8]),
    .prog_clk_1_S_out(prog_clk_1_wires[13]),
    .prog_clk_1_N_out(prog_clk_1_wires[12]),
    .prog_clk_1_W_in(prog_clk_1_wires[8]),
    .prog_clk_0_N_in(prog_clk_0_wires[72]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[13]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[13]),
    .SC_OUT_TOP(scff_Wires[34]),
    .SC_IN_BOT(scff_Wires[33]),
    .chanx_left_in(sb_1__1__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__13_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__13_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__13_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__13_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__13_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__13_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__13_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__13_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__13_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__13_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__13_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__13_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__13_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__13_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__13_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__13_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__13_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__13_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__13_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__13_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__13_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__4_
  (
    .clk_2_E_in(clk_2_wires[7]),
    .clk_2_W_out(clk_2_wires[6]),
    .prog_clk_2_E_in(prog_clk_2_wires[7]),
    .prog_clk_2_W_out(prog_clk_2_wires[6]),
    .prog_clk_0_N_in(prog_clk_0_wires[75]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[14]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[14]),
    .SC_OUT_TOP(scff_Wires[36]),
    .SC_IN_BOT(scff_Wires[35]),
    .chanx_left_in(sb_1__1__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__14_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__14_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__14_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__14_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__14_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__14_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__14_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__14_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__14_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__14_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__14_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__14_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__14_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__14_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__14_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__14_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__14_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__14_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__14_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__14_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__14_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__5_
  (
    .clk_1_S_out(clk_1_wires[20]),
    .clk_1_N_out(clk_1_wires[19]),
    .clk_1_W_in(clk_1_wires[15]),
    .prog_clk_1_S_out(prog_clk_1_wires[20]),
    .prog_clk_1_N_out(prog_clk_1_wires[19]),
    .prog_clk_1_W_in(prog_clk_1_wires[15]),
    .prog_clk_0_N_in(prog_clk_0_wires[78]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[15]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[15]),
    .SC_OUT_TOP(scff_Wires[38]),
    .SC_IN_BOT(scff_Wires[37]),
    .chanx_left_in(sb_1__1__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__15_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__15_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__15_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__15_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__15_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__15_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__15_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__15_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__15_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__15_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__15_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__15_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__15_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__15_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__15_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__15_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__15_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__15_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__15_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__15_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__15_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[81]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[16]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[16]),
    .SC_OUT_TOP(scff_Wires[40]),
    .SC_IN_BOT(scff_Wires[39]),
    .chanx_left_in(sb_1__1__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__16_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__16_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__16_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__16_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__16_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__16_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__16_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__16_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__16_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__16_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__16_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__16_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__16_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__16_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__16_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__16_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__16_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__16_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__16_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__16_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__16_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__7_
  (
    .clk_1_S_out(clk_1_wires[27]),
    .clk_1_N_out(clk_1_wires[26]),
    .clk_1_W_in(clk_1_wires[22]),
    .prog_clk_1_S_out(prog_clk_1_wires[27]),
    .prog_clk_1_N_out(prog_clk_1_wires[26]),
    .prog_clk_1_W_in(prog_clk_1_wires[22]),
    .prog_clk_0_N_in(prog_clk_0_wires[84]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[17]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[17]),
    .SC_OUT_TOP(scff_Wires[42]),
    .SC_IN_BOT(scff_Wires[41]),
    .chanx_left_in(sb_1__1__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__17_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__17_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__17_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__17_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__17_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__17_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__17_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__17_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__17_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__17_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__17_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__17_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__17_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__17_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__17_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__17_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__17_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__17_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__17_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__17_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__17_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__8_
  (
    .clk_2_E_in(clk_2_wires[14]),
    .clk_2_W_out(clk_2_wires[13]),
    .prog_clk_2_E_in(prog_clk_2_wires[14]),
    .prog_clk_2_W_out(prog_clk_2_wires[13]),
    .prog_clk_0_N_in(prog_clk_0_wires[87]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[18]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[18]),
    .SC_OUT_TOP(scff_Wires[44]),
    .SC_IN_BOT(scff_Wires[43]),
    .chanx_left_in(sb_1__1__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__18_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__18_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__18_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__18_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__18_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__18_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__18_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__18_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__18_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__18_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__18_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__18_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__18_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__18_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__18_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__18_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__18_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__18_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__18_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__18_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__18_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__9_
  (
    .clk_1_S_out(clk_1_wires[34]),
    .clk_1_N_out(clk_1_wires[33]),
    .clk_1_W_in(clk_1_wires[29]),
    .prog_clk_1_S_out(prog_clk_1_wires[34]),
    .prog_clk_1_N_out(prog_clk_1_wires[33]),
    .prog_clk_1_W_in(prog_clk_1_wires[29]),
    .prog_clk_0_N_in(prog_clk_0_wires[90]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[19]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[19]),
    .SC_OUT_TOP(scff_Wires[46]),
    .SC_IN_BOT(scff_Wires[45]),
    .chanx_left_in(sb_1__1__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__19_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__19_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__19_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__19_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__19_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__19_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__19_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__19_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__19_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__19_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__19_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__19_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__19_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__19_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__19_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__19_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__19_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__19_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__19_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__19_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__19_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__10_
  (
    .clk_2_E_in(clk_2_wires[21]),
    .clk_2_W_out(clk_2_wires[20]),
    .prog_clk_2_E_in(prog_clk_2_wires[21]),
    .prog_clk_2_W_out(prog_clk_2_wires[20]),
    .prog_clk_0_N_in(prog_clk_0_wires[93]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[20]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[20]),
    .SC_OUT_TOP(scff_Wires[48]),
    .SC_IN_BOT(scff_Wires[47]),
    .chanx_left_in(sb_1__1__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__20_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__20_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__20_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__20_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__20_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__20_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__20_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__20_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__20_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__20_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__20_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__20_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__20_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__20_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__20_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__20_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__20_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__20_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__20_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__20_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__20_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__11_
  (
    .clk_1_S_out(clk_1_wires[41]),
    .clk_1_N_out(clk_1_wires[40]),
    .clk_1_W_in(clk_1_wires[36]),
    .prog_clk_1_S_out(prog_clk_1_wires[41]),
    .prog_clk_1_N_out(prog_clk_1_wires[40]),
    .prog_clk_1_W_in(prog_clk_1_wires[36]),
    .prog_clk_0_N_in(prog_clk_0_wires[96]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[21]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[21]),
    .SC_OUT_TOP(scff_Wires[50]),
    .SC_IN_BOT(scff_Wires[49]),
    .chanx_left_in(sb_1__1__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__21_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__21_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__21_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__21_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__21_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__21_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__21_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__21_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__21_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__21_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__21_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__21_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__21_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__21_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__21_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__21_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__21_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__21_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__21_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__21_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__21_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__1_
  (
    .clk_1_S_out(clk_1_wires[46]),
    .clk_1_N_out(clk_1_wires[45]),
    .clk_1_E_in(clk_1_wires[44]),
    .prog_clk_1_S_out(prog_clk_1_wires[46]),
    .prog_clk_1_N_out(prog_clk_1_wires[45]),
    .prog_clk_1_E_in(prog_clk_1_wires[44]),
    .prog_clk_0_N_in(prog_clk_0_wires[104]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[22]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[22]),
    .SC_OUT_BOT(scff_Wires[76]),
    .SC_IN_TOP(scff_Wires[75]),
    .chanx_left_in(sb_1__1__11_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__22_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__22_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__22_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__22_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__22_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__22_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__22_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__22_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__22_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__22_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__22_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__22_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__22_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__22_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__22_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__22_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__22_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__22_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__22_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__22_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__22_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[107]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[23]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[23]),
    .SC_OUT_BOT(scff_Wires[74]),
    .SC_IN_TOP(scff_Wires[73]),
    .chanx_left_in(sb_1__1__12_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__23_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__23_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__23_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__23_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__23_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__23_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__23_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__23_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__23_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__23_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__23_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__23_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__23_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__23_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__23_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__23_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__23_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__23_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__23_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__23_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__23_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__3_
  (
    .clk_1_S_out(clk_1_wires[53]),
    .clk_1_N_out(clk_1_wires[52]),
    .clk_1_E_in(clk_1_wires[51]),
    .prog_clk_1_S_out(prog_clk_1_wires[53]),
    .prog_clk_1_N_out(prog_clk_1_wires[52]),
    .prog_clk_1_E_in(prog_clk_1_wires[51]),
    .prog_clk_0_N_in(prog_clk_0_wires[110]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[24]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[24]),
    .SC_OUT_BOT(scff_Wires[72]),
    .SC_IN_TOP(scff_Wires[71]),
    .chanx_left_in(sb_1__1__13_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__24_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__24_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__24_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__24_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__24_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__24_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__24_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__24_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__24_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__24_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__24_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__24_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__24_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__24_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__24_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__24_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__24_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__24_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__24_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__24_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__24_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[113]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[25]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[25]),
    .SC_OUT_BOT(scff_Wires[70]),
    .SC_IN_TOP(scff_Wires[69]),
    .chanx_left_in(sb_1__1__14_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__25_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__25_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__25_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__25_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__25_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__25_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__25_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__25_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__25_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__25_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__25_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__25_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__25_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__25_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__25_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__25_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__25_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__25_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__25_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__25_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__25_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__5_
  (
    .clk_1_S_out(clk_1_wires[60]),
    .clk_1_N_out(clk_1_wires[59]),
    .clk_1_E_in(clk_1_wires[58]),
    .prog_clk_1_S_out(prog_clk_1_wires[60]),
    .prog_clk_1_N_out(prog_clk_1_wires[59]),
    .prog_clk_1_E_in(prog_clk_1_wires[58]),
    .prog_clk_0_N_in(prog_clk_0_wires[116]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[26]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[26]),
    .SC_OUT_BOT(scff_Wires[68]),
    .SC_IN_TOP(scff_Wires[67]),
    .chanx_left_in(sb_1__1__15_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__26_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__26_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__26_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__26_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__26_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__26_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__26_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__26_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__26_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__26_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__26_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__26_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__26_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__26_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__26_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__26_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__26_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__26_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__26_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__26_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__26_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__6_
  (
    .clk_3_W_out(clk_3_wires[51]),
    .clk_3_E_in(clk_3_wires[50]),
    .prog_clk_3_W_out(prog_clk_3_wires[51]),
    .prog_clk_3_E_in(prog_clk_3_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[119]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[27]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[27]),
    .SC_OUT_BOT(scff_Wires[66]),
    .SC_IN_TOP(scff_Wires[65]),
    .chanx_left_in(sb_1__1__16_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__27_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__27_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__27_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__27_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__27_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__27_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__27_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__27_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__27_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__27_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__27_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__27_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__27_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__27_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__27_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__27_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__27_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__27_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__27_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__27_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__27_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__7_
  (
    .clk_1_S_out(clk_1_wires[67]),
    .clk_1_N_out(clk_1_wires[66]),
    .clk_1_E_in(clk_1_wires[65]),
    .prog_clk_1_S_out(prog_clk_1_wires[67]),
    .prog_clk_1_N_out(prog_clk_1_wires[66]),
    .prog_clk_1_E_in(prog_clk_1_wires[65]),
    .prog_clk_0_N_in(prog_clk_0_wires[122]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[28]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[28]),
    .SC_OUT_BOT(scff_Wires[64]),
    .SC_IN_TOP(scff_Wires[63]),
    .chanx_left_in(sb_1__1__17_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__28_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__28_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__28_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__28_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__28_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__28_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__28_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__28_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__28_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__28_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__28_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__28_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__28_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__28_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__28_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__28_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__28_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__28_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__28_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__28_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__28_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[125]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[29]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[29]),
    .SC_OUT_BOT(scff_Wires[62]),
    .SC_IN_TOP(scff_Wires[61]),
    .chanx_left_in(sb_1__1__18_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__29_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__29_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__29_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__29_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__29_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__29_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__29_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__29_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__29_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__29_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__29_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__29_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__29_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__29_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__29_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__29_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__29_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__29_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__29_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__29_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__29_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__9_
  (
    .clk_1_S_out(clk_1_wires[74]),
    .clk_1_N_out(clk_1_wires[73]),
    .clk_1_E_in(clk_1_wires[72]),
    .prog_clk_1_S_out(prog_clk_1_wires[74]),
    .prog_clk_1_N_out(prog_clk_1_wires[73]),
    .prog_clk_1_E_in(prog_clk_1_wires[72]),
    .prog_clk_0_N_in(prog_clk_0_wires[128]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[30]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[30]),
    .SC_OUT_BOT(scff_Wires[60]),
    .SC_IN_TOP(scff_Wires[59]),
    .chanx_left_in(sb_1__1__19_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__30_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__30_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__30_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__30_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__30_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__30_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__30_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__30_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__30_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__30_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__30_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__30_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__30_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__30_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__30_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__30_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__30_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__30_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__30_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__30_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__30_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[131]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[31]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[31]),
    .SC_OUT_BOT(scff_Wires[58]),
    .SC_IN_TOP(scff_Wires[57]),
    .chanx_left_in(sb_1__1__20_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__31_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__31_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__31_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__31_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__31_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__31_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__31_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__31_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__31_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__31_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__31_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__31_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__31_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__31_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__31_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__31_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__31_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__31_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__31_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__31_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__31_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__11_
  (
    .clk_1_S_out(clk_1_wires[81]),
    .clk_1_N_out(clk_1_wires[80]),
    .clk_1_E_in(clk_1_wires[79]),
    .prog_clk_1_S_out(prog_clk_1_wires[81]),
    .prog_clk_1_N_out(prog_clk_1_wires[80]),
    .prog_clk_1_E_in(prog_clk_1_wires[79]),
    .prog_clk_0_N_in(prog_clk_0_wires[134]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[32]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[32]),
    .SC_OUT_BOT(scff_Wires[56]),
    .SC_IN_TOP(scff_Wires[55]),
    .chanx_left_in(sb_1__1__21_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__32_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__32_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__32_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__32_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__32_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__32_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__32_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__32_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__32_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__32_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__32_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__32_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__32_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__32_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__32_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__32_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__32_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__32_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__32_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__32_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__32_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__1_
  (
    .clk_1_S_out(clk_1_wires[48]),
    .clk_1_N_out(clk_1_wires[47]),
    .clk_1_W_in(clk_1_wires[43]),
    .prog_clk_1_S_out(prog_clk_1_wires[48]),
    .prog_clk_1_N_out(prog_clk_1_wires[47]),
    .prog_clk_1_W_in(prog_clk_1_wires[43]),
    .prog_clk_0_N_in(prog_clk_0_wires[142]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[33]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[33]),
    .SC_OUT_TOP(scff_Wires[83]),
    .SC_IN_BOT(scff_Wires[82]),
    .chanx_left_in(sb_1__1__22_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__33_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__33_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__33_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__33_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__33_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__33_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__33_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__33_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__33_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__33_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__33_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__33_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__33_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__33_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__33_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__33_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__33_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__33_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__33_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__33_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__33_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__2_
  (
    .clk_2_W_out(clk_2_wires[28]),
    .clk_2_E_in(clk_2_wires[27]),
    .prog_clk_2_W_out(prog_clk_2_wires[28]),
    .prog_clk_2_E_in(prog_clk_2_wires[27]),
    .prog_clk_0_N_in(prog_clk_0_wires[145]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[34]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[34]),
    .SC_OUT_TOP(scff_Wires[85]),
    .SC_IN_BOT(scff_Wires[84]),
    .chanx_left_in(sb_1__1__23_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__34_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__34_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__34_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__34_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__34_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__34_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__34_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__34_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__34_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__34_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__34_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__34_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__34_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__34_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__34_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__34_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__34_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__34_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__34_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__34_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__34_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__3_
  (
    .clk_1_S_out(clk_1_wires[55]),
    .clk_1_N_out(clk_1_wires[54]),
    .clk_1_W_in(clk_1_wires[50]),
    .prog_clk_1_S_out(prog_clk_1_wires[55]),
    .prog_clk_1_N_out(prog_clk_1_wires[54]),
    .prog_clk_1_W_in(prog_clk_1_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[148]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[35]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[35]),
    .SC_OUT_TOP(scff_Wires[87]),
    .SC_IN_BOT(scff_Wires[86]),
    .chanx_left_in(sb_1__1__24_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__35_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__35_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__35_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__35_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__35_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__35_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__35_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__35_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__35_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__35_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__35_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__35_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__35_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__35_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__35_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__35_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__35_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__35_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__35_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__35_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__35_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__4_
  (
    .clk_2_W_out(clk_2_wires[37]),
    .clk_2_E_in(clk_2_wires[36]),
    .prog_clk_2_W_out(prog_clk_2_wires[37]),
    .prog_clk_2_E_in(prog_clk_2_wires[36]),
    .prog_clk_0_N_in(prog_clk_0_wires[151]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[36]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[36]),
    .SC_OUT_TOP(scff_Wires[89]),
    .SC_IN_BOT(scff_Wires[88]),
    .chanx_left_in(sb_1__1__25_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__36_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__36_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__36_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__36_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__36_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__36_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__36_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__36_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__36_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__36_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__36_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__36_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__36_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__36_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__36_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__36_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__36_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__36_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__36_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__36_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__36_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__5_
  (
    .clk_1_S_out(clk_1_wires[62]),
    .clk_1_N_out(clk_1_wires[61]),
    .clk_1_W_in(clk_1_wires[57]),
    .prog_clk_1_S_out(prog_clk_1_wires[62]),
    .prog_clk_1_N_out(prog_clk_1_wires[61]),
    .prog_clk_1_W_in(prog_clk_1_wires[57]),
    .prog_clk_0_N_in(prog_clk_0_wires[154]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[37]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[37]),
    .SC_OUT_TOP(scff_Wires[91]),
    .SC_IN_BOT(scff_Wires[90]),
    .chanx_left_in(sb_1__1__26_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__37_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__37_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__37_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__37_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__37_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__37_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__37_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__37_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__37_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__37_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__37_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__37_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__37_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__37_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__37_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__37_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__37_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__37_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__37_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__37_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__37_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__6_
  (
    .clk_3_W_out(clk_3_wires[47]),
    .clk_3_E_in(clk_3_wires[46]),
    .prog_clk_3_W_out(prog_clk_3_wires[47]),
    .prog_clk_3_E_in(prog_clk_3_wires[46]),
    .prog_clk_0_N_in(prog_clk_0_wires[157]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[38]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[38]),
    .SC_OUT_TOP(scff_Wires[93]),
    .SC_IN_BOT(scff_Wires[92]),
    .chanx_left_in(sb_1__1__27_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__38_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__38_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__38_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__38_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__38_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__38_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__38_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__38_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__38_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__38_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__38_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__38_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__38_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__38_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__38_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__38_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__38_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__38_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__38_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__38_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__38_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__7_
  (
    .clk_1_S_out(clk_1_wires[69]),
    .clk_1_N_out(clk_1_wires[68]),
    .clk_1_W_in(clk_1_wires[64]),
    .prog_clk_1_S_out(prog_clk_1_wires[69]),
    .prog_clk_1_N_out(prog_clk_1_wires[68]),
    .prog_clk_1_W_in(prog_clk_1_wires[64]),
    .prog_clk_0_N_in(prog_clk_0_wires[160]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[39]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[39]),
    .SC_OUT_TOP(scff_Wires[95]),
    .SC_IN_BOT(scff_Wires[94]),
    .chanx_left_in(sb_1__1__28_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__39_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__39_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__39_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__39_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__39_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__39_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__39_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__39_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__39_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__39_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__39_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__39_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__39_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__39_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__39_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__39_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__39_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__39_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__39_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__39_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__39_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__8_
  (
    .clk_2_W_out(clk_2_wires[50]),
    .clk_2_E_in(clk_2_wires[49]),
    .prog_clk_2_W_out(prog_clk_2_wires[50]),
    .prog_clk_2_E_in(prog_clk_2_wires[49]),
    .prog_clk_0_N_in(prog_clk_0_wires[163]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[40]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[40]),
    .SC_OUT_TOP(scff_Wires[97]),
    .SC_IN_BOT(scff_Wires[96]),
    .chanx_left_in(sb_1__1__29_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__40_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__40_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__40_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__40_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__40_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__40_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__40_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__40_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__40_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__40_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__40_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__40_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__40_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__40_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__40_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__40_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__40_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__40_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__40_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__40_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__40_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__9_
  (
    .clk_1_S_out(clk_1_wires[76]),
    .clk_1_N_out(clk_1_wires[75]),
    .clk_1_W_in(clk_1_wires[71]),
    .prog_clk_1_S_out(prog_clk_1_wires[76]),
    .prog_clk_1_N_out(prog_clk_1_wires[75]),
    .prog_clk_1_W_in(prog_clk_1_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[166]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[41]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[41]),
    .SC_OUT_TOP(scff_Wires[99]),
    .SC_IN_BOT(scff_Wires[98]),
    .chanx_left_in(sb_1__1__30_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__41_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__41_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__41_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__41_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__41_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__41_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__41_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__41_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__41_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__41_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__41_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__41_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__41_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__41_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__41_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__41_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__41_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__41_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__41_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__41_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__41_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__10_
  (
    .clk_2_W_out(clk_2_wires[63]),
    .clk_2_E_in(clk_2_wires[62]),
    .prog_clk_2_W_out(prog_clk_2_wires[63]),
    .prog_clk_2_E_in(prog_clk_2_wires[62]),
    .prog_clk_0_N_in(prog_clk_0_wires[169]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[42]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[42]),
    .SC_OUT_TOP(scff_Wires[101]),
    .SC_IN_BOT(scff_Wires[100]),
    .chanx_left_in(sb_1__1__31_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__42_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__42_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__42_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__42_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__42_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__42_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__42_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__42_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__42_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__42_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__42_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__42_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__42_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__42_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__42_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__42_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__42_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__42_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__42_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__42_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__42_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__11_
  (
    .clk_1_S_out(clk_1_wires[83]),
    .clk_1_N_out(clk_1_wires[82]),
    .clk_1_W_in(clk_1_wires[78]),
    .prog_clk_1_S_out(prog_clk_1_wires[83]),
    .prog_clk_1_N_out(prog_clk_1_wires[82]),
    .prog_clk_1_W_in(prog_clk_1_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[172]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[43]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[43]),
    .SC_OUT_TOP(scff_Wires[103]),
    .SC_IN_BOT(scff_Wires[102]),
    .chanx_left_in(sb_1__1__32_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__43_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__43_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__43_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__43_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__43_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__43_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__43_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__43_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__43_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__43_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__43_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__43_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__43_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__43_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__43_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__43_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__43_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__43_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__43_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__43_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__43_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__1_
  (
    .clk_1_S_out(clk_1_wires[88]),
    .clk_1_N_out(clk_1_wires[87]),
    .clk_1_E_in(clk_1_wires[86]),
    .prog_clk_1_S_out(prog_clk_1_wires[88]),
    .prog_clk_1_N_out(prog_clk_1_wires[87]),
    .prog_clk_1_E_in(prog_clk_1_wires[86]),
    .prog_clk_0_N_in(prog_clk_0_wires[180]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[44]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[44]),
    .SC_OUT_BOT(scff_Wires[129]),
    .SC_IN_TOP(scff_Wires[128]),
    .chanx_left_in(sb_1__1__33_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__44_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__44_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__44_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__44_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__44_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__44_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__44_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__44_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__44_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__44_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__44_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__44_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__44_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__44_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__44_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__44_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__44_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__44_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__44_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__44_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__44_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__2_
  (
    .clk_2_E_out(clk_2_wires[26]),
    .clk_2_W_in(clk_2_wires[25]),
    .prog_clk_2_E_out(prog_clk_2_wires[26]),
    .prog_clk_2_W_in(prog_clk_2_wires[25]),
    .prog_clk_0_N_in(prog_clk_0_wires[183]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[45]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[45]),
    .SC_OUT_BOT(scff_Wires[127]),
    .SC_IN_TOP(scff_Wires[126]),
    .chanx_left_in(sb_1__1__34_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__45_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__45_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__45_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__45_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__45_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__45_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__45_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__45_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__45_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__45_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__45_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__45_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__45_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__45_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__45_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__45_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__45_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__45_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__45_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__45_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__45_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__3_
  (
    .clk_1_S_out(clk_1_wires[95]),
    .clk_1_N_out(clk_1_wires[94]),
    .clk_1_E_in(clk_1_wires[93]),
    .prog_clk_1_S_out(prog_clk_1_wires[95]),
    .prog_clk_1_N_out(prog_clk_1_wires[94]),
    .prog_clk_1_E_in(prog_clk_1_wires[93]),
    .prog_clk_0_N_in(prog_clk_0_wires[186]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[46]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[46]),
    .SC_OUT_BOT(scff_Wires[125]),
    .SC_IN_TOP(scff_Wires[124]),
    .chanx_left_in(sb_1__1__35_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__46_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__46_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__46_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__46_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__46_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__46_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__46_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__46_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__46_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__46_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__46_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__46_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__46_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__46_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__46_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__46_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__46_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__46_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__46_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__46_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__46_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__4_
  (
    .clk_2_E_out(clk_2_wires[35]),
    .clk_2_W_in(clk_2_wires[34]),
    .prog_clk_2_E_out(prog_clk_2_wires[35]),
    .prog_clk_2_W_in(prog_clk_2_wires[34]),
    .prog_clk_0_N_in(prog_clk_0_wires[189]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[47]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[47]),
    .SC_OUT_BOT(scff_Wires[123]),
    .SC_IN_TOP(scff_Wires[122]),
    .chanx_left_in(sb_1__1__36_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__47_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__47_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__47_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__47_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__47_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__47_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__47_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__47_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__47_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__47_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__47_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__47_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__47_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__47_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__47_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__47_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__47_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__47_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__47_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__47_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__47_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__5_
  (
    .clk_1_S_out(clk_1_wires[102]),
    .clk_1_N_out(clk_1_wires[101]),
    .clk_1_E_in(clk_1_wires[100]),
    .prog_clk_1_S_out(prog_clk_1_wires[102]),
    .prog_clk_1_N_out(prog_clk_1_wires[101]),
    .prog_clk_1_E_in(prog_clk_1_wires[100]),
    .prog_clk_0_N_in(prog_clk_0_wires[192]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[48]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[48]),
    .SC_OUT_BOT(scff_Wires[121]),
    .SC_IN_TOP(scff_Wires[120]),
    .chanx_left_in(sb_1__1__37_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__48_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__48_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__48_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__48_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__48_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__48_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__48_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__48_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__48_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__48_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__48_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__48_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__48_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__48_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__48_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__48_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__48_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__48_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__48_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__48_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__48_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__6_
  (
    .clk_3_W_out(clk_3_wires[7]),
    .clk_3_E_in(clk_3_wires[6]),
    .prog_clk_3_W_out(prog_clk_3_wires[7]),
    .prog_clk_3_E_in(prog_clk_3_wires[6]),
    .prog_clk_0_N_in(prog_clk_0_wires[195]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[49]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[49]),
    .SC_OUT_BOT(scff_Wires[119]),
    .SC_IN_TOP(scff_Wires[118]),
    .chanx_left_in(sb_1__1__38_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__49_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__49_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__49_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__49_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__49_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__49_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__49_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__49_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__49_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__49_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__49_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__49_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__49_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__49_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__49_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__49_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__49_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__49_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__49_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__49_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__49_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__7_
  (
    .clk_1_S_out(clk_1_wires[109]),
    .clk_1_N_out(clk_1_wires[108]),
    .clk_1_E_in(clk_1_wires[107]),
    .prog_clk_1_S_out(prog_clk_1_wires[109]),
    .prog_clk_1_N_out(prog_clk_1_wires[108]),
    .prog_clk_1_E_in(prog_clk_1_wires[107]),
    .prog_clk_0_N_in(prog_clk_0_wires[198]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[50]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[50]),
    .SC_OUT_BOT(scff_Wires[117]),
    .SC_IN_TOP(scff_Wires[116]),
    .chanx_left_in(sb_1__1__39_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__50_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__50_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__50_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__50_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__50_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__50_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__50_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__50_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__50_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__50_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__50_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__50_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__50_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__50_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__50_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__50_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__50_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__50_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__50_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__50_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__50_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__8_
  (
    .clk_2_E_out(clk_2_wires[48]),
    .clk_2_W_in(clk_2_wires[47]),
    .prog_clk_2_E_out(prog_clk_2_wires[48]),
    .prog_clk_2_W_in(prog_clk_2_wires[47]),
    .prog_clk_0_N_in(prog_clk_0_wires[201]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[51]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[51]),
    .SC_OUT_BOT(scff_Wires[115]),
    .SC_IN_TOP(scff_Wires[114]),
    .chanx_left_in(sb_1__1__40_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__51_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__51_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__51_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__51_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__51_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__51_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__51_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__51_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__51_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__51_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__51_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__51_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__51_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__51_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__51_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__51_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__51_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__51_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__51_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__51_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__51_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__9_
  (
    .clk_1_S_out(clk_1_wires[116]),
    .clk_1_N_out(clk_1_wires[115]),
    .clk_1_E_in(clk_1_wires[114]),
    .prog_clk_1_S_out(prog_clk_1_wires[116]),
    .prog_clk_1_N_out(prog_clk_1_wires[115]),
    .prog_clk_1_E_in(prog_clk_1_wires[114]),
    .prog_clk_0_N_in(prog_clk_0_wires[204]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[52]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[52]),
    .SC_OUT_BOT(scff_Wires[113]),
    .SC_IN_TOP(scff_Wires[112]),
    .chanx_left_in(sb_1__1__41_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__52_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__52_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__52_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__52_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__52_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__52_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__52_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__52_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__52_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__52_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__52_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__52_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__52_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__52_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__52_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__52_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__52_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__52_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__52_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__52_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__52_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__10_
  (
    .clk_2_E_out(clk_2_wires[61]),
    .clk_2_W_in(clk_2_wires[60]),
    .prog_clk_2_E_out(prog_clk_2_wires[61]),
    .prog_clk_2_W_in(prog_clk_2_wires[60]),
    .prog_clk_0_N_in(prog_clk_0_wires[207]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[53]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[53]),
    .SC_OUT_BOT(scff_Wires[111]),
    .SC_IN_TOP(scff_Wires[110]),
    .chanx_left_in(sb_1__1__42_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__53_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__53_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__53_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__53_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__53_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__53_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__53_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__53_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__53_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__53_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__53_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__53_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__53_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__53_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__53_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__53_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__53_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__53_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__53_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__53_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__53_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__11_
  (
    .clk_1_S_out(clk_1_wires[123]),
    .clk_1_N_out(clk_1_wires[122]),
    .clk_1_E_in(clk_1_wires[121]),
    .prog_clk_1_S_out(prog_clk_1_wires[123]),
    .prog_clk_1_N_out(prog_clk_1_wires[122]),
    .prog_clk_1_E_in(prog_clk_1_wires[121]),
    .prog_clk_0_N_in(prog_clk_0_wires[210]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[54]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[54]),
    .SC_OUT_BOT(scff_Wires[109]),
    .SC_IN_TOP(scff_Wires[108]),
    .chanx_left_in(sb_1__1__43_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__54_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__54_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__54_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__54_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__54_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__54_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__54_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__54_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__54_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__54_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__54_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__54_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__54_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__54_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__54_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__54_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__54_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__54_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__54_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__54_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__54_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__1_
  (
    .clk_1_S_out(clk_1_wires[90]),
    .clk_1_N_out(clk_1_wires[89]),
    .clk_1_W_in(clk_1_wires[85]),
    .prog_clk_1_S_out(prog_clk_1_wires[90]),
    .prog_clk_1_N_out(prog_clk_1_wires[89]),
    .prog_clk_1_W_in(prog_clk_1_wires[85]),
    .prog_clk_0_N_in(prog_clk_0_wires[218]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[55]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[55]),
    .SC_OUT_TOP(scff_Wires[136]),
    .SC_IN_BOT(scff_Wires[135]),
    .chanx_left_in(sb_1__1__44_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__55_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__55_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__55_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__55_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__55_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__55_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__55_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__55_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__55_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__55_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__55_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__55_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__55_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__55_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__55_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__55_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__55_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__55_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__55_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__55_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__55_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[221]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[56]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[56]),
    .SC_OUT_TOP(scff_Wires[138]),
    .SC_IN_BOT(scff_Wires[137]),
    .chanx_left_in(sb_1__1__45_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__56_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__56_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__56_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__56_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__56_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__56_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__56_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__56_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__56_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__56_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__56_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__56_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__56_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__56_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__56_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__56_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__56_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__56_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__56_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__56_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__56_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__3_
  (
    .clk_1_S_out(clk_1_wires[97]),
    .clk_1_N_out(clk_1_wires[96]),
    .clk_1_W_in(clk_1_wires[92]),
    .prog_clk_1_S_out(prog_clk_1_wires[97]),
    .prog_clk_1_N_out(prog_clk_1_wires[96]),
    .prog_clk_1_W_in(prog_clk_1_wires[92]),
    .prog_clk_0_N_in(prog_clk_0_wires[224]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[57]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[57]),
    .SC_OUT_TOP(scff_Wires[140]),
    .SC_IN_BOT(scff_Wires[139]),
    .chanx_left_in(sb_1__1__46_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__57_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__57_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__57_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__57_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__57_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__57_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__57_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__57_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__57_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__57_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__57_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__57_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__57_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__57_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__57_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__57_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__57_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__57_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__57_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__57_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__57_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[227]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[58]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[58]),
    .SC_OUT_TOP(scff_Wires[142]),
    .SC_IN_BOT(scff_Wires[141]),
    .chanx_left_in(sb_1__1__47_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__58_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__58_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__58_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__58_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__58_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__58_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__58_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__58_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__58_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__58_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__58_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__58_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__58_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__58_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__58_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__58_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__58_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__58_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__58_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__58_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__58_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__5_
  (
    .clk_1_S_out(clk_1_wires[104]),
    .clk_1_N_out(clk_1_wires[103]),
    .clk_1_W_in(clk_1_wires[99]),
    .prog_clk_1_S_out(prog_clk_1_wires[104]),
    .prog_clk_1_N_out(prog_clk_1_wires[103]),
    .prog_clk_1_W_in(prog_clk_1_wires[99]),
    .prog_clk_0_N_in(prog_clk_0_wires[230]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[59]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[59]),
    .SC_OUT_TOP(scff_Wires[144]),
    .SC_IN_BOT(scff_Wires[143]),
    .chanx_left_in(sb_1__1__48_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__59_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__59_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__59_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__59_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__59_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__59_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__59_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__59_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__59_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__59_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__59_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__59_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__59_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__59_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__59_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__59_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__59_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__59_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__59_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__59_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__59_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__6_
  (
    .clk_3_W_out(clk_3_wires[3]),
    .clk_3_E_in(clk_3_wires[2]),
    .prog_clk_3_W_out(prog_clk_3_wires[3]),
    .prog_clk_3_E_in(prog_clk_3_wires[2]),
    .prog_clk_0_N_in(prog_clk_0_wires[233]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[60]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[60]),
    .SC_OUT_TOP(scff_Wires[146]),
    .SC_IN_BOT(scff_Wires[145]),
    .chanx_left_in(sb_1__1__49_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__60_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__60_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__60_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__60_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__60_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__60_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__60_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__60_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__60_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__60_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__60_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__60_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__60_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__60_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__60_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__60_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__60_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__60_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__60_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__60_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__60_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__7_
  (
    .clk_1_S_out(clk_1_wires[111]),
    .clk_1_N_out(clk_1_wires[110]),
    .clk_1_W_in(clk_1_wires[106]),
    .prog_clk_1_S_out(prog_clk_1_wires[111]),
    .prog_clk_1_N_out(prog_clk_1_wires[110]),
    .prog_clk_1_W_in(prog_clk_1_wires[106]),
    .prog_clk_0_N_in(prog_clk_0_wires[236]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[61]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[61]),
    .SC_OUT_TOP(scff_Wires[148]),
    .SC_IN_BOT(scff_Wires[147]),
    .chanx_left_in(sb_1__1__50_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__61_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__61_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__61_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__61_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__61_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__61_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__61_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__61_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__61_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__61_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__61_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__61_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__61_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__61_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__61_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__61_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__61_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__61_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__61_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__61_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__61_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[239]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[62]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[62]),
    .SC_OUT_TOP(scff_Wires[150]),
    .SC_IN_BOT(scff_Wires[149]),
    .chanx_left_in(sb_1__1__51_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__62_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__62_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__62_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__62_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__62_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__62_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__62_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__62_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__62_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__62_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__62_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__62_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__62_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__62_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__62_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__62_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__62_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__62_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__62_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__62_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__62_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__9_
  (
    .clk_1_S_out(clk_1_wires[118]),
    .clk_1_N_out(clk_1_wires[117]),
    .clk_1_W_in(clk_1_wires[113]),
    .prog_clk_1_S_out(prog_clk_1_wires[118]),
    .prog_clk_1_N_out(prog_clk_1_wires[117]),
    .prog_clk_1_W_in(prog_clk_1_wires[113]),
    .prog_clk_0_N_in(prog_clk_0_wires[242]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[63]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[63]),
    .SC_OUT_TOP(scff_Wires[152]),
    .SC_IN_BOT(scff_Wires[151]),
    .chanx_left_in(sb_1__1__52_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__63_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__63_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__63_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__63_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__63_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__63_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__63_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__63_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__63_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__63_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__63_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__63_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__63_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__63_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__63_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__63_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__63_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__63_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__63_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__63_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__63_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[245]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[64]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[64]),
    .SC_OUT_TOP(scff_Wires[154]),
    .SC_IN_BOT(scff_Wires[153]),
    .chanx_left_in(sb_1__1__53_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__64_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__64_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__64_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__64_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__64_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__64_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__64_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__64_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__64_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__64_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__64_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__64_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__64_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__64_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__64_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__64_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__64_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__64_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__64_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__64_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__64_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__11_
  (
    .clk_1_S_out(clk_1_wires[125]),
    .clk_1_N_out(clk_1_wires[124]),
    .clk_1_W_in(clk_1_wires[120]),
    .prog_clk_1_S_out(prog_clk_1_wires[125]),
    .prog_clk_1_N_out(prog_clk_1_wires[124]),
    .prog_clk_1_W_in(prog_clk_1_wires[120]),
    .prog_clk_0_N_in(prog_clk_0_wires[248]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[65]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[65]),
    .SC_OUT_TOP(scff_Wires[156]),
    .SC_IN_BOT(scff_Wires[155]),
    .chanx_left_in(sb_1__1__54_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__65_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__65_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__65_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__65_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__65_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__65_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__65_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__65_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__65_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__65_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__65_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__65_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__65_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__65_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__65_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__65_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__65_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__65_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__65_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__65_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__65_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__1_
  (
    .clk_1_S_out(clk_1_wires[130]),
    .clk_1_N_out(clk_1_wires[129]),
    .clk_1_E_in(clk_1_wires[128]),
    .prog_clk_1_S_out(prog_clk_1_wires[130]),
    .prog_clk_1_N_out(prog_clk_1_wires[129]),
    .prog_clk_1_E_in(prog_clk_1_wires[128]),
    .prog_clk_0_N_in(prog_clk_0_wires[256]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[66]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[66]),
    .SC_OUT_BOT(scff_Wires[182]),
    .SC_IN_TOP(scff_Wires[181]),
    .chanx_left_in(sb_1__1__55_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__66_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__66_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__66_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__66_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__66_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__66_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__66_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__66_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__66_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__66_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__66_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__66_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__66_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__66_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__66_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__66_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__66_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__66_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__66_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__66_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__66_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[259]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[67]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[67]),
    .SC_OUT_BOT(scff_Wires[180]),
    .SC_IN_TOP(scff_Wires[179]),
    .chanx_left_in(sb_1__1__56_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__67_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__67_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__67_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__67_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__67_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__67_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__67_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__67_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__67_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__67_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__67_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__67_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__67_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__67_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__67_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__67_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__67_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__67_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__67_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__67_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__67_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__3_
  (
    .clk_1_S_out(clk_1_wires[137]),
    .clk_1_N_out(clk_1_wires[136]),
    .clk_1_E_in(clk_1_wires[135]),
    .prog_clk_1_S_out(prog_clk_1_wires[137]),
    .prog_clk_1_N_out(prog_clk_1_wires[136]),
    .prog_clk_1_E_in(prog_clk_1_wires[135]),
    .prog_clk_0_N_in(prog_clk_0_wires[262]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[68]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[68]),
    .SC_OUT_BOT(scff_Wires[178]),
    .SC_IN_TOP(scff_Wires[177]),
    .chanx_left_in(sb_1__1__57_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__68_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__68_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__68_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__68_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__68_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__68_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__68_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__68_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__68_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__68_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__68_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__68_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__68_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__68_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__68_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__68_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__68_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__68_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__68_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__68_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__68_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[265]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[69]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[69]),
    .SC_OUT_BOT(scff_Wires[176]),
    .SC_IN_TOP(scff_Wires[175]),
    .chanx_left_in(sb_1__1__58_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__69_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__69_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__69_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__69_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__69_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__69_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__69_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__69_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__69_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__69_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__69_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__69_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__69_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__69_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__69_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__69_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__69_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__69_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__69_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__69_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__69_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__5_
  (
    .clk_1_S_out(clk_1_wires[144]),
    .clk_1_N_out(clk_1_wires[143]),
    .clk_1_E_in(clk_1_wires[142]),
    .prog_clk_1_S_out(prog_clk_1_wires[144]),
    .prog_clk_1_N_out(prog_clk_1_wires[143]),
    .prog_clk_1_E_in(prog_clk_1_wires[142]),
    .prog_clk_0_N_in(prog_clk_0_wires[268]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[70]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[70]),
    .SC_OUT_BOT(scff_Wires[174]),
    .SC_IN_TOP(scff_Wires[173]),
    .chanx_left_in(sb_1__1__59_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__70_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__70_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__70_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__70_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__70_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__70_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__70_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__70_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__70_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__70_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__70_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__70_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__70_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__70_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__70_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__70_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__70_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__70_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__70_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__70_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__70_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__6_
  (
    .clk_3_E_out(clk_3_wires[1]),
    .clk_3_W_in(clk_3_wires[0]),
    .prog_clk_3_E_out(prog_clk_3_wires[1]),
    .prog_clk_3_W_in(prog_clk_3_wires[0]),
    .prog_clk_0_N_in(prog_clk_0_wires[271]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[71]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[71]),
    .SC_OUT_BOT(scff_Wires[172]),
    .SC_IN_TOP(scff_Wires[171]),
    .chanx_left_in(sb_1__1__60_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__71_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__71_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__71_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__71_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__71_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__71_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__71_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__71_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__71_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__71_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__71_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__71_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__71_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__71_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__71_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__71_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__71_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__71_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__71_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__71_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__71_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__7_
  (
    .clk_1_S_out(clk_1_wires[151]),
    .clk_1_N_out(clk_1_wires[150]),
    .clk_1_E_in(clk_1_wires[149]),
    .prog_clk_1_S_out(prog_clk_1_wires[151]),
    .prog_clk_1_N_out(prog_clk_1_wires[150]),
    .prog_clk_1_E_in(prog_clk_1_wires[149]),
    .prog_clk_0_N_in(prog_clk_0_wires[274]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[72]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[72]),
    .SC_OUT_BOT(scff_Wires[170]),
    .SC_IN_TOP(scff_Wires[169]),
    .chanx_left_in(sb_1__1__61_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__72_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__72_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__72_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__72_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__72_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__72_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__72_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__72_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__72_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__72_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__72_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__72_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__72_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__72_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__72_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__72_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__72_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__72_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__72_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__72_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__72_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[277]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[73]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[73]),
    .SC_OUT_BOT(scff_Wires[168]),
    .SC_IN_TOP(scff_Wires[167]),
    .chanx_left_in(sb_1__1__62_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__73_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__73_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__73_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__73_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__73_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__73_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__73_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__73_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__73_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__73_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__73_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__73_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__73_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__73_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__73_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__73_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__73_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__73_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__73_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__73_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__73_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__9_
  (
    .clk_1_S_out(clk_1_wires[158]),
    .clk_1_N_out(clk_1_wires[157]),
    .clk_1_E_in(clk_1_wires[156]),
    .prog_clk_1_S_out(prog_clk_1_wires[158]),
    .prog_clk_1_N_out(prog_clk_1_wires[157]),
    .prog_clk_1_E_in(prog_clk_1_wires[156]),
    .prog_clk_0_N_in(prog_clk_0_wires[280]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[74]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[74]),
    .SC_OUT_BOT(scff_Wires[166]),
    .SC_IN_TOP(scff_Wires[165]),
    .chanx_left_in(sb_1__1__63_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__74_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__74_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__74_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__74_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__74_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__74_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__74_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__74_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__74_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__74_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__74_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__74_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__74_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__74_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__74_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__74_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__74_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__74_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__74_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__74_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__74_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[283]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[75]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[75]),
    .SC_OUT_BOT(scff_Wires[164]),
    .SC_IN_TOP(scff_Wires[163]),
    .chanx_left_in(sb_1__1__64_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__75_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__75_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__75_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__75_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__75_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__75_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__75_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__75_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__75_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__75_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__75_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__75_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__75_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__75_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__75_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__75_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__75_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__75_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__75_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__75_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__75_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__11_
  (
    .clk_1_S_out(clk_1_wires[165]),
    .clk_1_N_out(clk_1_wires[164]),
    .clk_1_E_in(clk_1_wires[163]),
    .prog_clk_1_S_out(prog_clk_1_wires[165]),
    .prog_clk_1_N_out(prog_clk_1_wires[164]),
    .prog_clk_1_E_in(prog_clk_1_wires[163]),
    .prog_clk_0_N_in(prog_clk_0_wires[286]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[76]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[76]),
    .SC_OUT_BOT(scff_Wires[162]),
    .SC_IN_TOP(scff_Wires[161]),
    .chanx_left_in(sb_1__1__65_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__76_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__76_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__76_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__76_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__76_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__76_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__76_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__76_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__76_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__76_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__76_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__76_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__76_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__76_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__76_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__76_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__76_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__76_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__76_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__76_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__76_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__1_
  (
    .clk_1_S_out(clk_1_wires[132]),
    .clk_1_N_out(clk_1_wires[131]),
    .clk_1_W_in(clk_1_wires[127]),
    .prog_clk_1_S_out(prog_clk_1_wires[132]),
    .prog_clk_1_N_out(prog_clk_1_wires[131]),
    .prog_clk_1_W_in(prog_clk_1_wires[127]),
    .prog_clk_0_N_in(prog_clk_0_wires[294]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[77]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[77]),
    .SC_OUT_TOP(scff_Wires[189]),
    .SC_IN_BOT(scff_Wires[188]),
    .chanx_left_in(sb_1__1__66_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__77_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__77_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__77_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__77_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__77_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__77_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__77_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__77_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__77_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__77_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__77_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__77_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__77_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__77_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__77_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__77_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__77_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__77_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__77_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__77_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__77_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__2_
  (
    .clk_2_W_out(clk_2_wires[72]),
    .clk_2_E_in(clk_2_wires[71]),
    .prog_clk_2_W_out(prog_clk_2_wires[72]),
    .prog_clk_2_E_in(prog_clk_2_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[297]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[78]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[78]),
    .SC_OUT_TOP(scff_Wires[191]),
    .SC_IN_BOT(scff_Wires[190]),
    .chanx_left_in(sb_1__1__67_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__78_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__78_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__78_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__78_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__78_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__78_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__78_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__78_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__78_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__78_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__78_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__78_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__78_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__78_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__78_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__78_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__78_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__78_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__78_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__78_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__78_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__3_
  (
    .clk_1_S_out(clk_1_wires[139]),
    .clk_1_N_out(clk_1_wires[138]),
    .clk_1_W_in(clk_1_wires[134]),
    .prog_clk_1_S_out(prog_clk_1_wires[139]),
    .prog_clk_1_N_out(prog_clk_1_wires[138]),
    .prog_clk_1_W_in(prog_clk_1_wires[134]),
    .prog_clk_0_N_in(prog_clk_0_wires[300]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[79]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[79]),
    .SC_OUT_TOP(scff_Wires[193]),
    .SC_IN_BOT(scff_Wires[192]),
    .chanx_left_in(sb_1__1__68_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__79_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__79_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__79_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__79_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__79_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__79_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__79_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__79_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__79_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__79_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__79_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__79_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__79_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__79_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__79_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__79_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__79_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__79_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__79_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__79_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__79_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__4_
  (
    .clk_2_W_out(clk_2_wires[81]),
    .clk_2_E_in(clk_2_wires[80]),
    .prog_clk_2_W_out(prog_clk_2_wires[81]),
    .prog_clk_2_E_in(prog_clk_2_wires[80]),
    .prog_clk_0_N_in(prog_clk_0_wires[303]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[80]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[80]),
    .SC_OUT_TOP(scff_Wires[195]),
    .SC_IN_BOT(scff_Wires[194]),
    .chanx_left_in(sb_1__1__69_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__80_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__80_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__80_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__80_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__80_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__80_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__80_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__80_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__80_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__80_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__80_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__80_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__80_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__80_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__80_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__80_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__80_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__80_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__80_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__80_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__80_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__5_
  (
    .clk_1_S_out(clk_1_wires[146]),
    .clk_1_N_out(clk_1_wires[145]),
    .clk_1_W_in(clk_1_wires[141]),
    .prog_clk_1_S_out(prog_clk_1_wires[146]),
    .prog_clk_1_N_out(prog_clk_1_wires[145]),
    .prog_clk_1_W_in(prog_clk_1_wires[141]),
    .prog_clk_0_N_in(prog_clk_0_wires[306]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[81]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[81]),
    .SC_OUT_TOP(scff_Wires[197]),
    .SC_IN_BOT(scff_Wires[196]),
    .chanx_left_in(sb_1__1__70_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__81_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__81_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__81_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__81_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__81_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__81_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__81_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__81_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__81_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__81_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__81_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__81_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__81_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__81_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__81_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__81_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__81_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__81_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__81_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__81_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__81_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__6_
  (
    .clk_3_E_out(clk_3_wires[5]),
    .clk_3_W_in(clk_3_wires[4]),
    .prog_clk_3_E_out(prog_clk_3_wires[5]),
    .prog_clk_3_W_in(prog_clk_3_wires[4]),
    .prog_clk_0_N_in(prog_clk_0_wires[309]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[82]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[82]),
    .SC_OUT_TOP(scff_Wires[199]),
    .SC_IN_BOT(scff_Wires[198]),
    .chanx_left_in(sb_1__1__71_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__82_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__82_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__82_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__82_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__82_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__82_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__82_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__82_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__82_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__82_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__82_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__82_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__82_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__82_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__82_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__82_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__82_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__82_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__82_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__82_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__82_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__7_
  (
    .clk_1_S_out(clk_1_wires[153]),
    .clk_1_N_out(clk_1_wires[152]),
    .clk_1_W_in(clk_1_wires[148]),
    .prog_clk_1_S_out(prog_clk_1_wires[153]),
    .prog_clk_1_N_out(prog_clk_1_wires[152]),
    .prog_clk_1_W_in(prog_clk_1_wires[148]),
    .prog_clk_0_N_in(prog_clk_0_wires[312]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[83]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[83]),
    .SC_OUT_TOP(scff_Wires[201]),
    .SC_IN_BOT(scff_Wires[200]),
    .chanx_left_in(sb_1__1__72_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__83_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__83_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__83_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__83_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__83_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__83_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__83_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__83_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__83_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__83_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__83_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__83_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__83_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__83_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__83_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__83_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__83_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__83_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__83_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__83_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__83_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__8_
  (
    .clk_2_W_out(clk_2_wires[94]),
    .clk_2_E_in(clk_2_wires[93]),
    .prog_clk_2_W_out(prog_clk_2_wires[94]),
    .prog_clk_2_E_in(prog_clk_2_wires[93]),
    .prog_clk_0_N_in(prog_clk_0_wires[315]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[84]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[84]),
    .SC_OUT_TOP(scff_Wires[203]),
    .SC_IN_BOT(scff_Wires[202]),
    .chanx_left_in(sb_1__1__73_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__84_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__84_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__84_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__84_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__84_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__84_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__84_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__84_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__84_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__84_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__84_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__84_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__84_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__84_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__84_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__84_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__84_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__84_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__84_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__84_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__84_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__9_
  (
    .clk_1_S_out(clk_1_wires[160]),
    .clk_1_N_out(clk_1_wires[159]),
    .clk_1_W_in(clk_1_wires[155]),
    .prog_clk_1_S_out(prog_clk_1_wires[160]),
    .prog_clk_1_N_out(prog_clk_1_wires[159]),
    .prog_clk_1_W_in(prog_clk_1_wires[155]),
    .prog_clk_0_N_in(prog_clk_0_wires[318]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[85]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[85]),
    .SC_OUT_TOP(scff_Wires[205]),
    .SC_IN_BOT(scff_Wires[204]),
    .chanx_left_in(sb_1__1__74_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__85_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__85_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__85_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__85_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__85_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__85_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__85_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__85_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__85_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__85_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__85_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__85_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__85_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__85_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__85_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__85_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__85_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__85_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__85_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__85_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__85_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__10_
  (
    .clk_2_W_out(clk_2_wires[107]),
    .clk_2_E_in(clk_2_wires[106]),
    .prog_clk_2_W_out(prog_clk_2_wires[107]),
    .prog_clk_2_E_in(prog_clk_2_wires[106]),
    .prog_clk_0_N_in(prog_clk_0_wires[321]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[86]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[86]),
    .SC_OUT_TOP(scff_Wires[207]),
    .SC_IN_BOT(scff_Wires[206]),
    .chanx_left_in(sb_1__1__75_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__86_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__86_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__86_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__86_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__86_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__86_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__86_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__86_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__86_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__86_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__86_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__86_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__86_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__86_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__86_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__86_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__86_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__86_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__86_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__86_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__86_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__11_
  (
    .clk_1_S_out(clk_1_wires[167]),
    .clk_1_N_out(clk_1_wires[166]),
    .clk_1_W_in(clk_1_wires[162]),
    .prog_clk_1_S_out(prog_clk_1_wires[167]),
    .prog_clk_1_N_out(prog_clk_1_wires[166]),
    .prog_clk_1_W_in(prog_clk_1_wires[162]),
    .prog_clk_0_N_in(prog_clk_0_wires[324]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[87]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[87]),
    .SC_OUT_TOP(scff_Wires[209]),
    .SC_IN_BOT(scff_Wires[208]),
    .chanx_left_in(sb_1__1__76_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__87_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__87_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__87_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__87_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__87_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__87_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__87_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__87_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__87_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__87_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__87_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__87_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__87_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__87_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__87_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__87_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__87_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__87_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__87_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__87_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__87_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__1_
  (
    .clk_1_S_out(clk_1_wires[172]),
    .clk_1_N_out(clk_1_wires[171]),
    .clk_1_E_in(clk_1_wires[170]),
    .prog_clk_1_S_out(prog_clk_1_wires[172]),
    .prog_clk_1_N_out(prog_clk_1_wires[171]),
    .prog_clk_1_E_in(prog_clk_1_wires[170]),
    .prog_clk_0_N_in(prog_clk_0_wires[332]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[88]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[88]),
    .SC_OUT_BOT(scff_Wires[235]),
    .SC_IN_TOP(scff_Wires[234]),
    .chanx_left_in(sb_1__1__77_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__88_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__88_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__88_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__88_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__88_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__88_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__88_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__88_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__88_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__88_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__88_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__88_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__88_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__88_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__88_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__88_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__88_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__88_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__88_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__88_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__88_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__2_
  (
    .clk_2_E_out(clk_2_wires[70]),
    .clk_2_W_in(clk_2_wires[69]),
    .prog_clk_2_E_out(prog_clk_2_wires[70]),
    .prog_clk_2_W_in(prog_clk_2_wires[69]),
    .prog_clk_0_N_in(prog_clk_0_wires[335]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[89]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[89]),
    .SC_OUT_BOT(scff_Wires[233]),
    .SC_IN_TOP(scff_Wires[232]),
    .chanx_left_in(sb_1__1__78_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__89_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__89_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__89_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__89_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__89_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__89_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__89_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__89_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__89_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__89_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__89_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__89_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__89_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__89_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__89_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__89_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__89_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__89_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__89_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__89_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__89_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__3_
  (
    .clk_1_S_out(clk_1_wires[179]),
    .clk_1_N_out(clk_1_wires[178]),
    .clk_1_E_in(clk_1_wires[177]),
    .prog_clk_1_S_out(prog_clk_1_wires[179]),
    .prog_clk_1_N_out(prog_clk_1_wires[178]),
    .prog_clk_1_E_in(prog_clk_1_wires[177]),
    .prog_clk_0_N_in(prog_clk_0_wires[338]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[90]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[90]),
    .SC_OUT_BOT(scff_Wires[231]),
    .SC_IN_TOP(scff_Wires[230]),
    .chanx_left_in(sb_1__1__79_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__90_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__90_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__90_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__90_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__90_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__90_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__90_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__90_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__90_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__90_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__90_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__90_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__90_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__90_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__90_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__90_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__90_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__90_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__90_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__90_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__90_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__4_
  (
    .clk_2_E_out(clk_2_wires[79]),
    .clk_2_W_in(clk_2_wires[78]),
    .prog_clk_2_E_out(prog_clk_2_wires[79]),
    .prog_clk_2_W_in(prog_clk_2_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[341]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[91]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[91]),
    .SC_OUT_BOT(scff_Wires[229]),
    .SC_IN_TOP(scff_Wires[228]),
    .chanx_left_in(sb_1__1__80_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__91_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__91_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__91_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__91_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__91_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__91_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__91_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__91_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__91_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__91_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__91_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__91_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__91_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__91_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__91_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__91_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__91_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__91_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__91_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__91_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__91_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__5_
  (
    .clk_1_S_out(clk_1_wires[186]),
    .clk_1_N_out(clk_1_wires[185]),
    .clk_1_E_in(clk_1_wires[184]),
    .prog_clk_1_S_out(prog_clk_1_wires[186]),
    .prog_clk_1_N_out(prog_clk_1_wires[185]),
    .prog_clk_1_E_in(prog_clk_1_wires[184]),
    .prog_clk_0_N_in(prog_clk_0_wires[344]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[92]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[92]),
    .SC_OUT_BOT(scff_Wires[227]),
    .SC_IN_TOP(scff_Wires[226]),
    .chanx_left_in(sb_1__1__81_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__92_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__92_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__92_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__92_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__92_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__92_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__92_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__92_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__92_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__92_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__92_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__92_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__92_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__92_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__92_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__92_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__92_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__92_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__92_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__92_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__92_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__6_
  (
    .clk_3_E_out(clk_3_wires[45]),
    .clk_3_W_in(clk_3_wires[44]),
    .prog_clk_3_E_out(prog_clk_3_wires[45]),
    .prog_clk_3_W_in(prog_clk_3_wires[44]),
    .prog_clk_0_N_in(prog_clk_0_wires[347]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[93]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[93]),
    .SC_OUT_BOT(scff_Wires[225]),
    .SC_IN_TOP(scff_Wires[224]),
    .chanx_left_in(sb_1__1__82_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__93_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__93_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__93_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__93_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__93_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__93_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__93_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__93_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__93_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__93_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__93_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__93_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__93_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__93_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__93_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__93_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__93_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__93_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__93_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__93_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__93_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__7_
  (
    .clk_1_S_out(clk_1_wires[193]),
    .clk_1_N_out(clk_1_wires[192]),
    .clk_1_E_in(clk_1_wires[191]),
    .prog_clk_1_S_out(prog_clk_1_wires[193]),
    .prog_clk_1_N_out(prog_clk_1_wires[192]),
    .prog_clk_1_E_in(prog_clk_1_wires[191]),
    .prog_clk_0_N_in(prog_clk_0_wires[350]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[94]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[94]),
    .SC_OUT_BOT(scff_Wires[223]),
    .SC_IN_TOP(scff_Wires[222]),
    .chanx_left_in(sb_1__1__83_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__94_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__94_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__94_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__94_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__94_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__94_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__94_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__94_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__94_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__94_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__94_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__94_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__94_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__94_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__94_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__94_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__94_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__94_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__94_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__94_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__94_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__8_
  (
    .clk_2_E_out(clk_2_wires[92]),
    .clk_2_W_in(clk_2_wires[91]),
    .prog_clk_2_E_out(prog_clk_2_wires[92]),
    .prog_clk_2_W_in(prog_clk_2_wires[91]),
    .prog_clk_0_N_in(prog_clk_0_wires[353]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[95]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[95]),
    .SC_OUT_BOT(scff_Wires[221]),
    .SC_IN_TOP(scff_Wires[220]),
    .chanx_left_in(sb_1__1__84_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__95_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__95_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__95_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__95_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__95_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__95_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__95_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__95_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__95_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__95_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__95_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__95_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__95_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__95_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__95_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__95_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__95_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__95_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__95_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__95_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__95_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__9_
  (
    .clk_1_S_out(clk_1_wires[200]),
    .clk_1_N_out(clk_1_wires[199]),
    .clk_1_E_in(clk_1_wires[198]),
    .prog_clk_1_S_out(prog_clk_1_wires[200]),
    .prog_clk_1_N_out(prog_clk_1_wires[199]),
    .prog_clk_1_E_in(prog_clk_1_wires[198]),
    .prog_clk_0_N_in(prog_clk_0_wires[356]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[96]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[96]),
    .SC_OUT_BOT(scff_Wires[219]),
    .SC_IN_TOP(scff_Wires[218]),
    .chanx_left_in(sb_1__1__85_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__96_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__96_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__96_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__96_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__96_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__96_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__96_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__96_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__96_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__96_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__96_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__96_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__96_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__96_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__96_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__96_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__96_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__96_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__96_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__96_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__96_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__10_
  (
    .clk_2_E_out(clk_2_wires[105]),
    .clk_2_W_in(clk_2_wires[104]),
    .prog_clk_2_E_out(prog_clk_2_wires[105]),
    .prog_clk_2_W_in(prog_clk_2_wires[104]),
    .prog_clk_0_N_in(prog_clk_0_wires[359]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[97]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[97]),
    .SC_OUT_BOT(scff_Wires[217]),
    .SC_IN_TOP(scff_Wires[216]),
    .chanx_left_in(sb_1__1__86_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__97_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__97_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__97_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__97_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__97_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__97_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__97_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__97_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__97_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__97_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__97_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__97_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__97_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__97_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__97_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__97_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__97_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__97_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__97_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__97_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__97_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__11_
  (
    .clk_1_S_out(clk_1_wires[207]),
    .clk_1_N_out(clk_1_wires[206]),
    .clk_1_E_in(clk_1_wires[205]),
    .prog_clk_1_S_out(prog_clk_1_wires[207]),
    .prog_clk_1_N_out(prog_clk_1_wires[206]),
    .prog_clk_1_E_in(prog_clk_1_wires[205]),
    .prog_clk_0_N_in(prog_clk_0_wires[362]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[98]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[98]),
    .SC_OUT_BOT(scff_Wires[215]),
    .SC_IN_TOP(scff_Wires[214]),
    .chanx_left_in(sb_1__1__87_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__98_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__98_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__98_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__98_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__98_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__98_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__98_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__98_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__98_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__98_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__98_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__98_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__98_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__98_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__98_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__98_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__98_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__98_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__98_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__98_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__98_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__1_
  (
    .clk_1_S_out(clk_1_wires[174]),
    .clk_1_N_out(clk_1_wires[173]),
    .clk_1_W_in(clk_1_wires[169]),
    .prog_clk_1_S_out(prog_clk_1_wires[174]),
    .prog_clk_1_N_out(prog_clk_1_wires[173]),
    .prog_clk_1_W_in(prog_clk_1_wires[169]),
    .prog_clk_0_N_in(prog_clk_0_wires[370]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[99]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[99]),
    .SC_OUT_TOP(scff_Wires[242]),
    .SC_IN_BOT(scff_Wires[241]),
    .chanx_left_in(sb_1__1__88_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__99_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__99_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__99_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__99_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__99_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__99_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__99_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__99_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__99_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__99_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__99_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__99_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__99_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__99_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__99_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__99_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__99_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__99_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__99_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__99_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__99_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[373]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[100]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[100]),
    .SC_OUT_TOP(scff_Wires[244]),
    .SC_IN_BOT(scff_Wires[243]),
    .chanx_left_in(sb_1__1__89_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__100_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__100_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__100_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__100_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__100_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__100_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__100_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__100_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__100_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__100_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__100_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__100_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__100_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__100_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__100_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__100_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__100_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__100_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__100_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__100_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__100_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__3_
  (
    .clk_1_S_out(clk_1_wires[181]),
    .clk_1_N_out(clk_1_wires[180]),
    .clk_1_W_in(clk_1_wires[176]),
    .prog_clk_1_S_out(prog_clk_1_wires[181]),
    .prog_clk_1_N_out(prog_clk_1_wires[180]),
    .prog_clk_1_W_in(prog_clk_1_wires[176]),
    .prog_clk_0_N_in(prog_clk_0_wires[376]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[101]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[101]),
    .SC_OUT_TOP(scff_Wires[246]),
    .SC_IN_BOT(scff_Wires[245]),
    .chanx_left_in(sb_1__1__90_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__101_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__101_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__101_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__101_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__101_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__101_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__101_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__101_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__101_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__101_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__101_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__101_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__101_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__101_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__101_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__101_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__101_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__101_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__101_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__101_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__101_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[379]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[102]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[102]),
    .SC_OUT_TOP(scff_Wires[248]),
    .SC_IN_BOT(scff_Wires[247]),
    .chanx_left_in(sb_1__1__91_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__102_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__102_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__102_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__102_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__102_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__102_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__102_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__102_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__102_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__102_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__102_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__102_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__102_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__102_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__102_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__102_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__102_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__102_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__102_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__102_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__102_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__5_
  (
    .clk_1_S_out(clk_1_wires[188]),
    .clk_1_N_out(clk_1_wires[187]),
    .clk_1_W_in(clk_1_wires[183]),
    .prog_clk_1_S_out(prog_clk_1_wires[188]),
    .prog_clk_1_N_out(prog_clk_1_wires[187]),
    .prog_clk_1_W_in(prog_clk_1_wires[183]),
    .prog_clk_0_N_in(prog_clk_0_wires[382]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[103]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[103]),
    .SC_OUT_TOP(scff_Wires[250]),
    .SC_IN_BOT(scff_Wires[249]),
    .chanx_left_in(sb_1__1__92_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__103_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__103_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__103_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__103_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__103_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__103_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__103_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__103_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__103_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__103_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__103_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__103_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__103_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__103_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__103_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__103_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__103_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__103_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__103_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__103_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__103_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__6_
  (
    .clk_3_E_out(clk_3_wires[49]),
    .clk_3_W_in(clk_3_wires[48]),
    .prog_clk_3_E_out(prog_clk_3_wires[49]),
    .prog_clk_3_W_in(prog_clk_3_wires[48]),
    .prog_clk_0_N_in(prog_clk_0_wires[385]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[104]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[104]),
    .SC_OUT_TOP(scff_Wires[252]),
    .SC_IN_BOT(scff_Wires[251]),
    .chanx_left_in(sb_1__1__93_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__104_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__104_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__104_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__104_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__104_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__104_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__104_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__104_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__104_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__104_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__104_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__104_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__104_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__104_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__104_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__104_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__104_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__104_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__104_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__104_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__104_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__7_
  (
    .clk_1_S_out(clk_1_wires[195]),
    .clk_1_N_out(clk_1_wires[194]),
    .clk_1_W_in(clk_1_wires[190]),
    .prog_clk_1_S_out(prog_clk_1_wires[195]),
    .prog_clk_1_N_out(prog_clk_1_wires[194]),
    .prog_clk_1_W_in(prog_clk_1_wires[190]),
    .prog_clk_0_N_in(prog_clk_0_wires[388]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[105]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[105]),
    .SC_OUT_TOP(scff_Wires[254]),
    .SC_IN_BOT(scff_Wires[253]),
    .chanx_left_in(sb_1__1__94_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__105_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__105_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__105_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__105_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__105_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__105_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__105_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__105_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__105_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__105_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__105_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__105_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__105_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__105_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__105_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__105_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__105_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__105_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__105_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__105_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__105_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[391]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[106]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[106]),
    .SC_OUT_TOP(scff_Wires[256]),
    .SC_IN_BOT(scff_Wires[255]),
    .chanx_left_in(sb_1__1__95_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__106_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__106_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__106_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__106_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__106_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__106_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__106_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__106_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__106_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__106_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__106_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__106_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__106_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__106_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__106_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__106_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__106_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__106_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__106_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__106_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__106_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__9_
  (
    .clk_1_S_out(clk_1_wires[202]),
    .clk_1_N_out(clk_1_wires[201]),
    .clk_1_W_in(clk_1_wires[197]),
    .prog_clk_1_S_out(prog_clk_1_wires[202]),
    .prog_clk_1_N_out(prog_clk_1_wires[201]),
    .prog_clk_1_W_in(prog_clk_1_wires[197]),
    .prog_clk_0_N_in(prog_clk_0_wires[394]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[107]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[107]),
    .SC_OUT_TOP(scff_Wires[258]),
    .SC_IN_BOT(scff_Wires[257]),
    .chanx_left_in(sb_1__1__96_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__107_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__107_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__107_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__107_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__107_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__107_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__107_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__107_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__107_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__107_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__107_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__107_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__107_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__107_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__107_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__107_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__107_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__107_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__107_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__107_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__107_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[397]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[108]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[108]),
    .SC_OUT_TOP(scff_Wires[260]),
    .SC_IN_BOT(scff_Wires[259]),
    .chanx_left_in(sb_1__1__97_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__108_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__108_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__108_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__108_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__108_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__108_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__108_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__108_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__108_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__108_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__108_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__108_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__108_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__108_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__108_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__108_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__108_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__108_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__108_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__108_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__108_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__11_
  (
    .clk_1_S_out(clk_1_wires[209]),
    .clk_1_N_out(clk_1_wires[208]),
    .clk_1_W_in(clk_1_wires[204]),
    .prog_clk_1_S_out(prog_clk_1_wires[209]),
    .prog_clk_1_N_out(prog_clk_1_wires[208]),
    .prog_clk_1_W_in(prog_clk_1_wires[204]),
    .prog_clk_0_N_in(prog_clk_0_wires[400]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[109]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[109]),
    .SC_OUT_TOP(scff_Wires[262]),
    .SC_IN_BOT(scff_Wires[261]),
    .chanx_left_in(sb_1__1__98_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__109_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__109_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__109_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__109_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__109_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__109_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__109_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__109_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__109_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__109_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__109_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__109_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__109_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__109_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__109_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__109_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__109_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__109_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__109_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__109_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__109_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__1_
  (
    .clk_1_S_out(clk_1_wires[214]),
    .clk_1_N_out(clk_1_wires[213]),
    .clk_1_E_in(clk_1_wires[212]),
    .prog_clk_1_S_out(prog_clk_1_wires[214]),
    .prog_clk_1_N_out(prog_clk_1_wires[213]),
    .prog_clk_1_E_in(prog_clk_1_wires[212]),
    .prog_clk_0_N_in(prog_clk_0_wires[408]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[110]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[110]),
    .SC_OUT_BOT(scff_Wires[288]),
    .SC_IN_TOP(scff_Wires[287]),
    .chanx_left_in(sb_1__1__99_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__110_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__110_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__110_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__110_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__110_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__110_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__110_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__110_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__110_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__110_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__110_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__110_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__110_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__110_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__110_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__110_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__110_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__110_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__110_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__110_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__110_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__2_
  (
    .clk_2_W_in(clk_2_wires[114]),
    .clk_2_E_out(clk_2_wires[113]),
    .prog_clk_2_W_in(prog_clk_2_wires[114]),
    .prog_clk_2_E_out(prog_clk_2_wires[113]),
    .prog_clk_0_N_in(prog_clk_0_wires[411]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[111]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[111]),
    .SC_OUT_BOT(scff_Wires[286]),
    .SC_IN_TOP(scff_Wires[285]),
    .chanx_left_in(sb_1__1__100_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__111_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__111_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__111_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__111_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__111_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__111_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__111_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__111_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__111_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__111_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__111_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__111_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__111_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__111_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__111_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__111_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__111_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__111_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__111_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__111_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__111_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__3_
  (
    .clk_1_S_out(clk_1_wires[221]),
    .clk_1_N_out(clk_1_wires[220]),
    .clk_1_E_in(clk_1_wires[219]),
    .prog_clk_1_S_out(prog_clk_1_wires[221]),
    .prog_clk_1_N_out(prog_clk_1_wires[220]),
    .prog_clk_1_E_in(prog_clk_1_wires[219]),
    .prog_clk_0_N_in(prog_clk_0_wires[414]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[112]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[112]),
    .SC_OUT_BOT(scff_Wires[284]),
    .SC_IN_TOP(scff_Wires[283]),
    .chanx_left_in(sb_1__1__101_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__112_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__112_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__112_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__112_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__112_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__112_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__112_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__112_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__112_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__112_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__112_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__112_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__112_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__112_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__112_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__112_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__112_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__112_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__112_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__112_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__112_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__4_
  (
    .clk_2_W_in(clk_2_wires[119]),
    .clk_2_E_out(clk_2_wires[118]),
    .prog_clk_2_W_in(prog_clk_2_wires[119]),
    .prog_clk_2_E_out(prog_clk_2_wires[118]),
    .prog_clk_0_N_in(prog_clk_0_wires[417]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[113]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[113]),
    .SC_OUT_BOT(scff_Wires[282]),
    .SC_IN_TOP(scff_Wires[281]),
    .chanx_left_in(sb_1__1__102_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__113_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__113_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__113_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__113_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__113_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__113_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__113_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__113_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__113_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__113_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__113_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__113_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__113_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__113_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__113_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__113_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__113_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__113_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__113_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__113_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__113_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__5_
  (
    .clk_1_S_out(clk_1_wires[228]),
    .clk_1_N_out(clk_1_wires[227]),
    .clk_1_E_in(clk_1_wires[226]),
    .prog_clk_1_S_out(prog_clk_1_wires[228]),
    .prog_clk_1_N_out(prog_clk_1_wires[227]),
    .prog_clk_1_E_in(prog_clk_1_wires[226]),
    .prog_clk_0_N_in(prog_clk_0_wires[420]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[114]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[114]),
    .SC_OUT_BOT(scff_Wires[280]),
    .SC_IN_TOP(scff_Wires[279]),
    .chanx_left_in(sb_1__1__103_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__114_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__114_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__114_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__114_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__114_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__114_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__114_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__114_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__114_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__114_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__114_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__114_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__114_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__114_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__114_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__114_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__114_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__114_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__114_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__114_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__114_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[423]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[115]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[115]),
    .SC_OUT_BOT(scff_Wires[278]),
    .SC_IN_TOP(scff_Wires[277]),
    .chanx_left_in(sb_1__1__104_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__115_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__115_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__115_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__115_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__115_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__115_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__115_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__115_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__115_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__115_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__115_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__115_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__115_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__115_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__115_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__115_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__115_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__115_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__115_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__115_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__115_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__7_
  (
    .clk_1_S_out(clk_1_wires[235]),
    .clk_1_N_out(clk_1_wires[234]),
    .clk_1_E_in(clk_1_wires[233]),
    .prog_clk_1_S_out(prog_clk_1_wires[235]),
    .prog_clk_1_N_out(prog_clk_1_wires[234]),
    .prog_clk_1_E_in(prog_clk_1_wires[233]),
    .prog_clk_0_N_in(prog_clk_0_wires[426]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[116]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[116]),
    .SC_OUT_BOT(scff_Wires[276]),
    .SC_IN_TOP(scff_Wires[275]),
    .chanx_left_in(sb_1__1__105_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__116_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__116_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__116_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__116_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__116_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__116_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__116_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__116_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__116_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__116_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__116_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__116_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__116_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__116_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__116_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__116_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__116_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__116_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__116_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__116_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__116_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__8_
  (
    .clk_2_W_in(clk_2_wires[126]),
    .clk_2_E_out(clk_2_wires[125]),
    .prog_clk_2_W_in(prog_clk_2_wires[126]),
    .prog_clk_2_E_out(prog_clk_2_wires[125]),
    .prog_clk_0_N_in(prog_clk_0_wires[429]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[117]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[117]),
    .SC_OUT_BOT(scff_Wires[274]),
    .SC_IN_TOP(scff_Wires[273]),
    .chanx_left_in(sb_1__1__106_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__117_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__117_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__117_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__117_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__117_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__117_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__117_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__117_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__117_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__117_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__117_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__117_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__117_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__117_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__117_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__117_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__117_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__117_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__117_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__117_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__117_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__9_
  (
    .clk_1_S_out(clk_1_wires[242]),
    .clk_1_N_out(clk_1_wires[241]),
    .clk_1_E_in(clk_1_wires[240]),
    .prog_clk_1_S_out(prog_clk_1_wires[242]),
    .prog_clk_1_N_out(prog_clk_1_wires[241]),
    .prog_clk_1_E_in(prog_clk_1_wires[240]),
    .prog_clk_0_N_in(prog_clk_0_wires[432]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[118]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[118]),
    .SC_OUT_BOT(scff_Wires[272]),
    .SC_IN_TOP(scff_Wires[271]),
    .chanx_left_in(sb_1__1__107_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__118_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__118_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__118_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__118_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__118_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__118_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__118_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__118_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__118_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__118_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__118_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__118_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__118_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__118_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__118_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__118_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__118_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__118_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__118_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__118_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__118_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__10_
  (
    .clk_2_W_in(clk_2_wires[133]),
    .clk_2_E_out(clk_2_wires[132]),
    .prog_clk_2_W_in(prog_clk_2_wires[133]),
    .prog_clk_2_E_out(prog_clk_2_wires[132]),
    .prog_clk_0_N_in(prog_clk_0_wires[435]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[119]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[119]),
    .SC_OUT_BOT(scff_Wires[270]),
    .SC_IN_TOP(scff_Wires[269]),
    .chanx_left_in(sb_1__1__108_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__119_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__119_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__119_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__119_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__119_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__119_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__119_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__119_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__119_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__119_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__119_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__119_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__119_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__119_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__119_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__119_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__119_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__119_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__119_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__119_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__119_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__11_
  (
    .clk_1_S_out(clk_1_wires[249]),
    .clk_1_N_out(clk_1_wires[248]),
    .clk_1_E_in(clk_1_wires[247]),
    .prog_clk_1_S_out(prog_clk_1_wires[249]),
    .prog_clk_1_N_out(prog_clk_1_wires[248]),
    .prog_clk_1_E_in(prog_clk_1_wires[247]),
    .prog_clk_0_N_in(prog_clk_0_wires[438]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[120]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[120]),
    .SC_OUT_BOT(scff_Wires[268]),
    .SC_IN_TOP(scff_Wires[267]),
    .chanx_left_in(sb_1__1__109_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__120_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__120_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__120_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__120_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__120_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__120_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__120_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__120_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__120_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__120_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__120_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__120_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__120_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__120_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__120_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__120_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__120_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__120_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__120_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__120_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__120_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__1_
  (
    .clk_1_S_out(clk_1_wires[216]),
    .clk_1_N_out(clk_1_wires[215]),
    .clk_1_W_in(clk_1_wires[211]),
    .prog_clk_1_S_out(prog_clk_1_wires[216]),
    .prog_clk_1_N_out(prog_clk_1_wires[215]),
    .prog_clk_1_W_in(prog_clk_1_wires[211]),
    .prog_clk_0_N_in(prog_clk_0_wires[446]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[121]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[121]),
    .SC_OUT_TOP(scff_Wires[295]),
    .SC_IN_BOT(scff_Wires[294]),
    .chanx_left_in(sb_1__1__110_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__0_chanx_left_out[0:19]),
    .ccff_head(sb_12__1__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__121_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__121_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__121_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__121_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__121_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__121_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__121_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__121_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__121_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__121_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__121_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__121_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__121_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__121_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__121_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__121_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__121_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__121_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__121_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[449]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[122]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[122]),
    .SC_OUT_TOP(scff_Wires[297]),
    .SC_IN_BOT(scff_Wires[296]),
    .chanx_left_in(sb_1__1__111_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__1_chanx_left_out[0:19]),
    .ccff_head(sb_12__1__1_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__122_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__122_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__122_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__122_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__122_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__122_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__122_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__122_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__122_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__122_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__122_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__122_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__122_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__122_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__122_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__122_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__122_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__122_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__122_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__3_
  (
    .clk_1_S_out(clk_1_wires[223]),
    .clk_1_N_out(clk_1_wires[222]),
    .clk_1_W_in(clk_1_wires[218]),
    .prog_clk_1_S_out(prog_clk_1_wires[223]),
    .prog_clk_1_N_out(prog_clk_1_wires[222]),
    .prog_clk_1_W_in(prog_clk_1_wires[218]),
    .prog_clk_0_N_in(prog_clk_0_wires[452]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[123]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[123]),
    .SC_OUT_TOP(scff_Wires[299]),
    .SC_IN_BOT(scff_Wires[298]),
    .chanx_left_in(sb_1__1__112_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__2_chanx_left_out[0:19]),
    .ccff_head(sb_12__1__2_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__123_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__123_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__123_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__123_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__123_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__123_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__123_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__123_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__123_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__123_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__123_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__123_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__123_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__123_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__123_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__123_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__123_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__123_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__123_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[455]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[124]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[124]),
    .SC_OUT_TOP(scff_Wires[301]),
    .SC_IN_BOT(scff_Wires[300]),
    .chanx_left_in(sb_1__1__113_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__3_chanx_left_out[0:19]),
    .ccff_head(sb_12__1__3_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__124_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__124_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__124_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__124_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__124_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__124_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__124_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__124_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__124_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__124_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__124_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__124_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__124_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__124_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__124_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__124_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__124_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__124_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__124_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__5_
  (
    .clk_1_S_out(clk_1_wires[230]),
    .clk_1_N_out(clk_1_wires[229]),
    .clk_1_W_in(clk_1_wires[225]),
    .prog_clk_1_S_out(prog_clk_1_wires[230]),
    .prog_clk_1_N_out(prog_clk_1_wires[229]),
    .prog_clk_1_W_in(prog_clk_1_wires[225]),
    .prog_clk_0_N_in(prog_clk_0_wires[458]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[125]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[125]),
    .SC_OUT_TOP(scff_Wires[303]),
    .SC_IN_BOT(scff_Wires[302]),
    .chanx_left_in(sb_1__1__114_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__4_chanx_left_out[0:19]),
    .ccff_head(sb_12__1__4_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__125_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__125_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__125_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__125_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__125_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__125_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__125_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__125_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__125_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__125_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__125_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__125_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__125_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__125_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__125_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__125_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__125_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__125_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__125_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[461]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[126]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[126]),
    .SC_OUT_TOP(scff_Wires[305]),
    .SC_IN_BOT(scff_Wires[304]),
    .chanx_left_in(sb_1__1__115_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__5_chanx_left_out[0:19]),
    .ccff_head(sb_12__1__5_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__126_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__126_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__126_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__126_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__126_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__126_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__126_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__126_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__126_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__126_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__126_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__126_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__126_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__126_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__126_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__126_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__126_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__126_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__126_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__7_
  (
    .clk_1_S_out(clk_1_wires[237]),
    .clk_1_N_out(clk_1_wires[236]),
    .clk_1_W_in(clk_1_wires[232]),
    .prog_clk_1_S_out(prog_clk_1_wires[237]),
    .prog_clk_1_N_out(prog_clk_1_wires[236]),
    .prog_clk_1_W_in(prog_clk_1_wires[232]),
    .prog_clk_0_N_in(prog_clk_0_wires[464]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[127]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[127]),
    .SC_OUT_TOP(scff_Wires[307]),
    .SC_IN_BOT(scff_Wires[306]),
    .chanx_left_in(sb_1__1__116_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__6_chanx_left_out[0:19]),
    .ccff_head(sb_12__1__6_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__127_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__127_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__127_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__127_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__127_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__127_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__127_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__127_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__127_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__127_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__127_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__127_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__127_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__127_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__127_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__127_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__127_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__127_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__127_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[467]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[128]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[128]),
    .SC_OUT_TOP(scff_Wires[309]),
    .SC_IN_BOT(scff_Wires[308]),
    .chanx_left_in(sb_1__1__117_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__7_chanx_left_out[0:19]),
    .ccff_head(sb_12__1__7_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__128_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__128_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__128_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__128_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__128_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__128_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__128_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__128_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__128_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__128_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__128_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__128_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__128_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__128_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__128_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__128_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__128_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__128_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__128_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__9_
  (
    .clk_1_S_out(clk_1_wires[244]),
    .clk_1_N_out(clk_1_wires[243]),
    .clk_1_W_in(clk_1_wires[239]),
    .prog_clk_1_S_out(prog_clk_1_wires[244]),
    .prog_clk_1_N_out(prog_clk_1_wires[243]),
    .prog_clk_1_W_in(prog_clk_1_wires[239]),
    .prog_clk_0_N_in(prog_clk_0_wires[470]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[129]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[129]),
    .SC_OUT_TOP(scff_Wires[311]),
    .SC_IN_BOT(scff_Wires[310]),
    .chanx_left_in(sb_1__1__118_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__8_chanx_left_out[0:19]),
    .ccff_head(sb_12__1__8_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__129_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__129_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__129_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__129_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__129_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__129_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__129_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__129_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__129_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__129_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__129_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__129_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__129_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__129_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__129_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__129_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__129_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__129_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__129_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[473]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[130]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[130]),
    .SC_OUT_TOP(scff_Wires[313]),
    .SC_IN_BOT(scff_Wires[312]),
    .chanx_left_in(sb_1__1__119_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__9_chanx_left_out[0:19]),
    .ccff_head(sb_12__1__9_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__130_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__130_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__130_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__130_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__130_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__130_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__130_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__130_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__130_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__130_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__130_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__130_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__130_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__130_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__130_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__130_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__130_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__130_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__130_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__11_
  (
    .clk_1_S_out(clk_1_wires[251]),
    .clk_1_N_out(clk_1_wires[250]),
    .clk_1_W_in(clk_1_wires[246]),
    .prog_clk_1_S_out(prog_clk_1_wires[251]),
    .prog_clk_1_N_out(prog_clk_1_wires[250]),
    .prog_clk_1_W_in(prog_clk_1_wires[246]),
    .prog_clk_0_N_in(prog_clk_0_wires[476]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[131]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[131]),
    .SC_OUT_TOP(scff_Wires[315]),
    .SC_IN_BOT(scff_Wires[314]),
    .chanx_left_in(sb_1__1__120_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__1__10_chanx_left_out[0:19]),
    .ccff_head(sb_12__1__10_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__131_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__131_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__131_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__131_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__131_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__131_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__131_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__131_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__131_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__131_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__131_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__131_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__131_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__131_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__131_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__131_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__131_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__131_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__131_ccff_tail[0])
  );


  cbx_1__2_
  cbx_1__12_
  (
    .prog_clk_0_W_out(prog_clk_0_wires[62]),
    .prog_clk_0_S_in(prog_clk_0_wires[59]),
    .SC_OUT_BOT(scff_Wires[1]),
    .SC_IN_TOP(scff_Wires[0]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_0_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_0_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__0_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_0__12__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__12__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__0_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__12__0_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__0_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__0_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__0_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__0_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__0_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__0_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__0_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__0_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__0_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__0_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__0_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__0_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__0_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__0_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__0_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__0_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_0_ccff_tail[0])
  );


  cbx_1__2_
  cbx_2__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[99]),
    .SC_OUT_TOP(scff_Wires[52]),
    .SC_IN_BOT(scff_Wires[51]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_1_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_1_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__1_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__12__1_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__1_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__12__1_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__1_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__1_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__1_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__1_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__1_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__1_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__1_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__1_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__1_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__1_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__1_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__1_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__1_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__1_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__1_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__1_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_1_ccff_tail[0])
  );


  cbx_1__2_
  cbx_3__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[137]),
    .SC_OUT_BOT(scff_Wires[54]),
    .SC_IN_TOP(scff_Wires[53]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_2_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_2_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__2_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__12__2_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__2_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__12__2_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__2_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__2_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__2_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__2_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__2_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__2_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__2_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__2_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__2_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__2_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__2_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__2_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__2_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__2_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__2_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__2_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_2_ccff_tail[0])
  );


  cbx_1__2_
  cbx_4__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[175]),
    .SC_OUT_TOP(scff_Wires[105]),
    .SC_IN_BOT(scff_Wires[104]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_3_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_3_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__3_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__12__3_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__3_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__12__3_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__3_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__3_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__3_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__3_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__3_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__3_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__3_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__3_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__3_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__3_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__3_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__3_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__3_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__3_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__3_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__3_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_3_ccff_tail[0])
  );


  cbx_1__2_
  cbx_5__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[213]),
    .SC_OUT_BOT(scff_Wires[107]),
    .SC_IN_TOP(scff_Wires[106]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_4_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_4_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__4_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__12__4_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__4_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__12__4_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__4_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__4_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__4_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__4_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__4_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__4_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__4_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__4_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__4_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__4_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__4_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__4_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__4_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__4_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__4_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__4_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_4_ccff_tail[0])
  );


  cbx_1__2_
  cbx_6__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[251]),
    .SC_OUT_TOP(scff_Wires[158]),
    .SC_IN_BOT(scff_Wires[157]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_5_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_5_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__5_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__12__5_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__5_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__12__5_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__5_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__5_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__5_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__5_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__5_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__5_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__5_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__5_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__5_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__5_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__5_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__5_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__5_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__5_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__5_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__5_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_5_ccff_tail[0])
  );


  cbx_1__2_
  cbx_7__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[289]),
    .SC_OUT_BOT(scff_Wires[160]),
    .SC_IN_TOP(scff_Wires[159]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_6_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_6_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__6_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__12__6_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__6_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__12__6_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__6_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__6_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__6_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__6_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__6_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__6_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__6_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__6_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__6_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__6_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__6_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__6_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__6_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__6_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__6_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__6_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_6_ccff_tail[0])
  );


  cbx_1__2_
  cbx_8__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[327]),
    .SC_OUT_TOP(scff_Wires[211]),
    .SC_IN_BOT(scff_Wires[210]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_7_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_7_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__7_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__7_chanx_left_out[0:19]),
    .ccff_head(sb_1__12__7_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__7_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__12__7_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__7_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__7_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__7_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__7_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__7_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__7_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__7_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__7_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__7_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__7_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__7_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__7_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__7_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__7_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__7_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__7_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_7_ccff_tail[0])
  );


  cbx_1__2_
  cbx_9__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[365]),
    .SC_OUT_BOT(scff_Wires[213]),
    .SC_IN_TOP(scff_Wires[212]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_8_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_8_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__8_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__8_chanx_left_out[0:19]),
    .ccff_head(sb_1__12__8_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__8_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__12__8_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__8_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__8_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__8_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__8_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__8_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__8_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__8_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__8_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__8_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__8_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__8_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__8_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__8_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__8_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__8_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__8_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_8_ccff_tail[0])
  );


  cbx_1__2_
  cbx_10__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[403]),
    .SC_OUT_TOP(scff_Wires[264]),
    .SC_IN_BOT(scff_Wires[263]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_9_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_9_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__9_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__9_chanx_left_out[0:19]),
    .ccff_head(sb_1__12__9_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__9_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__12__9_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__9_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__9_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__9_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__9_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__9_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__9_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__9_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__9_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__9_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__9_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__9_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__9_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__9_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__9_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__9_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__9_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_9_ccff_tail[0])
  );


  cbx_1__2_
  cbx_11__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[441]),
    .SC_OUT_BOT(scff_Wires[266]),
    .SC_IN_TOP(scff_Wires[265]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_10_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_10_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__10_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__12__10_chanx_left_out[0:19]),
    .ccff_head(sb_1__12__10_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__10_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__12__10_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__10_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__10_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__10_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__10_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__10_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__10_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__10_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__10_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__10_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__10_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__10_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__10_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__10_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__10_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__10_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__10_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_10_ccff_tail[0])
  );


  cbx_1__2_
  cbx_12__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[479]),
    .SC_OUT_TOP(scff_Wires[317]),
    .SC_IN_BOT(scff_Wires[316]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_11_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_11_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__11_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_12__12__0_chanx_left_out[0:19]),
    .ccff_head(sb_12__12__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__12__11_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__12__11_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__11_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__11_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__11_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__11_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__11_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__11_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__11_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__11_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__11_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__11_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__11_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__11_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__11_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__11_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__11_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__11_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_11_ccff_tail[0])
  );


  cby_0__1_
  cby_0__1_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[3]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_0_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_0_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__0_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[132]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[132]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[132]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__0__0_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__0_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__0_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__0_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__0_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_0_ccff_tail[0])
  );


  cby_0__1_
  cby_0__2_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[9]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_1_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_1_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__1_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[133]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[133]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[133]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__0_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__1_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__1_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__1_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__1_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_1_ccff_tail[0])
  );


  cby_0__1_
  cby_0__3_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[14]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_2_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_2_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__2_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[134]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[134]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[134]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__1_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__2_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__2_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__2_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__2_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_2_ccff_tail[0])
  );


  cby_0__1_
  cby_0__4_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[19]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_3_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_3_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__3_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[135]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[135]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[135]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__2_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__3_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__3_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__3_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__3_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_3_ccff_tail[0])
  );


  cby_0__1_
  cby_0__5_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[24]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_4_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_4_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__4_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[136]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[136]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[136]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__3_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__4_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__4_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__4_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__4_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_4_ccff_tail[0])
  );


  cby_0__1_
  cby_0__6_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[29]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_5_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_5_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__5_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[137]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[137]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[137]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__4_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__5_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__5_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__5_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__5_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_5_ccff_tail[0])
  );


  cby_0__1_
  cby_0__7_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[34]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_6_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_6_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__6_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[138]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[138]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[138]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__5_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__6_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__6_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__6_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__6_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_6_ccff_tail[0])
  );


  cby_0__1_
  cby_0__8_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[39]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_7_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_7_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__7_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[139]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[139]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[139]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__6_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__7_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__7_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__7_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__7_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_7_ccff_tail[0])
  );


  cby_0__1_
  cby_0__9_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[44]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_8_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_8_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__8_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[140]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[140]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[140]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__7_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__8_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__8_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__8_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__8_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__8_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_8_ccff_tail[0])
  );


  cby_0__1_
  cby_0__10_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[49]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_9_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_9_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__9_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[141]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[141]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[141]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__8_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__9_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__9_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__9_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__9_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__9_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_9_ccff_tail[0])
  );


  cby_0__1_
  cby_0__11_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[54]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_10_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_10_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__10_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[142]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[142]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[142]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__9_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__10_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__10_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__10_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__10_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__10_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_10_ccff_tail[0])
  );


  cby_0__1_
  cby_0__12_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[61]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_11_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_11_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__11_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[143]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[143]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[143]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__10_chany_top_out[0:19]),
    .chany_top_in(sb_0__12__0_chany_bottom_out[0:19]),
    .ccff_head(sb_0__12__0_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__11_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__11_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__11_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_11_ccff_tail[0])
  );


  cby_1__1_
  cby_1__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[2]),
    .prog_clk_0_W_in(prog_clk_0_wires[1]),
    .Test_en_E_in(Test_enWires[26]),
    .Test_en_W_out(Test_enWires[24]),
    .chany_bottom_in(sb_1__0__0_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_0_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__0_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__0_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__0_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__0_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__0_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__0_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__0_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__0_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__0_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__0_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__0_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__0_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__0_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__0_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__0_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__0_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__0_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__0_ccff_tail[0])
  );


  cby_1__1_
  cby_1__2_
  (
    .clk_2_S_out(clk_2_wires[4]),
    .clk_2_N_in(clk_2_wires[3]),
    .prog_clk_2_S_out(prog_clk_2_wires[4]),
    .prog_clk_2_N_in(prog_clk_2_wires[3]),
    .prog_clk_0_S_out(prog_clk_0_wires[8]),
    .prog_clk_0_W_in(prog_clk_0_wires[7]),
    .Test_en_E_in(Test_enWires[48]),
    .Test_en_W_out(Test_enWires[46]),
    .chany_bottom_in(sb_1__1__0_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_1_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__1_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__1_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__1_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__1_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__1_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__1_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__1_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__1_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__1_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__1_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__1_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__1_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__1_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__1_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__1_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__1_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__1_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__1_ccff_tail[0])
  );


  cby_1__1_
  cby_1__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[13]),
    .prog_clk_0_W_in(prog_clk_0_wires[12]),
    .Test_en_E_in(Test_enWires[70]),
    .Test_en_W_out(Test_enWires[68]),
    .chany_bottom_in(sb_1__1__1_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_2_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__2_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__2_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__2_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__2_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__2_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__2_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__2_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__2_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__2_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__2_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__2_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__2_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__2_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__2_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__2_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__2_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__2_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__2_ccff_tail[0])
  );


  cby_1__1_
  cby_1__4_
  (
    .clk_2_S_out(clk_2_wires[11]),
    .clk_2_N_in(clk_2_wires[10]),
    .prog_clk_2_S_out(prog_clk_2_wires[11]),
    .prog_clk_2_N_in(prog_clk_2_wires[10]),
    .prog_clk_0_S_out(prog_clk_0_wires[18]),
    .prog_clk_0_W_in(prog_clk_0_wires[17]),
    .Test_en_E_in(Test_enWires[92]),
    .Test_en_W_out(Test_enWires[90]),
    .chany_bottom_in(sb_1__1__2_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_3_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__3_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__3_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__3_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__3_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__3_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__3_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__3_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__3_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__3_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__3_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__3_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__3_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__3_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__3_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__3_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__3_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__3_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__3_ccff_tail[0])
  );


  cby_1__1_
  cby_1__5_
  (
    .clk_2_N_out(clk_2_wires[9]),
    .clk_2_S_in(clk_2_wires[8]),
    .prog_clk_2_N_out(prog_clk_2_wires[9]),
    .prog_clk_2_S_in(prog_clk_2_wires[8]),
    .prog_clk_0_S_out(prog_clk_0_wires[23]),
    .prog_clk_0_W_in(prog_clk_0_wires[22]),
    .Test_en_E_in(Test_enWires[114]),
    .Test_en_W_out(Test_enWires[112]),
    .chany_bottom_in(sb_1__1__3_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_4_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__4_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__4_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__4_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__4_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__4_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__4_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__4_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__4_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__4_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__4_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__4_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__4_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__4_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__4_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__4_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__4_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__4_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__4_ccff_tail[0])
  );


  cby_1__1_
  cby_1__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[28]),
    .prog_clk_0_W_in(prog_clk_0_wires[27]),
    .Test_en_E_in(Test_enWires[136]),
    .Test_en_W_out(Test_enWires[134]),
    .chany_bottom_in(sb_1__1__4_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_5_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__5_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__5_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__5_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__5_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__5_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__5_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__5_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__5_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__5_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__5_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__5_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__5_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__5_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__5_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__5_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__5_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__5_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__5_ccff_tail[0])
  );


  cby_1__1_
  cby_1__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[33]),
    .prog_clk_0_W_in(prog_clk_0_wires[32]),
    .Test_en_E_in(Test_enWires[158]),
    .Test_en_W_out(Test_enWires[156]),
    .chany_bottom_in(sb_1__1__5_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_6_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__6_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__6_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__6_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__6_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__6_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__6_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__6_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__6_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__6_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__6_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__6_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__6_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__6_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__6_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__6_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__6_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__6_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__6_ccff_tail[0])
  );


  cby_1__1_
  cby_1__8_
  (
    .clk_2_S_out(clk_2_wires[18]),
    .clk_2_N_in(clk_2_wires[17]),
    .prog_clk_2_S_out(prog_clk_2_wires[18]),
    .prog_clk_2_N_in(prog_clk_2_wires[17]),
    .prog_clk_0_S_out(prog_clk_0_wires[38]),
    .prog_clk_0_W_in(prog_clk_0_wires[37]),
    .Test_en_E_in(Test_enWires[180]),
    .Test_en_W_out(Test_enWires[178]),
    .chany_bottom_in(sb_1__1__6_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__7_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_7_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__7_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__7_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__7_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__7_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__7_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__7_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__7_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__7_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__7_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__7_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__7_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__7_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__7_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__7_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__7_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__7_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__7_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__7_ccff_tail[0])
  );


  cby_1__1_
  cby_1__9_
  (
    .clk_2_N_out(clk_2_wires[16]),
    .clk_2_S_in(clk_2_wires[15]),
    .prog_clk_2_N_out(prog_clk_2_wires[16]),
    .prog_clk_2_S_in(prog_clk_2_wires[15]),
    .prog_clk_0_S_out(prog_clk_0_wires[43]),
    .prog_clk_0_W_in(prog_clk_0_wires[42]),
    .Test_en_E_in(Test_enWires[202]),
    .Test_en_W_out(Test_enWires[200]),
    .chany_bottom_in(sb_1__1__7_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__8_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_8_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__8_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__8_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__8_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__8_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__8_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__8_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__8_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__8_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__8_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__8_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__8_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__8_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__8_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__8_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__8_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__8_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__8_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__8_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__8_ccff_tail[0])
  );


  cby_1__1_
  cby_1__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[48]),
    .prog_clk_0_W_in(prog_clk_0_wires[47]),
    .Test_en_E_in(Test_enWires[224]),
    .Test_en_W_out(Test_enWires[222]),
    .chany_bottom_in(sb_1__1__8_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__9_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_9_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__9_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__9_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__9_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__9_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__9_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__9_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__9_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__9_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__9_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__9_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__9_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__9_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__9_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__9_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__9_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__9_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__9_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__9_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__9_ccff_tail[0])
  );


  cby_1__1_
  cby_1__11_
  (
    .clk_2_N_out(clk_2_wires[23]),
    .clk_2_S_in(clk_2_wires[22]),
    .prog_clk_2_N_out(prog_clk_2_wires[23]),
    .prog_clk_2_S_in(prog_clk_2_wires[22]),
    .prog_clk_0_S_out(prog_clk_0_wires[53]),
    .prog_clk_0_W_in(prog_clk_0_wires[52]),
    .Test_en_E_in(Test_enWires[246]),
    .Test_en_W_out(Test_enWires[244]),
    .chany_bottom_in(sb_1__1__9_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__10_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_10_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__10_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__10_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__10_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__10_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__10_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__10_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__10_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__10_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__10_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__10_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__10_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__10_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__10_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__10_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__10_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__10_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__10_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__10_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__10_ccff_tail[0])
  );


  cby_1__1_
  cby_1__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[60]),
    .prog_clk_0_S_out(prog_clk_0_wires[58]),
    .prog_clk_0_W_in(prog_clk_0_wires[57]),
    .Test_en_E_in(Test_enWires[268]),
    .Test_en_W_out(Test_enWires[266]),
    .chany_bottom_in(sb_1__1__10_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_11_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__11_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__11_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__11_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__11_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__11_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__11_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__11_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__11_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__11_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__11_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__11_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__11_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__11_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__11_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__11_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__11_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__11_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__11_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__11_ccff_tail[0])
  );


  cby_1__1_
  cby_2__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[65]),
    .prog_clk_0_W_in(prog_clk_0_wires[64]),
    .Test_en_E_in(Test_enWires[28]),
    .Test_en_W_out(Test_enWires[25]),
    .chany_bottom_in(sb_1__0__1_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__11_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_12_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__12_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__12_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__12_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__12_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__12_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__12_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__12_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__12_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__12_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__12_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__12_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__12_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__12_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__12_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__12_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__12_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__12_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__12_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__12_ccff_tail[0])
  );


  cby_1__1_
  cby_2__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[68]),
    .prog_clk_0_W_in(prog_clk_0_wires[67]),
    .Test_en_E_in(Test_enWires[50]),
    .Test_en_W_out(Test_enWires[47]),
    .chany_bottom_in(sb_1__1__11_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__12_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_13_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__13_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__13_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__13_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__13_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__13_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__13_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__13_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__13_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__13_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__13_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__13_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__13_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__13_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__13_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__13_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__13_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__13_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__13_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__13_ccff_tail[0])
  );


  cby_1__1_
  cby_2__3_
  (
    .clk_3_S_out(clk_3_wires[69]),
    .clk_3_N_in(clk_3_wires[68]),
    .prog_clk_3_S_out(prog_clk_3_wires[69]),
    .prog_clk_3_N_in(prog_clk_3_wires[68]),
    .prog_clk_0_S_out(prog_clk_0_wires[71]),
    .prog_clk_0_W_in(prog_clk_0_wires[70]),
    .Test_en_E_in(Test_enWires[72]),
    .Test_en_W_out(Test_enWires[69]),
    .chany_bottom_in(sb_1__1__12_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__13_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_14_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__14_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__14_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__14_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__14_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__14_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__14_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__14_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__14_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__14_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__14_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__14_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__14_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__14_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__14_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__14_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__14_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__14_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__14_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__14_ccff_tail[0])
  );


  cby_1__1_
  cby_2__4_
  (
    .clk_3_S_out(clk_3_wires[65]),
    .clk_3_N_in(clk_3_wires[64]),
    .prog_clk_3_S_out(prog_clk_3_wires[65]),
    .prog_clk_3_N_in(prog_clk_3_wires[64]),
    .prog_clk_0_S_out(prog_clk_0_wires[74]),
    .prog_clk_0_W_in(prog_clk_0_wires[73]),
    .Test_en_E_in(Test_enWires[94]),
    .Test_en_W_out(Test_enWires[91]),
    .chany_bottom_in(sb_1__1__13_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__14_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_15_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__15_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__15_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__15_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__15_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__15_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__15_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__15_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__15_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__15_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__15_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__15_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__15_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__15_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__15_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__15_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__15_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__15_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__15_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__15_ccff_tail[0])
  );


  cby_1__1_
  cby_2__5_
  (
    .clk_3_S_out(clk_3_wires[59]),
    .clk_3_N_in(clk_3_wires[58]),
    .prog_clk_3_S_out(prog_clk_3_wires[59]),
    .prog_clk_3_N_in(prog_clk_3_wires[58]),
    .prog_clk_0_S_out(prog_clk_0_wires[77]),
    .prog_clk_0_W_in(prog_clk_0_wires[76]),
    .Test_en_E_in(Test_enWires[116]),
    .Test_en_W_out(Test_enWires[113]),
    .chany_bottom_in(sb_1__1__14_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__15_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_16_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__16_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__16_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__16_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__16_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__16_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__16_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__16_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__16_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__16_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__16_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__16_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__16_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__16_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__16_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__16_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__16_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__16_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__16_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__16_ccff_tail[0])
  );


  cby_1__1_
  cby_2__6_
  (
    .clk_3_S_out(clk_3_wires[55]),
    .clk_3_N_in(clk_3_wires[54]),
    .prog_clk_3_S_out(prog_clk_3_wires[55]),
    .prog_clk_3_N_in(prog_clk_3_wires[54]),
    .prog_clk_0_S_out(prog_clk_0_wires[80]),
    .prog_clk_0_W_in(prog_clk_0_wires[79]),
    .Test_en_E_in(Test_enWires[138]),
    .Test_en_W_out(Test_enWires[135]),
    .chany_bottom_in(sb_1__1__15_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__16_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_17_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__17_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__17_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__17_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__17_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__17_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__17_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__17_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__17_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__17_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__17_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__17_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__17_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__17_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__17_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__17_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__17_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__17_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__17_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__17_ccff_tail[0])
  );


  cby_1__1_
  cby_2__7_
  (
    .clk_3_N_out(clk_3_wires[53]),
    .clk_3_S_in(clk_3_wires[52]),
    .prog_clk_3_N_out(prog_clk_3_wires[53]),
    .prog_clk_3_S_in(prog_clk_3_wires[52]),
    .prog_clk_0_S_out(prog_clk_0_wires[83]),
    .prog_clk_0_W_in(prog_clk_0_wires[82]),
    .Test_en_E_in(Test_enWires[160]),
    .Test_en_W_out(Test_enWires[157]),
    .chany_bottom_in(sb_1__1__16_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__17_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_18_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__18_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__18_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__18_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__18_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__18_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__18_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__18_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__18_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__18_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__18_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__18_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__18_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__18_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__18_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__18_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__18_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__18_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__18_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__18_ccff_tail[0])
  );


  cby_1__1_
  cby_2__8_
  (
    .clk_3_N_out(clk_3_wires[57]),
    .clk_3_S_in(clk_3_wires[56]),
    .prog_clk_3_N_out(prog_clk_3_wires[57]),
    .prog_clk_3_S_in(prog_clk_3_wires[56]),
    .prog_clk_0_S_out(prog_clk_0_wires[86]),
    .prog_clk_0_W_in(prog_clk_0_wires[85]),
    .Test_en_E_in(Test_enWires[182]),
    .Test_en_W_out(Test_enWires[179]),
    .chany_bottom_in(sb_1__1__17_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__18_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_19_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__19_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__19_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__19_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__19_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__19_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__19_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__19_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__19_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__19_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__19_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__19_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__19_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__19_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__19_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__19_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__19_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__19_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__19_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__19_ccff_tail[0])
  );


  cby_1__1_
  cby_2__9_
  (
    .clk_3_N_out(clk_3_wires[63]),
    .clk_3_S_in(clk_3_wires[62]),
    .prog_clk_3_N_out(prog_clk_3_wires[63]),
    .prog_clk_3_S_in(prog_clk_3_wires[62]),
    .prog_clk_0_S_out(prog_clk_0_wires[89]),
    .prog_clk_0_W_in(prog_clk_0_wires[88]),
    .Test_en_E_in(Test_enWires[204]),
    .Test_en_W_out(Test_enWires[201]),
    .chany_bottom_in(sb_1__1__18_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__19_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_20_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__20_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__20_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__20_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__20_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__20_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__20_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__20_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__20_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__20_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__20_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__20_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__20_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__20_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__20_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__20_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__20_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__20_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__20_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__20_ccff_tail[0])
  );


  cby_1__1_
  cby_2__10_
  (
    .clk_3_N_out(clk_3_wires[67]),
    .clk_3_S_in(clk_3_wires[66]),
    .prog_clk_3_N_out(prog_clk_3_wires[67]),
    .prog_clk_3_S_in(prog_clk_3_wires[66]),
    .prog_clk_0_S_out(prog_clk_0_wires[92]),
    .prog_clk_0_W_in(prog_clk_0_wires[91]),
    .Test_en_E_in(Test_enWires[226]),
    .Test_en_W_out(Test_enWires[223]),
    .chany_bottom_in(sb_1__1__19_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__20_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_21_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__21_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__21_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__21_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__21_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__21_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__21_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__21_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__21_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__21_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__21_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__21_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__21_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__21_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__21_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__21_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__21_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__21_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__21_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__21_ccff_tail[0])
  );


  cby_1__1_
  cby_2__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[95]),
    .prog_clk_0_W_in(prog_clk_0_wires[94]),
    .Test_en_E_in(Test_enWires[248]),
    .Test_en_W_out(Test_enWires[245]),
    .chany_bottom_in(sb_1__1__20_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__21_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_22_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__22_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__22_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__22_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__22_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__22_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__22_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__22_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__22_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__22_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__22_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__22_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__22_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__22_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__22_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__22_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__22_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__22_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__22_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__22_ccff_tail[0])
  );


  cby_1__1_
  cby_2__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[100]),
    .prog_clk_0_S_out(prog_clk_0_wires[98]),
    .prog_clk_0_W_in(prog_clk_0_wires[97]),
    .Test_en_E_in(Test_enWires[270]),
    .Test_en_W_out(Test_enWires[267]),
    .chany_bottom_in(sb_1__1__21_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_23_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__23_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__23_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__23_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__23_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__23_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__23_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__23_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__23_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__23_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__23_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__23_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__23_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__23_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__23_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__23_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__23_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__23_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__23_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__23_ccff_tail[0])
  );


  cby_1__1_
  cby_3__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[103]),
    .prog_clk_0_W_in(prog_clk_0_wires[102]),
    .Test_en_E_in(Test_enWires[30]),
    .Test_en_W_out(Test_enWires[27]),
    .chany_bottom_in(sb_1__0__2_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__22_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_24_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__24_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__24_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__24_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__24_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__24_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__24_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__24_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__24_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__24_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__24_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__24_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__24_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__24_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__24_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__24_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__24_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__24_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__24_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__24_ccff_tail[0])
  );


  cby_1__1_
  cby_3__2_
  (
    .clk_2_S_out(clk_2_wires[30]),
    .clk_2_N_in(clk_2_wires[29]),
    .prog_clk_2_S_out(prog_clk_2_wires[30]),
    .prog_clk_2_N_in(prog_clk_2_wires[29]),
    .prog_clk_0_S_out(prog_clk_0_wires[106]),
    .prog_clk_0_W_in(prog_clk_0_wires[105]),
    .Test_en_E_in(Test_enWires[52]),
    .Test_en_W_out(Test_enWires[49]),
    .chany_bottom_in(sb_1__1__22_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__23_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_25_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__25_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__25_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__25_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__25_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__25_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__25_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__25_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__25_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__25_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__25_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__25_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__25_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__25_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__25_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__25_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__25_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__25_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__25_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__25_ccff_tail[0])
  );


  cby_1__1_
  cby_3__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[109]),
    .prog_clk_0_W_in(prog_clk_0_wires[108]),
    .Test_en_E_in(Test_enWires[74]),
    .Test_en_W_out(Test_enWires[71]),
    .chany_bottom_in(sb_1__1__23_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__24_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_26_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__26_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__26_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__26_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__26_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__26_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__26_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__26_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__26_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__26_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__26_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__26_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__26_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__26_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__26_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__26_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__26_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__26_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__26_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__26_ccff_tail[0])
  );


  cby_1__1_
  cby_3__4_
  (
    .clk_2_S_out(clk_2_wires[41]),
    .clk_2_N_in(clk_2_wires[40]),
    .prog_clk_2_S_out(prog_clk_2_wires[41]),
    .prog_clk_2_N_in(prog_clk_2_wires[40]),
    .prog_clk_0_S_out(prog_clk_0_wires[112]),
    .prog_clk_0_W_in(prog_clk_0_wires[111]),
    .Test_en_E_in(Test_enWires[96]),
    .Test_en_W_out(Test_enWires[93]),
    .chany_bottom_in(sb_1__1__24_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__25_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_27_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__27_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__27_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__27_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__27_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__27_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__27_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__27_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__27_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__27_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__27_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__27_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__27_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__27_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__27_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__27_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__27_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__27_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__27_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__27_ccff_tail[0])
  );


  cby_1__1_
  cby_3__5_
  (
    .clk_2_N_out(clk_2_wires[39]),
    .clk_2_S_in(clk_2_wires[38]),
    .prog_clk_2_N_out(prog_clk_2_wires[39]),
    .prog_clk_2_S_in(prog_clk_2_wires[38]),
    .prog_clk_0_S_out(prog_clk_0_wires[115]),
    .prog_clk_0_W_in(prog_clk_0_wires[114]),
    .Test_en_E_in(Test_enWires[118]),
    .Test_en_W_out(Test_enWires[115]),
    .chany_bottom_in(sb_1__1__25_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__26_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_28_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__28_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__28_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__28_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__28_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__28_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__28_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__28_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__28_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__28_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__28_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__28_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__28_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__28_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__28_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__28_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__28_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__28_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__28_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__28_ccff_tail[0])
  );


  cby_1__1_
  cby_3__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[118]),
    .prog_clk_0_W_in(prog_clk_0_wires[117]),
    .Test_en_E_in(Test_enWires[140]),
    .Test_en_W_out(Test_enWires[137]),
    .chany_bottom_in(sb_1__1__26_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__27_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_29_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__29_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__29_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__29_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__29_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__29_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__29_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__29_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__29_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__29_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__29_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__29_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__29_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__29_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__29_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__29_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__29_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__29_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__29_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__29_ccff_tail[0])
  );


  cby_1__1_
  cby_3__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[121]),
    .prog_clk_0_W_in(prog_clk_0_wires[120]),
    .Test_en_E_in(Test_enWires[162]),
    .Test_en_W_out(Test_enWires[159]),
    .chany_bottom_in(sb_1__1__27_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__28_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_30_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__30_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__30_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__30_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__30_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__30_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__30_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__30_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__30_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__30_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__30_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__30_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__30_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__30_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__30_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__30_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__30_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__30_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__30_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__30_ccff_tail[0])
  );


  cby_1__1_
  cby_3__8_
  (
    .clk_2_S_out(clk_2_wires[54]),
    .clk_2_N_in(clk_2_wires[53]),
    .prog_clk_2_S_out(prog_clk_2_wires[54]),
    .prog_clk_2_N_in(prog_clk_2_wires[53]),
    .prog_clk_0_S_out(prog_clk_0_wires[124]),
    .prog_clk_0_W_in(prog_clk_0_wires[123]),
    .Test_en_E_in(Test_enWires[184]),
    .Test_en_W_out(Test_enWires[181]),
    .chany_bottom_in(sb_1__1__28_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__29_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_31_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__31_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__31_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__31_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__31_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__31_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__31_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__31_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__31_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__31_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__31_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__31_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__31_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__31_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__31_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__31_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__31_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__31_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__31_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__31_ccff_tail[0])
  );


  cby_1__1_
  cby_3__9_
  (
    .clk_2_N_out(clk_2_wires[52]),
    .clk_2_S_in(clk_2_wires[51]),
    .prog_clk_2_N_out(prog_clk_2_wires[52]),
    .prog_clk_2_S_in(prog_clk_2_wires[51]),
    .prog_clk_0_S_out(prog_clk_0_wires[127]),
    .prog_clk_0_W_in(prog_clk_0_wires[126]),
    .Test_en_E_in(Test_enWires[206]),
    .Test_en_W_out(Test_enWires[203]),
    .chany_bottom_in(sb_1__1__29_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__30_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_32_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__32_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__32_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__32_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__32_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__32_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__32_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__32_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__32_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__32_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__32_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__32_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__32_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__32_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__32_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__32_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__32_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__32_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__32_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__32_ccff_tail[0])
  );


  cby_1__1_
  cby_3__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[130]),
    .prog_clk_0_W_in(prog_clk_0_wires[129]),
    .Test_en_E_in(Test_enWires[228]),
    .Test_en_W_out(Test_enWires[225]),
    .chany_bottom_in(sb_1__1__30_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__31_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_33_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__33_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__33_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__33_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__33_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__33_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__33_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__33_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__33_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__33_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__33_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__33_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__33_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__33_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__33_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__33_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__33_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__33_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__33_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__33_ccff_tail[0])
  );


  cby_1__1_
  cby_3__11_
  (
    .clk_2_N_out(clk_2_wires[65]),
    .clk_2_S_in(clk_2_wires[64]),
    .prog_clk_2_N_out(prog_clk_2_wires[65]),
    .prog_clk_2_S_in(prog_clk_2_wires[64]),
    .prog_clk_0_S_out(prog_clk_0_wires[133]),
    .prog_clk_0_W_in(prog_clk_0_wires[132]),
    .Test_en_E_in(Test_enWires[250]),
    .Test_en_W_out(Test_enWires[247]),
    .chany_bottom_in(sb_1__1__31_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__32_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_34_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__34_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__34_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__34_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__34_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__34_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__34_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__34_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__34_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__34_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__34_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__34_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__34_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__34_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__34_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__34_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__34_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__34_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__34_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__34_ccff_tail[0])
  );


  cby_1__1_
  cby_3__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[138]),
    .prog_clk_0_S_out(prog_clk_0_wires[136]),
    .prog_clk_0_W_in(prog_clk_0_wires[135]),
    .Test_en_E_in(Test_enWires[272]),
    .Test_en_W_out(Test_enWires[269]),
    .chany_bottom_in(sb_1__1__32_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_35_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__35_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__35_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__35_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__35_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__35_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__35_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__35_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__35_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__35_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__35_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__35_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__35_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__35_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__35_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__35_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__35_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__35_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__35_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__35_ccff_tail[0])
  );


  cby_1__1_
  cby_4__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[141]),
    .prog_clk_0_W_in(prog_clk_0_wires[140]),
    .Test_en_E_in(Test_enWires[32]),
    .Test_en_W_out(Test_enWires[29]),
    .chany_bottom_in(sb_1__0__3_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__33_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_36_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__36_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__36_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__36_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__36_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__36_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__36_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__36_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__36_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__36_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__36_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__36_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__36_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__36_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__36_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__36_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__36_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__36_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__36_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__36_ccff_tail[0])
  );


  cby_1__1_
  cby_4__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[144]),
    .prog_clk_0_W_in(prog_clk_0_wires[143]),
    .Test_en_E_in(Test_enWires[54]),
    .Test_en_W_out(Test_enWires[51]),
    .chany_bottom_in(sb_1__1__33_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__34_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_37_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__37_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__37_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__37_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__37_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__37_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__37_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__37_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__37_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__37_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__37_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__37_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__37_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__37_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__37_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__37_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__37_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__37_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__37_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__37_ccff_tail[0])
  );


  cby_1__1_
  cby_4__3_
  (
    .clk_3_S_out(clk_3_wires[25]),
    .clk_3_N_in(clk_3_wires[24]),
    .prog_clk_3_S_out(prog_clk_3_wires[25]),
    .prog_clk_3_N_in(prog_clk_3_wires[24]),
    .prog_clk_0_S_out(prog_clk_0_wires[147]),
    .prog_clk_0_W_in(prog_clk_0_wires[146]),
    .Test_en_E_in(Test_enWires[76]),
    .Test_en_W_out(Test_enWires[73]),
    .chany_bottom_in(sb_1__1__34_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__35_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_38_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__38_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__38_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__38_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__38_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__38_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__38_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__38_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__38_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__38_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__38_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__38_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__38_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__38_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__38_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__38_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__38_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__38_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__38_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__38_ccff_tail[0])
  );


  cby_1__1_
  cby_4__4_
  (
    .clk_3_S_out(clk_3_wires[21]),
    .clk_3_N_in(clk_3_wires[20]),
    .prog_clk_3_S_out(prog_clk_3_wires[21]),
    .prog_clk_3_N_in(prog_clk_3_wires[20]),
    .prog_clk_0_S_out(prog_clk_0_wires[150]),
    .prog_clk_0_W_in(prog_clk_0_wires[149]),
    .Test_en_E_in(Test_enWires[98]),
    .Test_en_W_out(Test_enWires[95]),
    .chany_bottom_in(sb_1__1__35_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__36_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_39_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__39_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__39_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__39_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__39_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__39_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__39_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__39_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__39_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__39_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__39_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__39_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__39_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__39_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__39_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__39_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__39_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__39_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__39_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__39_ccff_tail[0])
  );


  cby_1__1_
  cby_4__5_
  (
    .clk_3_S_out(clk_3_wires[15]),
    .clk_3_N_in(clk_3_wires[14]),
    .prog_clk_3_S_out(prog_clk_3_wires[15]),
    .prog_clk_3_N_in(prog_clk_3_wires[14]),
    .prog_clk_0_S_out(prog_clk_0_wires[153]),
    .prog_clk_0_W_in(prog_clk_0_wires[152]),
    .Test_en_E_in(Test_enWires[120]),
    .Test_en_W_out(Test_enWires[117]),
    .chany_bottom_in(sb_1__1__36_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__37_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_40_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__40_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__40_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__40_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__40_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__40_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__40_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__40_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__40_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__40_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__40_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__40_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__40_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__40_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__40_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__40_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__40_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__40_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__40_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__40_ccff_tail[0])
  );


  cby_1__1_
  cby_4__6_
  (
    .clk_3_S_out(clk_3_wires[11]),
    .clk_3_N_in(clk_3_wires[10]),
    .prog_clk_3_S_out(prog_clk_3_wires[11]),
    .prog_clk_3_N_in(prog_clk_3_wires[10]),
    .prog_clk_0_S_out(prog_clk_0_wires[156]),
    .prog_clk_0_W_in(prog_clk_0_wires[155]),
    .Test_en_E_in(Test_enWires[142]),
    .Test_en_W_out(Test_enWires[139]),
    .chany_bottom_in(sb_1__1__37_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__38_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_41_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__41_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__41_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__41_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__41_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__41_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__41_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__41_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__41_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__41_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__41_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__41_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__41_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__41_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__41_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__41_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__41_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__41_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__41_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__41_ccff_tail[0])
  );


  cby_1__1_
  cby_4__7_
  (
    .clk_3_N_out(clk_3_wires[9]),
    .clk_3_S_in(clk_3_wires[8]),
    .prog_clk_3_N_out(prog_clk_3_wires[9]),
    .prog_clk_3_S_in(prog_clk_3_wires[8]),
    .prog_clk_0_S_out(prog_clk_0_wires[159]),
    .prog_clk_0_W_in(prog_clk_0_wires[158]),
    .Test_en_E_in(Test_enWires[164]),
    .Test_en_W_out(Test_enWires[161]),
    .chany_bottom_in(sb_1__1__38_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__39_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_42_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__42_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__42_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__42_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__42_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__42_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__42_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__42_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__42_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__42_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__42_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__42_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__42_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__42_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__42_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__42_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__42_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__42_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__42_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__42_ccff_tail[0])
  );


  cby_1__1_
  cby_4__8_
  (
    .clk_3_N_out(clk_3_wires[13]),
    .clk_3_S_in(clk_3_wires[12]),
    .prog_clk_3_N_out(prog_clk_3_wires[13]),
    .prog_clk_3_S_in(prog_clk_3_wires[12]),
    .prog_clk_0_S_out(prog_clk_0_wires[162]),
    .prog_clk_0_W_in(prog_clk_0_wires[161]),
    .Test_en_E_in(Test_enWires[186]),
    .Test_en_W_out(Test_enWires[183]),
    .chany_bottom_in(sb_1__1__39_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__40_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_43_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__43_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__43_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__43_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__43_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__43_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__43_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__43_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__43_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__43_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__43_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__43_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__43_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__43_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__43_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__43_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__43_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__43_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__43_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__43_ccff_tail[0])
  );


  cby_1__1_
  cby_4__9_
  (
    .clk_3_N_out(clk_3_wires[19]),
    .clk_3_S_in(clk_3_wires[18]),
    .prog_clk_3_N_out(prog_clk_3_wires[19]),
    .prog_clk_3_S_in(prog_clk_3_wires[18]),
    .prog_clk_0_S_out(prog_clk_0_wires[165]),
    .prog_clk_0_W_in(prog_clk_0_wires[164]),
    .Test_en_E_in(Test_enWires[208]),
    .Test_en_W_out(Test_enWires[205]),
    .chany_bottom_in(sb_1__1__40_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__41_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_44_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__44_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__44_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__44_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__44_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__44_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__44_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__44_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__44_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__44_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__44_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__44_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__44_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__44_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__44_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__44_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__44_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__44_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__44_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__44_ccff_tail[0])
  );


  cby_1__1_
  cby_4__10_
  (
    .clk_3_N_out(clk_3_wires[23]),
    .clk_3_S_in(clk_3_wires[22]),
    .prog_clk_3_N_out(prog_clk_3_wires[23]),
    .prog_clk_3_S_in(prog_clk_3_wires[22]),
    .prog_clk_0_S_out(prog_clk_0_wires[168]),
    .prog_clk_0_W_in(prog_clk_0_wires[167]),
    .Test_en_E_in(Test_enWires[230]),
    .Test_en_W_out(Test_enWires[227]),
    .chany_bottom_in(sb_1__1__41_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__42_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_45_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__45_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__45_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__45_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__45_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__45_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__45_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__45_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__45_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__45_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__45_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__45_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__45_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__45_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__45_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__45_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__45_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__45_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__45_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__45_ccff_tail[0])
  );


  cby_1__1_
  cby_4__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[171]),
    .prog_clk_0_W_in(prog_clk_0_wires[170]),
    .Test_en_E_in(Test_enWires[252]),
    .Test_en_W_out(Test_enWires[249]),
    .chany_bottom_in(sb_1__1__42_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__43_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_46_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__46_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__46_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__46_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__46_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__46_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__46_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__46_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__46_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__46_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__46_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__46_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__46_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__46_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__46_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__46_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__46_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__46_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__46_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__46_ccff_tail[0])
  );


  cby_1__1_
  cby_4__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[176]),
    .prog_clk_0_S_out(prog_clk_0_wires[174]),
    .prog_clk_0_W_in(prog_clk_0_wires[173]),
    .Test_en_E_in(Test_enWires[274]),
    .Test_en_W_out(Test_enWires[271]),
    .chany_bottom_in(sb_1__1__43_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_47_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__47_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__47_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__47_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__47_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__47_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__47_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__47_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__47_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__47_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__47_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__47_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__47_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__47_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__47_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__47_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__47_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__47_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__47_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__47_ccff_tail[0])
  );


  cby_1__1_
  cby_5__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[179]),
    .prog_clk_0_W_in(prog_clk_0_wires[178]),
    .Test_en_E_in(Test_enWires[34]),
    .Test_en_W_out(Test_enWires[31]),
    .chany_bottom_in(sb_1__0__4_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__44_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_48_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__48_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__48_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__48_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__48_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__48_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__48_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__48_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__48_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__48_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__48_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__48_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__48_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__48_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__48_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__48_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__48_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__48_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__48_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__48_ccff_tail[0])
  );


  cby_1__1_
  cby_5__2_
  (
    .clk_2_S_out(clk_2_wires[32]),
    .clk_2_N_in(clk_2_wires[31]),
    .prog_clk_2_S_out(prog_clk_2_wires[32]),
    .prog_clk_2_N_in(prog_clk_2_wires[31]),
    .prog_clk_0_S_out(prog_clk_0_wires[182]),
    .prog_clk_0_W_in(prog_clk_0_wires[181]),
    .Test_en_E_in(Test_enWires[56]),
    .Test_en_W_out(Test_enWires[53]),
    .chany_bottom_in(sb_1__1__44_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__45_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_49_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__49_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__49_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__49_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__49_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__49_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__49_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__49_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__49_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__49_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__49_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__49_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__49_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__49_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__49_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__49_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__49_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__49_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__49_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__49_ccff_tail[0])
  );


  cby_1__1_
  cby_5__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[185]),
    .prog_clk_0_W_in(prog_clk_0_wires[184]),
    .Test_en_E_in(Test_enWires[78]),
    .Test_en_W_out(Test_enWires[75]),
    .chany_bottom_in(sb_1__1__45_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__46_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_50_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__50_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__50_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__50_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__50_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__50_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__50_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__50_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__50_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__50_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__50_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__50_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__50_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__50_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__50_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__50_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__50_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__50_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__50_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__50_ccff_tail[0])
  );


  cby_1__1_
  cby_5__4_
  (
    .clk_2_S_out(clk_2_wires[45]),
    .clk_2_N_in(clk_2_wires[44]),
    .prog_clk_2_S_out(prog_clk_2_wires[45]),
    .prog_clk_2_N_in(prog_clk_2_wires[44]),
    .prog_clk_0_S_out(prog_clk_0_wires[188]),
    .prog_clk_0_W_in(prog_clk_0_wires[187]),
    .Test_en_E_in(Test_enWires[100]),
    .Test_en_W_out(Test_enWires[97]),
    .chany_bottom_in(sb_1__1__46_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__47_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_51_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__51_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__51_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__51_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__51_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__51_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__51_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__51_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__51_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__51_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__51_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__51_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__51_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__51_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__51_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__51_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__51_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__51_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__51_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__51_ccff_tail[0])
  );


  cby_1__1_
  cby_5__5_
  (
    .clk_2_N_out(clk_2_wires[43]),
    .clk_2_S_in(clk_2_wires[42]),
    .prog_clk_2_N_out(prog_clk_2_wires[43]),
    .prog_clk_2_S_in(prog_clk_2_wires[42]),
    .prog_clk_0_S_out(prog_clk_0_wires[191]),
    .prog_clk_0_W_in(prog_clk_0_wires[190]),
    .Test_en_E_in(Test_enWires[122]),
    .Test_en_W_out(Test_enWires[119]),
    .chany_bottom_in(sb_1__1__47_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__48_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_52_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__52_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__52_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__52_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__52_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__52_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__52_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__52_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__52_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__52_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__52_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__52_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__52_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__52_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__52_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__52_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__52_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__52_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__52_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__52_ccff_tail[0])
  );


  cby_1__1_
  cby_5__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[194]),
    .prog_clk_0_W_in(prog_clk_0_wires[193]),
    .Test_en_E_in(Test_enWires[144]),
    .Test_en_W_out(Test_enWires[141]),
    .chany_bottom_in(sb_1__1__48_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__49_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_53_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__53_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__53_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__53_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__53_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__53_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__53_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__53_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__53_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__53_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__53_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__53_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__53_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__53_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__53_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__53_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__53_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__53_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__53_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__53_ccff_tail[0])
  );


  cby_1__1_
  cby_5__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[197]),
    .prog_clk_0_W_in(prog_clk_0_wires[196]),
    .Test_en_E_in(Test_enWires[166]),
    .Test_en_W_out(Test_enWires[163]),
    .chany_bottom_in(sb_1__1__49_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__50_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_54_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__54_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__54_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__54_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__54_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__54_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__54_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__54_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__54_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__54_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__54_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__54_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__54_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__54_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__54_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__54_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__54_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__54_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__54_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__54_ccff_tail[0])
  );


  cby_1__1_
  cby_5__8_
  (
    .clk_2_S_out(clk_2_wires[58]),
    .clk_2_N_in(clk_2_wires[57]),
    .prog_clk_2_S_out(prog_clk_2_wires[58]),
    .prog_clk_2_N_in(prog_clk_2_wires[57]),
    .prog_clk_0_S_out(prog_clk_0_wires[200]),
    .prog_clk_0_W_in(prog_clk_0_wires[199]),
    .Test_en_E_in(Test_enWires[188]),
    .Test_en_W_out(Test_enWires[185]),
    .chany_bottom_in(sb_1__1__50_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__51_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_55_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__55_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__55_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__55_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__55_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__55_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__55_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__55_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__55_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__55_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__55_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__55_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__55_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__55_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__55_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__55_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__55_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__55_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__55_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__55_ccff_tail[0])
  );


  cby_1__1_
  cby_5__9_
  (
    .clk_2_N_out(clk_2_wires[56]),
    .clk_2_S_in(clk_2_wires[55]),
    .prog_clk_2_N_out(prog_clk_2_wires[56]),
    .prog_clk_2_S_in(prog_clk_2_wires[55]),
    .prog_clk_0_S_out(prog_clk_0_wires[203]),
    .prog_clk_0_W_in(prog_clk_0_wires[202]),
    .Test_en_E_in(Test_enWires[210]),
    .Test_en_W_out(Test_enWires[207]),
    .chany_bottom_in(sb_1__1__51_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__52_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_56_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__56_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__56_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__56_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__56_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__56_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__56_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__56_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__56_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__56_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__56_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__56_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__56_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__56_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__56_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__56_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__56_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__56_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__56_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__56_ccff_tail[0])
  );


  cby_1__1_
  cby_5__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[206]),
    .prog_clk_0_W_in(prog_clk_0_wires[205]),
    .Test_en_E_in(Test_enWires[232]),
    .Test_en_W_out(Test_enWires[229]),
    .chany_bottom_in(sb_1__1__52_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__53_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_57_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__57_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__57_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__57_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__57_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__57_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__57_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__57_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__57_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__57_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__57_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__57_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__57_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__57_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__57_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__57_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__57_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__57_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__57_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__57_ccff_tail[0])
  );


  cby_1__1_
  cby_5__11_
  (
    .clk_2_N_out(clk_2_wires[67]),
    .clk_2_S_in(clk_2_wires[66]),
    .prog_clk_2_N_out(prog_clk_2_wires[67]),
    .prog_clk_2_S_in(prog_clk_2_wires[66]),
    .prog_clk_0_S_out(prog_clk_0_wires[209]),
    .prog_clk_0_W_in(prog_clk_0_wires[208]),
    .Test_en_E_in(Test_enWires[254]),
    .Test_en_W_out(Test_enWires[251]),
    .chany_bottom_in(sb_1__1__53_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__54_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_58_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__58_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__58_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__58_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__58_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__58_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__58_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__58_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__58_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__58_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__58_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__58_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__58_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__58_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__58_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__58_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__58_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__58_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__58_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__58_ccff_tail[0])
  );


  cby_1__1_
  cby_5__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[214]),
    .prog_clk_0_S_out(prog_clk_0_wires[212]),
    .prog_clk_0_W_in(prog_clk_0_wires[211]),
    .Test_en_E_in(Test_enWires[276]),
    .Test_en_W_out(Test_enWires[273]),
    .chany_bottom_in(sb_1__1__54_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_59_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__59_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__59_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__59_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__59_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__59_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__59_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__59_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__59_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__59_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__59_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__59_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__59_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__59_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__59_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__59_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__59_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__59_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__59_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__59_ccff_tail[0])
  );


  cby_1__1_
  cby_6__1_
  (
    .clk_3_S_in(clk_3_wires[90]),
    .clk_3_N_out(clk_3_wires[89]),
    .prog_clk_3_S_in(prog_clk_3_wires[90]),
    .prog_clk_3_N_out(prog_clk_3_wires[89]),
    .prog_clk_0_S_out(prog_clk_0_wires[217]),
    .prog_clk_0_W_in(prog_clk_0_wires[216]),
    .Test_en_E_out(Test_enWires[35]),
    .Test_en_W_out(Test_enWires[33]),
    .Test_en_N_out(Test_enWires[2]),
    .Test_en_S_in(Test_enWires[1]),
    .chany_bottom_in(sb_1__0__5_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__55_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_60_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__60_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__60_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__60_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__60_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__60_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__60_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__60_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__60_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__60_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__60_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__60_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__60_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__60_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__60_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__60_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__60_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__60_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__60_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__60_ccff_tail[0])
  );


  cby_1__1_
  cby_6__2_
  (
    .clk_3_S_in(clk_3_wires[92]),
    .clk_3_N_out(clk_3_wires[91]),
    .prog_clk_3_S_in(prog_clk_3_wires[92]),
    .prog_clk_3_N_out(prog_clk_3_wires[91]),
    .prog_clk_0_S_out(prog_clk_0_wires[220]),
    .prog_clk_0_W_in(prog_clk_0_wires[219]),
    .Test_en_E_out(Test_enWires[57]),
    .Test_en_W_out(Test_enWires[55]),
    .Test_en_N_out(Test_enWires[4]),
    .Test_en_S_in(Test_enWires[3]),
    .chany_bottom_in(sb_1__1__55_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__56_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_61_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__61_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__61_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__61_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__61_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__61_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__61_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__61_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__61_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__61_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__61_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__61_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__61_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__61_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__61_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__61_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__61_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__61_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__61_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__61_ccff_tail[0])
  );


  cby_1__1_
  cby_6__3_
  (
    .clk_3_S_in(clk_3_wires[94]),
    .clk_3_N_out(clk_3_wires[93]),
    .prog_clk_3_S_in(prog_clk_3_wires[94]),
    .prog_clk_3_N_out(prog_clk_3_wires[93]),
    .prog_clk_0_S_out(prog_clk_0_wires[223]),
    .prog_clk_0_W_in(prog_clk_0_wires[222]),
    .Test_en_E_out(Test_enWires[79]),
    .Test_en_W_out(Test_enWires[77]),
    .Test_en_N_out(Test_enWires[6]),
    .Test_en_S_in(Test_enWires[5]),
    .chany_bottom_in(sb_1__1__56_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__57_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_62_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__62_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__62_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__62_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__62_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__62_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__62_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__62_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__62_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__62_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__62_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__62_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__62_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__62_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__62_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__62_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__62_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__62_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__62_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__62_ccff_tail[0])
  );


  cby_1__1_
  cby_6__4_
  (
    .clk_3_S_in(clk_3_wires[96]),
    .clk_3_N_out(clk_3_wires[95]),
    .prog_clk_3_S_in(prog_clk_3_wires[96]),
    .prog_clk_3_N_out(prog_clk_3_wires[95]),
    .prog_clk_0_S_out(prog_clk_0_wires[226]),
    .prog_clk_0_W_in(prog_clk_0_wires[225]),
    .Test_en_E_out(Test_enWires[101]),
    .Test_en_W_out(Test_enWires[99]),
    .Test_en_N_out(Test_enWires[8]),
    .Test_en_S_in(Test_enWires[7]),
    .chany_bottom_in(sb_1__1__57_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__58_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_63_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__63_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__63_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__63_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__63_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__63_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__63_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__63_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__63_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__63_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__63_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__63_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__63_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__63_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__63_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__63_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__63_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__63_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__63_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__63_ccff_tail[0])
  );


  cby_1__1_
  cby_6__5_
  (
    .clk_3_S_in(clk_3_wires[98]),
    .clk_3_N_out(clk_3_wires[97]),
    .prog_clk_3_S_in(prog_clk_3_wires[98]),
    .prog_clk_3_N_out(prog_clk_3_wires[97]),
    .prog_clk_0_S_out(prog_clk_0_wires[229]),
    .prog_clk_0_W_in(prog_clk_0_wires[228]),
    .Test_en_E_out(Test_enWires[123]),
    .Test_en_W_out(Test_enWires[121]),
    .Test_en_N_out(Test_enWires[10]),
    .Test_en_S_in(Test_enWires[9]),
    .chany_bottom_in(sb_1__1__58_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__59_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_64_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__64_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__64_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__64_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__64_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__64_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__64_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__64_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__64_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__64_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__64_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__64_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__64_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__64_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__64_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__64_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__64_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__64_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__64_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__64_ccff_tail[0])
  );


  cby_1__1_
  cby_6__6_
  (
    .clk_3_S_in(clk_3_wires[100]),
    .clk_3_N_out(clk_3_wires[99]),
    .prog_clk_3_S_in(prog_clk_3_wires[100]),
    .prog_clk_3_N_out(prog_clk_3_wires[99]),
    .prog_clk_0_S_out(prog_clk_0_wires[232]),
    .prog_clk_0_W_in(prog_clk_0_wires[231]),
    .Test_en_E_out(Test_enWires[145]),
    .Test_en_W_out(Test_enWires[143]),
    .Test_en_N_out(Test_enWires[12]),
    .Test_en_S_in(Test_enWires[11]),
    .chany_bottom_in(sb_1__1__59_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__60_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_65_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__65_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__65_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__65_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__65_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__65_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__65_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__65_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__65_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__65_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__65_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__65_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__65_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__65_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__65_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__65_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__65_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__65_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__65_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__65_ccff_tail[0])
  );


  cby_1__1_
  cby_6__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[235]),
    .prog_clk_0_W_in(prog_clk_0_wires[234]),
    .Test_en_E_out(Test_enWires[167]),
    .Test_en_W_out(Test_enWires[165]),
    .Test_en_N_out(Test_enWires[14]),
    .Test_en_S_in(Test_enWires[13]),
    .chany_bottom_in(sb_1__1__60_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__61_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_66_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__66_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__66_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__66_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__66_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__66_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__66_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__66_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__66_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__66_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__66_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__66_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__66_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__66_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__66_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__66_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__66_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__66_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__66_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__66_ccff_tail[0])
  );


  cby_1__1_
  cby_6__8_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[238]),
    .prog_clk_0_W_in(prog_clk_0_wires[237]),
    .Test_en_E_out(Test_enWires[189]),
    .Test_en_W_out(Test_enWires[187]),
    .Test_en_N_out(Test_enWires[16]),
    .Test_en_S_in(Test_enWires[15]),
    .chany_bottom_in(sb_1__1__61_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__62_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_67_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__67_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__67_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__67_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__67_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__67_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__67_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__67_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__67_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__67_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__67_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__67_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__67_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__67_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__67_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__67_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__67_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__67_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__67_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__67_ccff_tail[0])
  );


  cby_1__1_
  cby_6__9_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[241]),
    .prog_clk_0_W_in(prog_clk_0_wires[240]),
    .Test_en_E_out(Test_enWires[211]),
    .Test_en_W_out(Test_enWires[209]),
    .Test_en_N_out(Test_enWires[18]),
    .Test_en_S_in(Test_enWires[17]),
    .chany_bottom_in(sb_1__1__62_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__63_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_68_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__68_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__68_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__68_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__68_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__68_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__68_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__68_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__68_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__68_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__68_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__68_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__68_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__68_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__68_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__68_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__68_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__68_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__68_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__68_ccff_tail[0])
  );


  cby_1__1_
  cby_6__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[244]),
    .prog_clk_0_W_in(prog_clk_0_wires[243]),
    .Test_en_E_out(Test_enWires[233]),
    .Test_en_W_out(Test_enWires[231]),
    .Test_en_N_out(Test_enWires[20]),
    .Test_en_S_in(Test_enWires[19]),
    .chany_bottom_in(sb_1__1__63_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__64_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_69_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__69_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__69_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__69_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__69_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__69_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__69_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__69_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__69_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__69_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__69_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__69_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__69_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__69_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__69_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__69_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__69_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__69_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__69_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__69_ccff_tail[0])
  );


  cby_1__1_
  cby_6__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[247]),
    .prog_clk_0_W_in(prog_clk_0_wires[246]),
    .Test_en_E_out(Test_enWires[255]),
    .Test_en_W_out(Test_enWires[253]),
    .Test_en_N_out(Test_enWires[22]),
    .Test_en_S_in(Test_enWires[21]),
    .chany_bottom_in(sb_1__1__64_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__65_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_70_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__70_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__70_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__70_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__70_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__70_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__70_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__70_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__70_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__70_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__70_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__70_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__70_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__70_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__70_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__70_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__70_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__70_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__70_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__70_ccff_tail[0])
  );


  cby_1__1_
  cby_6__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[252]),
    .prog_clk_0_S_out(prog_clk_0_wires[250]),
    .prog_clk_0_W_in(prog_clk_0_wires[249]),
    .Test_en_E_out(Test_enWires[277]),
    .Test_en_W_out(Test_enWires[275]),
    .Test_en_S_in(Test_enWires[23]),
    .chany_bottom_in(sb_1__1__65_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_71_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__71_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__71_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__71_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__71_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__71_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__71_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__71_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__71_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__71_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__71_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__71_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__71_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__71_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__71_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__71_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__71_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__71_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__71_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__71_ccff_tail[0])
  );


  cby_1__1_
  cby_7__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[255]),
    .prog_clk_0_W_in(prog_clk_0_wires[254]),
    .Test_en_E_out(Test_enWires[37]),
    .Test_en_W_in(Test_enWires[36]),
    .chany_bottom_in(sb_1__0__6_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__66_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_72_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__72_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__72_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__72_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__72_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__72_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__72_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__72_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__72_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__72_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__72_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__72_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__72_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__72_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__72_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__72_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__72_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__72_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__72_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__72_ccff_tail[0])
  );


  cby_1__1_
  cby_7__2_
  (
    .clk_2_S_out(clk_2_wires[74]),
    .clk_2_N_in(clk_2_wires[73]),
    .prog_clk_2_S_out(prog_clk_2_wires[74]),
    .prog_clk_2_N_in(prog_clk_2_wires[73]),
    .prog_clk_0_S_out(prog_clk_0_wires[258]),
    .prog_clk_0_W_in(prog_clk_0_wires[257]),
    .Test_en_E_out(Test_enWires[59]),
    .Test_en_W_in(Test_enWires[58]),
    .chany_bottom_in(sb_1__1__66_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__67_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_73_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__73_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__73_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__73_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__73_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__73_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__73_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__73_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__73_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__73_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__73_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__73_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__73_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__73_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__73_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__73_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__73_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__73_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__73_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__73_ccff_tail[0])
  );


  cby_1__1_
  cby_7__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[261]),
    .prog_clk_0_W_in(prog_clk_0_wires[260]),
    .Test_en_E_out(Test_enWires[81]),
    .Test_en_W_in(Test_enWires[80]),
    .chany_bottom_in(sb_1__1__67_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__68_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_74_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__74_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__74_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__74_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__74_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__74_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__74_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__74_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__74_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__74_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__74_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__74_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__74_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__74_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__74_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__74_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__74_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__74_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__74_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__74_ccff_tail[0])
  );


  cby_1__1_
  cby_7__4_
  (
    .clk_2_S_out(clk_2_wires[85]),
    .clk_2_N_in(clk_2_wires[84]),
    .prog_clk_2_S_out(prog_clk_2_wires[85]),
    .prog_clk_2_N_in(prog_clk_2_wires[84]),
    .prog_clk_0_S_out(prog_clk_0_wires[264]),
    .prog_clk_0_W_in(prog_clk_0_wires[263]),
    .Test_en_E_out(Test_enWires[103]),
    .Test_en_W_in(Test_enWires[102]),
    .chany_bottom_in(sb_1__1__68_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__69_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_75_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__75_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__75_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__75_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__75_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__75_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__75_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__75_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__75_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__75_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__75_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__75_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__75_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__75_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__75_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__75_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__75_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__75_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__75_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__75_ccff_tail[0])
  );


  cby_1__1_
  cby_7__5_
  (
    .clk_2_N_out(clk_2_wires[83]),
    .clk_2_S_in(clk_2_wires[82]),
    .prog_clk_2_N_out(prog_clk_2_wires[83]),
    .prog_clk_2_S_in(prog_clk_2_wires[82]),
    .prog_clk_0_S_out(prog_clk_0_wires[267]),
    .prog_clk_0_W_in(prog_clk_0_wires[266]),
    .Test_en_E_out(Test_enWires[125]),
    .Test_en_W_in(Test_enWires[124]),
    .chany_bottom_in(sb_1__1__69_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__70_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_76_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__76_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__76_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__76_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__76_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__76_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__76_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__76_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__76_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__76_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__76_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__76_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__76_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__76_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__76_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__76_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__76_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__76_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__76_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__76_ccff_tail[0])
  );


  cby_1__1_
  cby_7__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[270]),
    .prog_clk_0_W_in(prog_clk_0_wires[269]),
    .Test_en_E_out(Test_enWires[147]),
    .Test_en_W_in(Test_enWires[146]),
    .chany_bottom_in(sb_1__1__70_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__71_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_77_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__77_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__77_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__77_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__77_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__77_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__77_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__77_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__77_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__77_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__77_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__77_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__77_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__77_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__77_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__77_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__77_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__77_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__77_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__77_ccff_tail[0])
  );


  cby_1__1_
  cby_7__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[273]),
    .prog_clk_0_W_in(prog_clk_0_wires[272]),
    .Test_en_E_out(Test_enWires[169]),
    .Test_en_W_in(Test_enWires[168]),
    .chany_bottom_in(sb_1__1__71_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__72_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_78_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__78_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__78_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__78_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__78_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__78_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__78_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__78_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__78_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__78_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__78_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__78_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__78_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__78_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__78_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__78_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__78_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__78_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__78_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__78_ccff_tail[0])
  );


  cby_1__1_
  cby_7__8_
  (
    .clk_2_S_out(clk_2_wires[98]),
    .clk_2_N_in(clk_2_wires[97]),
    .prog_clk_2_S_out(prog_clk_2_wires[98]),
    .prog_clk_2_N_in(prog_clk_2_wires[97]),
    .prog_clk_0_S_out(prog_clk_0_wires[276]),
    .prog_clk_0_W_in(prog_clk_0_wires[275]),
    .Test_en_E_out(Test_enWires[191]),
    .Test_en_W_in(Test_enWires[190]),
    .chany_bottom_in(sb_1__1__72_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__73_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_79_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__79_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__79_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__79_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__79_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__79_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__79_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__79_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__79_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__79_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__79_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__79_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__79_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__79_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__79_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__79_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__79_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__79_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__79_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__79_ccff_tail[0])
  );


  cby_1__1_
  cby_7__9_
  (
    .clk_2_N_out(clk_2_wires[96]),
    .clk_2_S_in(clk_2_wires[95]),
    .prog_clk_2_N_out(prog_clk_2_wires[96]),
    .prog_clk_2_S_in(prog_clk_2_wires[95]),
    .prog_clk_0_S_out(prog_clk_0_wires[279]),
    .prog_clk_0_W_in(prog_clk_0_wires[278]),
    .Test_en_E_out(Test_enWires[213]),
    .Test_en_W_in(Test_enWires[212]),
    .chany_bottom_in(sb_1__1__73_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__74_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_80_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__80_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__80_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__80_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__80_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__80_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__80_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__80_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__80_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__80_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__80_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__80_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__80_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__80_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__80_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__80_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__80_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__80_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__80_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__80_ccff_tail[0])
  );


  cby_1__1_
  cby_7__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[282]),
    .prog_clk_0_W_in(prog_clk_0_wires[281]),
    .Test_en_E_out(Test_enWires[235]),
    .Test_en_W_in(Test_enWires[234]),
    .chany_bottom_in(sb_1__1__74_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__75_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_81_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__81_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__81_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__81_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__81_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__81_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__81_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__81_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__81_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__81_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__81_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__81_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__81_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__81_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__81_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__81_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__81_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__81_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__81_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__81_ccff_tail[0])
  );


  cby_1__1_
  cby_7__11_
  (
    .clk_2_N_out(clk_2_wires[109]),
    .clk_2_S_in(clk_2_wires[108]),
    .prog_clk_2_N_out(prog_clk_2_wires[109]),
    .prog_clk_2_S_in(prog_clk_2_wires[108]),
    .prog_clk_0_S_out(prog_clk_0_wires[285]),
    .prog_clk_0_W_in(prog_clk_0_wires[284]),
    .Test_en_E_out(Test_enWires[257]),
    .Test_en_W_in(Test_enWires[256]),
    .chany_bottom_in(sb_1__1__75_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__76_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_82_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__82_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__82_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__82_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__82_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__82_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__82_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__82_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__82_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__82_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__82_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__82_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__82_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__82_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__82_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__82_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__82_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__82_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__82_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__82_ccff_tail[0])
  );


  cby_1__1_
  cby_7__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[290]),
    .prog_clk_0_S_out(prog_clk_0_wires[288]),
    .prog_clk_0_W_in(prog_clk_0_wires[287]),
    .Test_en_E_out(Test_enWires[279]),
    .Test_en_W_in(Test_enWires[278]),
    .chany_bottom_in(sb_1__1__76_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_83_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__83_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__83_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__83_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__83_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__83_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__83_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__83_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__83_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__83_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__83_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__83_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__83_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__83_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__83_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__83_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__83_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__83_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__83_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__83_ccff_tail[0])
  );


  cby_1__1_
  cby_8__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[293]),
    .prog_clk_0_W_in(prog_clk_0_wires[292]),
    .Test_en_E_out(Test_enWires[39]),
    .Test_en_W_in(Test_enWires[38]),
    .chany_bottom_in(sb_1__0__7_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__77_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_84_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__84_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__84_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__84_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__84_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__84_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__84_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__84_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__84_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__84_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__84_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__84_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__84_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__84_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__84_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__84_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__84_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__84_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__84_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__84_ccff_tail[0])
  );


  cby_1__1_
  cby_8__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[296]),
    .prog_clk_0_W_in(prog_clk_0_wires[295]),
    .Test_en_E_out(Test_enWires[61]),
    .Test_en_W_in(Test_enWires[60]),
    .chany_bottom_in(sb_1__1__77_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__78_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_85_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__85_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__85_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__85_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__85_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__85_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__85_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__85_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__85_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__85_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__85_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__85_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__85_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__85_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__85_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__85_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__85_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__85_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__85_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__85_ccff_tail[0])
  );


  cby_1__1_
  cby_8__3_
  (
    .clk_3_S_out(clk_3_wires[43]),
    .clk_3_N_in(clk_3_wires[42]),
    .prog_clk_3_S_out(prog_clk_3_wires[43]),
    .prog_clk_3_N_in(prog_clk_3_wires[42]),
    .prog_clk_0_S_out(prog_clk_0_wires[299]),
    .prog_clk_0_W_in(prog_clk_0_wires[298]),
    .Test_en_E_out(Test_enWires[83]),
    .Test_en_W_in(Test_enWires[82]),
    .chany_bottom_in(sb_1__1__78_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__79_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_86_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__86_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__86_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__86_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__86_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__86_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__86_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__86_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__86_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__86_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__86_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__86_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__86_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__86_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__86_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__86_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__86_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__86_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__86_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__86_ccff_tail[0])
  );


  cby_1__1_
  cby_8__4_
  (
    .clk_3_S_out(clk_3_wires[39]),
    .clk_3_N_in(clk_3_wires[38]),
    .prog_clk_3_S_out(prog_clk_3_wires[39]),
    .prog_clk_3_N_in(prog_clk_3_wires[38]),
    .prog_clk_0_S_out(prog_clk_0_wires[302]),
    .prog_clk_0_W_in(prog_clk_0_wires[301]),
    .Test_en_E_out(Test_enWires[105]),
    .Test_en_W_in(Test_enWires[104]),
    .chany_bottom_in(sb_1__1__79_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__80_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_87_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__87_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__87_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__87_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__87_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__87_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__87_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__87_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__87_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__87_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__87_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__87_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__87_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__87_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__87_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__87_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__87_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__87_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__87_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__87_ccff_tail[0])
  );


  cby_1__1_
  cby_8__5_
  (
    .clk_3_S_out(clk_3_wires[33]),
    .clk_3_N_in(clk_3_wires[32]),
    .prog_clk_3_S_out(prog_clk_3_wires[33]),
    .prog_clk_3_N_in(prog_clk_3_wires[32]),
    .prog_clk_0_S_out(prog_clk_0_wires[305]),
    .prog_clk_0_W_in(prog_clk_0_wires[304]),
    .Test_en_E_out(Test_enWires[127]),
    .Test_en_W_in(Test_enWires[126]),
    .chany_bottom_in(sb_1__1__80_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__81_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_88_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__88_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__88_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__88_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__88_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__88_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__88_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__88_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__88_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__88_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__88_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__88_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__88_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__88_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__88_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__88_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__88_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__88_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__88_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__88_ccff_tail[0])
  );


  cby_1__1_
  cby_8__6_
  (
    .clk_3_S_out(clk_3_wires[29]),
    .clk_3_N_in(clk_3_wires[28]),
    .prog_clk_3_S_out(prog_clk_3_wires[29]),
    .prog_clk_3_N_in(prog_clk_3_wires[28]),
    .prog_clk_0_S_out(prog_clk_0_wires[308]),
    .prog_clk_0_W_in(prog_clk_0_wires[307]),
    .Test_en_E_out(Test_enWires[149]),
    .Test_en_W_in(Test_enWires[148]),
    .chany_bottom_in(sb_1__1__81_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__82_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_89_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__89_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__89_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__89_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__89_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__89_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__89_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__89_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__89_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__89_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__89_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__89_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__89_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__89_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__89_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__89_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__89_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__89_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__89_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__89_ccff_tail[0])
  );


  cby_1__1_
  cby_8__7_
  (
    .clk_3_N_out(clk_3_wires[27]),
    .clk_3_S_in(clk_3_wires[26]),
    .prog_clk_3_N_out(prog_clk_3_wires[27]),
    .prog_clk_3_S_in(prog_clk_3_wires[26]),
    .prog_clk_0_S_out(prog_clk_0_wires[311]),
    .prog_clk_0_W_in(prog_clk_0_wires[310]),
    .Test_en_E_out(Test_enWires[171]),
    .Test_en_W_in(Test_enWires[170]),
    .chany_bottom_in(sb_1__1__82_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__83_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_90_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__90_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__90_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__90_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__90_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__90_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__90_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__90_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__90_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__90_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__90_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__90_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__90_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__90_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__90_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__90_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__90_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__90_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__90_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__90_ccff_tail[0])
  );


  cby_1__1_
  cby_8__8_
  (
    .clk_3_N_out(clk_3_wires[31]),
    .clk_3_S_in(clk_3_wires[30]),
    .prog_clk_3_N_out(prog_clk_3_wires[31]),
    .prog_clk_3_S_in(prog_clk_3_wires[30]),
    .prog_clk_0_S_out(prog_clk_0_wires[314]),
    .prog_clk_0_W_in(prog_clk_0_wires[313]),
    .Test_en_E_out(Test_enWires[193]),
    .Test_en_W_in(Test_enWires[192]),
    .chany_bottom_in(sb_1__1__83_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__84_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_91_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__91_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__91_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__91_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__91_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__91_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__91_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__91_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__91_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__91_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__91_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__91_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__91_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__91_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__91_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__91_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__91_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__91_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__91_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__91_ccff_tail[0])
  );


  cby_1__1_
  cby_8__9_
  (
    .clk_3_N_out(clk_3_wires[37]),
    .clk_3_S_in(clk_3_wires[36]),
    .prog_clk_3_N_out(prog_clk_3_wires[37]),
    .prog_clk_3_S_in(prog_clk_3_wires[36]),
    .prog_clk_0_S_out(prog_clk_0_wires[317]),
    .prog_clk_0_W_in(prog_clk_0_wires[316]),
    .Test_en_E_out(Test_enWires[215]),
    .Test_en_W_in(Test_enWires[214]),
    .chany_bottom_in(sb_1__1__84_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__85_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_92_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__92_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__92_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__92_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__92_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__92_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__92_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__92_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__92_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__92_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__92_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__92_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__92_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__92_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__92_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__92_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__92_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__92_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__92_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__92_ccff_tail[0])
  );


  cby_1__1_
  cby_8__10_
  (
    .clk_3_N_out(clk_3_wires[41]),
    .clk_3_S_in(clk_3_wires[40]),
    .prog_clk_3_N_out(prog_clk_3_wires[41]),
    .prog_clk_3_S_in(prog_clk_3_wires[40]),
    .prog_clk_0_S_out(prog_clk_0_wires[320]),
    .prog_clk_0_W_in(prog_clk_0_wires[319]),
    .Test_en_E_out(Test_enWires[237]),
    .Test_en_W_in(Test_enWires[236]),
    .chany_bottom_in(sb_1__1__85_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__86_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_93_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__93_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__93_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__93_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__93_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__93_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__93_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__93_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__93_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__93_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__93_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__93_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__93_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__93_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__93_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__93_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__93_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__93_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__93_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__93_ccff_tail[0])
  );


  cby_1__1_
  cby_8__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[323]),
    .prog_clk_0_W_in(prog_clk_0_wires[322]),
    .Test_en_E_out(Test_enWires[259]),
    .Test_en_W_in(Test_enWires[258]),
    .chany_bottom_in(sb_1__1__86_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__87_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_94_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__94_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__94_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__94_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__94_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__94_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__94_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__94_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__94_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__94_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__94_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__94_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__94_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__94_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__94_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__94_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__94_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__94_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__94_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__94_ccff_tail[0])
  );


  cby_1__1_
  cby_8__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[328]),
    .prog_clk_0_S_out(prog_clk_0_wires[326]),
    .prog_clk_0_W_in(prog_clk_0_wires[325]),
    .Test_en_E_out(Test_enWires[281]),
    .Test_en_W_in(Test_enWires[280]),
    .chany_bottom_in(sb_1__1__87_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__7_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_95_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__95_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__95_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__95_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__95_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__95_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__95_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__95_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__95_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__95_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__95_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__95_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__95_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__95_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__95_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__95_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__95_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__95_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__95_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__95_ccff_tail[0])
  );


  cby_1__1_
  cby_9__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[331]),
    .prog_clk_0_W_in(prog_clk_0_wires[330]),
    .Test_en_E_out(Test_enWires[41]),
    .Test_en_W_in(Test_enWires[40]),
    .chany_bottom_in(sb_1__0__8_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__88_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_96_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__96_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__96_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__96_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__96_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__96_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__96_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__96_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__96_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__96_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__96_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__96_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__96_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__96_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__96_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__96_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__96_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__96_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__96_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__96_ccff_tail[0])
  );


  cby_1__1_
  cby_9__2_
  (
    .clk_2_S_out(clk_2_wires[76]),
    .clk_2_N_in(clk_2_wires[75]),
    .prog_clk_2_S_out(prog_clk_2_wires[76]),
    .prog_clk_2_N_in(prog_clk_2_wires[75]),
    .prog_clk_0_S_out(prog_clk_0_wires[334]),
    .prog_clk_0_W_in(prog_clk_0_wires[333]),
    .Test_en_E_out(Test_enWires[63]),
    .Test_en_W_in(Test_enWires[62]),
    .chany_bottom_in(sb_1__1__88_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__89_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_97_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__97_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__97_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__97_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__97_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__97_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__97_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__97_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__97_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__97_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__97_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__97_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__97_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__97_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__97_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__97_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__97_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__97_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__97_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__97_ccff_tail[0])
  );


  cby_1__1_
  cby_9__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[337]),
    .prog_clk_0_W_in(prog_clk_0_wires[336]),
    .Test_en_E_out(Test_enWires[85]),
    .Test_en_W_in(Test_enWires[84]),
    .chany_bottom_in(sb_1__1__89_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__90_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_98_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__98_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__98_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__98_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__98_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__98_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__98_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__98_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__98_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__98_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__98_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__98_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__98_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__98_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__98_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__98_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__98_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__98_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__98_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__98_ccff_tail[0])
  );


  cby_1__1_
  cby_9__4_
  (
    .clk_2_S_out(clk_2_wires[89]),
    .clk_2_N_in(clk_2_wires[88]),
    .prog_clk_2_S_out(prog_clk_2_wires[89]),
    .prog_clk_2_N_in(prog_clk_2_wires[88]),
    .prog_clk_0_S_out(prog_clk_0_wires[340]),
    .prog_clk_0_W_in(prog_clk_0_wires[339]),
    .Test_en_E_out(Test_enWires[107]),
    .Test_en_W_in(Test_enWires[106]),
    .chany_bottom_in(sb_1__1__90_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__91_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_99_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__99_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__99_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__99_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__99_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__99_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__99_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__99_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__99_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__99_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__99_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__99_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__99_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__99_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__99_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__99_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__99_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__99_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__99_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__99_ccff_tail[0])
  );


  cby_1__1_
  cby_9__5_
  (
    .clk_2_N_out(clk_2_wires[87]),
    .clk_2_S_in(clk_2_wires[86]),
    .prog_clk_2_N_out(prog_clk_2_wires[87]),
    .prog_clk_2_S_in(prog_clk_2_wires[86]),
    .prog_clk_0_S_out(prog_clk_0_wires[343]),
    .prog_clk_0_W_in(prog_clk_0_wires[342]),
    .Test_en_E_out(Test_enWires[129]),
    .Test_en_W_in(Test_enWires[128]),
    .chany_bottom_in(sb_1__1__91_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__92_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_100_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__100_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__100_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__100_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__100_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__100_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__100_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__100_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__100_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__100_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__100_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__100_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__100_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__100_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__100_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__100_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__100_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__100_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__100_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__100_ccff_tail[0])
  );


  cby_1__1_
  cby_9__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[346]),
    .prog_clk_0_W_in(prog_clk_0_wires[345]),
    .Test_en_E_out(Test_enWires[151]),
    .Test_en_W_in(Test_enWires[150]),
    .chany_bottom_in(sb_1__1__92_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__93_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_101_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__101_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__101_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__101_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__101_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__101_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__101_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__101_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__101_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__101_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__101_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__101_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__101_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__101_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__101_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__101_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__101_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__101_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__101_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__101_ccff_tail[0])
  );


  cby_1__1_
  cby_9__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[349]),
    .prog_clk_0_W_in(prog_clk_0_wires[348]),
    .Test_en_E_out(Test_enWires[173]),
    .Test_en_W_in(Test_enWires[172]),
    .chany_bottom_in(sb_1__1__93_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__94_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_102_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__102_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__102_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__102_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__102_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__102_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__102_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__102_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__102_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__102_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__102_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__102_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__102_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__102_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__102_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__102_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__102_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__102_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__102_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__102_ccff_tail[0])
  );


  cby_1__1_
  cby_9__8_
  (
    .clk_2_S_out(clk_2_wires[102]),
    .clk_2_N_in(clk_2_wires[101]),
    .prog_clk_2_S_out(prog_clk_2_wires[102]),
    .prog_clk_2_N_in(prog_clk_2_wires[101]),
    .prog_clk_0_S_out(prog_clk_0_wires[352]),
    .prog_clk_0_W_in(prog_clk_0_wires[351]),
    .Test_en_E_out(Test_enWires[195]),
    .Test_en_W_in(Test_enWires[194]),
    .chany_bottom_in(sb_1__1__94_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__95_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_103_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__103_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__103_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__103_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__103_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__103_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__103_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__103_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__103_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__103_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__103_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__103_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__103_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__103_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__103_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__103_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__103_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__103_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__103_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__103_ccff_tail[0])
  );


  cby_1__1_
  cby_9__9_
  (
    .clk_2_N_out(clk_2_wires[100]),
    .clk_2_S_in(clk_2_wires[99]),
    .prog_clk_2_N_out(prog_clk_2_wires[100]),
    .prog_clk_2_S_in(prog_clk_2_wires[99]),
    .prog_clk_0_S_out(prog_clk_0_wires[355]),
    .prog_clk_0_W_in(prog_clk_0_wires[354]),
    .Test_en_E_out(Test_enWires[217]),
    .Test_en_W_in(Test_enWires[216]),
    .chany_bottom_in(sb_1__1__95_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__96_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_104_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__104_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__104_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__104_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__104_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__104_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__104_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__104_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__104_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__104_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__104_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__104_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__104_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__104_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__104_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__104_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__104_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__104_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__104_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__104_ccff_tail[0])
  );


  cby_1__1_
  cby_9__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[358]),
    .prog_clk_0_W_in(prog_clk_0_wires[357]),
    .Test_en_E_out(Test_enWires[239]),
    .Test_en_W_in(Test_enWires[238]),
    .chany_bottom_in(sb_1__1__96_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__97_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_105_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__105_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__105_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__105_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__105_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__105_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__105_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__105_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__105_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__105_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__105_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__105_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__105_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__105_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__105_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__105_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__105_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__105_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__105_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__105_ccff_tail[0])
  );


  cby_1__1_
  cby_9__11_
  (
    .clk_2_N_out(clk_2_wires[111]),
    .clk_2_S_in(clk_2_wires[110]),
    .prog_clk_2_N_out(prog_clk_2_wires[111]),
    .prog_clk_2_S_in(prog_clk_2_wires[110]),
    .prog_clk_0_S_out(prog_clk_0_wires[361]),
    .prog_clk_0_W_in(prog_clk_0_wires[360]),
    .Test_en_E_out(Test_enWires[261]),
    .Test_en_W_in(Test_enWires[260]),
    .chany_bottom_in(sb_1__1__97_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__98_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_106_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__106_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__106_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__106_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__106_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__106_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__106_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__106_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__106_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__106_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__106_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__106_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__106_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__106_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__106_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__106_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__106_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__106_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__106_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__106_ccff_tail[0])
  );


  cby_1__1_
  cby_9__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[366]),
    .prog_clk_0_S_out(prog_clk_0_wires[364]),
    .prog_clk_0_W_in(prog_clk_0_wires[363]),
    .Test_en_E_out(Test_enWires[283]),
    .Test_en_W_in(Test_enWires[282]),
    .chany_bottom_in(sb_1__1__98_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__8_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_107_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__107_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__107_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__107_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__107_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__107_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__107_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__107_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__107_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__107_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__107_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__107_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__107_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__107_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__107_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__107_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__107_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__107_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__107_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__107_ccff_tail[0])
  );


  cby_1__1_
  cby_10__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[369]),
    .prog_clk_0_W_in(prog_clk_0_wires[368]),
    .Test_en_E_out(Test_enWires[43]),
    .Test_en_W_in(Test_enWires[42]),
    .chany_bottom_in(sb_1__0__9_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__99_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_108_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__108_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__108_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__108_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__108_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__108_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__108_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__108_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__108_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__108_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__108_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__108_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__108_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__108_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__108_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__108_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__108_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__108_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__108_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__108_ccff_tail[0])
  );


  cby_1__1_
  cby_10__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[372]),
    .prog_clk_0_W_in(prog_clk_0_wires[371]),
    .Test_en_E_out(Test_enWires[65]),
    .Test_en_W_in(Test_enWires[64]),
    .chany_bottom_in(sb_1__1__99_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__100_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_109_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__109_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__109_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__109_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__109_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__109_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__109_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__109_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__109_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__109_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__109_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__109_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__109_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__109_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__109_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__109_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__109_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__109_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__109_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__109_ccff_tail[0])
  );


  cby_1__1_
  cby_10__3_
  (
    .clk_3_S_out(clk_3_wires[87]),
    .clk_3_N_in(clk_3_wires[86]),
    .prog_clk_3_S_out(prog_clk_3_wires[87]),
    .prog_clk_3_N_in(prog_clk_3_wires[86]),
    .prog_clk_0_S_out(prog_clk_0_wires[375]),
    .prog_clk_0_W_in(prog_clk_0_wires[374]),
    .Test_en_E_out(Test_enWires[87]),
    .Test_en_W_in(Test_enWires[86]),
    .chany_bottom_in(sb_1__1__100_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__101_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_110_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__110_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__110_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__110_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__110_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__110_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__110_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__110_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__110_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__110_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__110_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__110_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__110_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__110_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__110_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__110_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__110_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__110_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__110_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__110_ccff_tail[0])
  );


  cby_1__1_
  cby_10__4_
  (
    .clk_3_S_out(clk_3_wires[83]),
    .clk_3_N_in(clk_3_wires[82]),
    .prog_clk_3_S_out(prog_clk_3_wires[83]),
    .prog_clk_3_N_in(prog_clk_3_wires[82]),
    .prog_clk_0_S_out(prog_clk_0_wires[378]),
    .prog_clk_0_W_in(prog_clk_0_wires[377]),
    .Test_en_E_out(Test_enWires[109]),
    .Test_en_W_in(Test_enWires[108]),
    .chany_bottom_in(sb_1__1__101_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__102_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_111_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__111_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__111_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__111_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__111_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__111_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__111_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__111_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__111_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__111_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__111_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__111_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__111_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__111_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__111_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__111_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__111_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__111_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__111_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__111_ccff_tail[0])
  );


  cby_1__1_
  cby_10__5_
  (
    .clk_3_S_out(clk_3_wires[77]),
    .clk_3_N_in(clk_3_wires[76]),
    .prog_clk_3_S_out(prog_clk_3_wires[77]),
    .prog_clk_3_N_in(prog_clk_3_wires[76]),
    .prog_clk_0_S_out(prog_clk_0_wires[381]),
    .prog_clk_0_W_in(prog_clk_0_wires[380]),
    .Test_en_E_out(Test_enWires[131]),
    .Test_en_W_in(Test_enWires[130]),
    .chany_bottom_in(sb_1__1__102_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__103_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_112_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__112_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__112_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__112_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__112_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__112_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__112_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__112_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__112_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__112_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__112_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__112_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__112_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__112_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__112_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__112_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__112_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__112_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__112_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__112_ccff_tail[0])
  );


  cby_1__1_
  cby_10__6_
  (
    .clk_3_S_out(clk_3_wires[73]),
    .clk_3_N_in(clk_3_wires[72]),
    .prog_clk_3_S_out(prog_clk_3_wires[73]),
    .prog_clk_3_N_in(prog_clk_3_wires[72]),
    .prog_clk_0_S_out(prog_clk_0_wires[384]),
    .prog_clk_0_W_in(prog_clk_0_wires[383]),
    .Test_en_E_out(Test_enWires[153]),
    .Test_en_W_in(Test_enWires[152]),
    .chany_bottom_in(sb_1__1__103_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__104_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_113_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__113_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__113_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__113_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__113_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__113_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__113_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__113_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__113_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__113_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__113_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__113_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__113_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__113_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__113_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__113_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__113_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__113_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__113_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__113_ccff_tail[0])
  );


  cby_1__1_
  cby_10__7_
  (
    .clk_3_N_out(clk_3_wires[71]),
    .clk_3_S_in(clk_3_wires[70]),
    .prog_clk_3_N_out(prog_clk_3_wires[71]),
    .prog_clk_3_S_in(prog_clk_3_wires[70]),
    .prog_clk_0_S_out(prog_clk_0_wires[387]),
    .prog_clk_0_W_in(prog_clk_0_wires[386]),
    .Test_en_E_out(Test_enWires[175]),
    .Test_en_W_in(Test_enWires[174]),
    .chany_bottom_in(sb_1__1__104_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__105_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_114_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__114_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__114_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__114_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__114_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__114_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__114_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__114_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__114_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__114_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__114_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__114_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__114_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__114_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__114_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__114_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__114_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__114_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__114_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__114_ccff_tail[0])
  );


  cby_1__1_
  cby_10__8_
  (
    .clk_3_N_out(clk_3_wires[75]),
    .clk_3_S_in(clk_3_wires[74]),
    .prog_clk_3_N_out(prog_clk_3_wires[75]),
    .prog_clk_3_S_in(prog_clk_3_wires[74]),
    .prog_clk_0_S_out(prog_clk_0_wires[390]),
    .prog_clk_0_W_in(prog_clk_0_wires[389]),
    .Test_en_E_out(Test_enWires[197]),
    .Test_en_W_in(Test_enWires[196]),
    .chany_bottom_in(sb_1__1__105_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__106_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_115_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__115_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__115_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__115_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__115_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__115_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__115_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__115_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__115_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__115_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__115_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__115_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__115_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__115_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__115_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__115_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__115_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__115_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__115_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__115_ccff_tail[0])
  );


  cby_1__1_
  cby_10__9_
  (
    .clk_3_N_out(clk_3_wires[81]),
    .clk_3_S_in(clk_3_wires[80]),
    .prog_clk_3_N_out(prog_clk_3_wires[81]),
    .prog_clk_3_S_in(prog_clk_3_wires[80]),
    .prog_clk_0_S_out(prog_clk_0_wires[393]),
    .prog_clk_0_W_in(prog_clk_0_wires[392]),
    .Test_en_E_out(Test_enWires[219]),
    .Test_en_W_in(Test_enWires[218]),
    .chany_bottom_in(sb_1__1__106_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__107_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_116_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__116_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__116_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__116_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__116_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__116_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__116_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__116_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__116_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__116_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__116_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__116_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__116_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__116_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__116_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__116_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__116_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__116_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__116_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__116_ccff_tail[0])
  );


  cby_1__1_
  cby_10__10_
  (
    .clk_3_N_out(clk_3_wires[85]),
    .clk_3_S_in(clk_3_wires[84]),
    .prog_clk_3_N_out(prog_clk_3_wires[85]),
    .prog_clk_3_S_in(prog_clk_3_wires[84]),
    .prog_clk_0_S_out(prog_clk_0_wires[396]),
    .prog_clk_0_W_in(prog_clk_0_wires[395]),
    .Test_en_E_out(Test_enWires[241]),
    .Test_en_W_in(Test_enWires[240]),
    .chany_bottom_in(sb_1__1__107_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__108_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_117_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__117_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__117_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__117_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__117_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__117_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__117_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__117_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__117_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__117_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__117_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__117_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__117_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__117_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__117_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__117_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__117_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__117_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__117_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__117_ccff_tail[0])
  );


  cby_1__1_
  cby_10__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[399]),
    .prog_clk_0_W_in(prog_clk_0_wires[398]),
    .Test_en_E_out(Test_enWires[263]),
    .Test_en_W_in(Test_enWires[262]),
    .chany_bottom_in(sb_1__1__108_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__109_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_118_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__118_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__118_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__118_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__118_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__118_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__118_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__118_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__118_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__118_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__118_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__118_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__118_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__118_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__118_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__118_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__118_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__118_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__118_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__118_ccff_tail[0])
  );


  cby_1__1_
  cby_10__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[404]),
    .prog_clk_0_S_out(prog_clk_0_wires[402]),
    .prog_clk_0_W_in(prog_clk_0_wires[401]),
    .Test_en_E_out(Test_enWires[285]),
    .Test_en_W_in(Test_enWires[284]),
    .chany_bottom_in(sb_1__1__109_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__9_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_119_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__119_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__119_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__119_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__119_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__119_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__119_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__119_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__119_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__119_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__119_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__119_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__119_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__119_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__119_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__119_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__119_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__119_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__119_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__119_ccff_tail[0])
  );


  cby_1__1_
  cby_11__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[407]),
    .prog_clk_0_W_in(prog_clk_0_wires[406]),
    .Test_en_E_out(Test_enWires[45]),
    .Test_en_W_in(Test_enWires[44]),
    .chany_bottom_in(sb_1__0__10_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__110_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_120_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__120_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__120_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__120_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__120_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__120_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__120_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__120_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__120_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__120_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__120_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__120_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__120_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__120_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__120_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__120_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__120_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__120_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__120_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__120_ccff_tail[0])
  );


  cby_1__1_
  cby_11__2_
  (
    .clk_2_S_out(clk_2_wires[116]),
    .clk_2_N_in(clk_2_wires[115]),
    .prog_clk_2_S_out(prog_clk_2_wires[116]),
    .prog_clk_2_N_in(prog_clk_2_wires[115]),
    .prog_clk_0_S_out(prog_clk_0_wires[410]),
    .prog_clk_0_W_in(prog_clk_0_wires[409]),
    .Test_en_E_out(Test_enWires[67]),
    .Test_en_W_in(Test_enWires[66]),
    .chany_bottom_in(sb_1__1__110_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__111_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_121_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__121_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__121_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__121_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__121_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__121_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__121_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__121_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__121_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__121_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__121_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__121_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__121_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__121_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__121_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__121_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__121_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__121_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__121_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__121_ccff_tail[0])
  );


  cby_1__1_
  cby_11__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[413]),
    .prog_clk_0_W_in(prog_clk_0_wires[412]),
    .Test_en_E_out(Test_enWires[89]),
    .Test_en_W_in(Test_enWires[88]),
    .chany_bottom_in(sb_1__1__111_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__112_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_122_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__122_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__122_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__122_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__122_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__122_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__122_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__122_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__122_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__122_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__122_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__122_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__122_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__122_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__122_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__122_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__122_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__122_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__122_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__122_ccff_tail[0])
  );


  cby_1__1_
  cby_11__4_
  (
    .clk_2_S_out(clk_2_wires[123]),
    .clk_2_N_in(clk_2_wires[122]),
    .prog_clk_2_S_out(prog_clk_2_wires[123]),
    .prog_clk_2_N_in(prog_clk_2_wires[122]),
    .prog_clk_0_S_out(prog_clk_0_wires[416]),
    .prog_clk_0_W_in(prog_clk_0_wires[415]),
    .Test_en_E_out(Test_enWires[111]),
    .Test_en_W_in(Test_enWires[110]),
    .chany_bottom_in(sb_1__1__112_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__113_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_123_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__123_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__123_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__123_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__123_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__123_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__123_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__123_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__123_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__123_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__123_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__123_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__123_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__123_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__123_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__123_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__123_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__123_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__123_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__123_ccff_tail[0])
  );


  cby_1__1_
  cby_11__5_
  (
    .clk_2_N_out(clk_2_wires[121]),
    .clk_2_S_in(clk_2_wires[120]),
    .prog_clk_2_N_out(prog_clk_2_wires[121]),
    .prog_clk_2_S_in(prog_clk_2_wires[120]),
    .prog_clk_0_S_out(prog_clk_0_wires[419]),
    .prog_clk_0_W_in(prog_clk_0_wires[418]),
    .Test_en_E_out(Test_enWires[133]),
    .Test_en_W_in(Test_enWires[132]),
    .chany_bottom_in(sb_1__1__113_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__114_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_124_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__124_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__124_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__124_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__124_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__124_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__124_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__124_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__124_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__124_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__124_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__124_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__124_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__124_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__124_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__124_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__124_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__124_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__124_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__124_ccff_tail[0])
  );


  cby_1__1_
  cby_11__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[422]),
    .prog_clk_0_W_in(prog_clk_0_wires[421]),
    .Test_en_E_out(Test_enWires[155]),
    .Test_en_W_in(Test_enWires[154]),
    .chany_bottom_in(sb_1__1__114_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__115_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_125_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__125_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__125_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__125_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__125_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__125_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__125_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__125_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__125_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__125_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__125_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__125_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__125_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__125_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__125_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__125_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__125_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__125_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__125_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__125_ccff_tail[0])
  );


  cby_1__1_
  cby_11__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[425]),
    .prog_clk_0_W_in(prog_clk_0_wires[424]),
    .Test_en_E_out(Test_enWires[177]),
    .Test_en_W_in(Test_enWires[176]),
    .chany_bottom_in(sb_1__1__115_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__116_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_126_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__126_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__126_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__126_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__126_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__126_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__126_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__126_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__126_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__126_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__126_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__126_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__126_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__126_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__126_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__126_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__126_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__126_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__126_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__126_ccff_tail[0])
  );


  cby_1__1_
  cby_11__8_
  (
    .clk_2_S_out(clk_2_wires[130]),
    .clk_2_N_in(clk_2_wires[129]),
    .prog_clk_2_S_out(prog_clk_2_wires[130]),
    .prog_clk_2_N_in(prog_clk_2_wires[129]),
    .prog_clk_0_S_out(prog_clk_0_wires[428]),
    .prog_clk_0_W_in(prog_clk_0_wires[427]),
    .Test_en_E_out(Test_enWires[199]),
    .Test_en_W_in(Test_enWires[198]),
    .chany_bottom_in(sb_1__1__116_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__117_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_127_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__127_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__127_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__127_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__127_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__127_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__127_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__127_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__127_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__127_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__127_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__127_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__127_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__127_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__127_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__127_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__127_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__127_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__127_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__127_ccff_tail[0])
  );


  cby_1__1_
  cby_11__9_
  (
    .clk_2_N_out(clk_2_wires[128]),
    .clk_2_S_in(clk_2_wires[127]),
    .prog_clk_2_N_out(prog_clk_2_wires[128]),
    .prog_clk_2_S_in(prog_clk_2_wires[127]),
    .prog_clk_0_S_out(prog_clk_0_wires[431]),
    .prog_clk_0_W_in(prog_clk_0_wires[430]),
    .Test_en_E_out(Test_enWires[221]),
    .Test_en_W_in(Test_enWires[220]),
    .chany_bottom_in(sb_1__1__117_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__118_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_128_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__128_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__128_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__128_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__128_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__128_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__128_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__128_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__128_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__128_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__128_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__128_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__128_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__128_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__128_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__128_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__128_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__128_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__128_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__128_ccff_tail[0])
  );


  cby_1__1_
  cby_11__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[434]),
    .prog_clk_0_W_in(prog_clk_0_wires[433]),
    .Test_en_E_out(Test_enWires[243]),
    .Test_en_W_in(Test_enWires[242]),
    .chany_bottom_in(sb_1__1__118_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__119_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_129_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__129_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__129_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__129_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__129_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__129_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__129_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__129_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__129_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__129_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__129_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__129_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__129_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__129_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__129_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__129_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__129_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__129_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__129_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__129_ccff_tail[0])
  );


  cby_1__1_
  cby_11__11_
  (
    .clk_2_N_out(clk_2_wires[135]),
    .clk_2_S_in(clk_2_wires[134]),
    .prog_clk_2_N_out(prog_clk_2_wires[135]),
    .prog_clk_2_S_in(prog_clk_2_wires[134]),
    .prog_clk_0_S_out(prog_clk_0_wires[437]),
    .prog_clk_0_W_in(prog_clk_0_wires[436]),
    .Test_en_E_out(Test_enWires[265]),
    .Test_en_W_in(Test_enWires[264]),
    .chany_bottom_in(sb_1__1__119_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__120_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_130_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__130_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__130_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__130_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__130_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__130_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__130_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__130_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__130_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__130_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__130_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__130_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__130_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__130_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__130_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__130_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__130_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__130_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__130_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__130_ccff_tail[0])
  );


  cby_1__1_
  cby_11__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[442]),
    .prog_clk_0_S_out(prog_clk_0_wires[440]),
    .prog_clk_0_W_in(prog_clk_0_wires[439]),
    .Test_en_E_out(Test_enWires[287]),
    .Test_en_W_in(Test_enWires[286]),
    .chany_bottom_in(sb_1__1__120_chany_top_out[0:19]),
    .chany_top_in(sb_1__12__10_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_131_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__131_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__131_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__131_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__131_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__131_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__131_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__131_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__131_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__131_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__131_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__131_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__131_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__131_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__131_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__131_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__131_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__131_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__131_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__131_ccff_tail[0])
  );


  cby_2__1_
  cby_12__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[445]),
    .prog_clk_0_W_in(prog_clk_0_wires[444]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_11_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_11_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__0_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__0__0_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_132_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__0_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_12__1__0_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__0_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__0_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__0_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__0_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__0_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__0_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__0_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__0_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__0_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__0_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__0_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__0_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__0_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__0_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__0_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__0_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_11_ccff_tail[0])
  );


  cby_2__1_
  cby_12__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[448]),
    .prog_clk_0_W_in(prog_clk_0_wires[447]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_10_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_10_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__1_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__0_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_133_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__1_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_12__1__1_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__1_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__1_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__1_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__1_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__1_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__1_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__1_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__1_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__1_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__1_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__1_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__1_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__1_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__1_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__1_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__1_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_10_ccff_tail[0])
  );


  cby_2__1_
  cby_12__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[451]),
    .prog_clk_0_W_in(prog_clk_0_wires[450]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_9_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_9_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__2_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__1_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_134_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__2_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_12__1__2_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__2_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__2_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__2_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__2_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__2_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__2_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__2_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__2_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__2_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__2_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__2_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__2_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__2_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__2_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__2_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__2_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_9_ccff_tail[0])
  );


  cby_2__1_
  cby_12__4_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[454]),
    .prog_clk_0_W_in(prog_clk_0_wires[453]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_8_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_8_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__3_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__2_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_135_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__3_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_12__1__3_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__3_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__3_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__3_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__3_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__3_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__3_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__3_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__3_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__3_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__3_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__3_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__3_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__3_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__3_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__3_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__3_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_8_ccff_tail[0])
  );


  cby_2__1_
  cby_12__5_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[457]),
    .prog_clk_0_W_in(prog_clk_0_wires[456]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_7_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_7_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__4_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__3_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_136_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__4_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_12__1__4_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__4_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__4_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__4_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__4_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__4_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__4_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__4_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__4_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__4_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__4_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__4_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__4_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__4_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__4_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__4_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__4_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_7_ccff_tail[0])
  );


  cby_2__1_
  cby_12__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[460]),
    .prog_clk_0_W_in(prog_clk_0_wires[459]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_6_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_6_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__5_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__4_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_137_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__5_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_12__1__5_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__5_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__5_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__5_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__5_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__5_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__5_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__5_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__5_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__5_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__5_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__5_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__5_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__5_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__5_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__5_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__5_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_6_ccff_tail[0])
  );


  cby_2__1_
  cby_12__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[463]),
    .prog_clk_0_W_in(prog_clk_0_wires[462]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_5_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_5_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__6_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__5_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_138_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__6_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_12__1__6_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__6_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__6_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__6_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__6_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__6_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__6_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__6_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__6_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__6_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__6_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__6_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__6_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__6_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__6_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__6_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__6_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_5_ccff_tail[0])
  );


  cby_2__1_
  cby_12__8_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[466]),
    .prog_clk_0_W_in(prog_clk_0_wires[465]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_4_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_4_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__7_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__6_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__7_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_139_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__7_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_12__1__7_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__7_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__7_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__7_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__7_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__7_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__7_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__7_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__7_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__7_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__7_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__7_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__7_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__7_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__7_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__7_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__7_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_4_ccff_tail[0])
  );


  cby_2__1_
  cby_12__9_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[469]),
    .prog_clk_0_W_in(prog_clk_0_wires[468]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_3_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_3_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__8_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__7_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__8_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_140_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__8_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__8_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_12__1__8_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__8_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__8_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__8_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__8_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__8_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__8_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__8_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__8_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__8_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__8_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__8_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__8_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__8_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__8_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__8_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__8_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_3_ccff_tail[0])
  );


  cby_2__1_
  cby_12__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[472]),
    .prog_clk_0_W_in(prog_clk_0_wires[471]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_2_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_2_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__9_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__8_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__9_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_141_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__9_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__9_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_12__1__9_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__9_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__9_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__9_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__9_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__9_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__9_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__9_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__9_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__9_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__9_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__9_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__9_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__9_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__9_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__9_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__9_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_2_ccff_tail[0])
  );


  cby_2__1_
  cby_12__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[475]),
    .prog_clk_0_W_in(prog_clk_0_wires[474]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_1_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_1_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__10_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__9_chany_top_out[0:19]),
    .chany_top_in(sb_12__1__10_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_142_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__10_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__10_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_12__1__10_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__10_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__10_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__10_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__10_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__10_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__10_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__10_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__10_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__10_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__10_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__10_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__10_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__10_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__10_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__10_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__10_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_1_ccff_tail[0])
  );


  cby_2__1_
  cby_12__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[480]),
    .prog_clk_0_S_out(prog_clk_0_wires[478]),
    .prog_clk_0_W_in(prog_clk_0_wires[477]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_0_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_0_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__11_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__10_chany_top_out[0:19]),
    .chany_top_in(sb_12__12__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_143_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__11_chany_bottom_out[0:19]),
    .chany_top_out(cby_12__1__11_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_12__1__11_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__11_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__11_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__11_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__11_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__11_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__11_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__11_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__11_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__11_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__11_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__11_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__11_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__11_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__11_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__11_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__11_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_0_ccff_tail[0])
  );


  direct_interc
  direct_interc_0_
  (
    .in(grid_clb_1_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_0_out[0])
  );


  direct_interc
  direct_interc_1_
  (
    .in(grid_clb_2_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_1_out[0])
  );


  direct_interc
  direct_interc_2_
  (
    .in(grid_clb_3_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_2_out[0])
  );


  direct_interc
  direct_interc_3_
  (
    .in(grid_clb_4_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_3_out[0])
  );


  direct_interc
  direct_interc_4_
  (
    .in(grid_clb_5_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_4_out[0])
  );


  direct_interc
  direct_interc_5_
  (
    .in(grid_clb_6_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_5_out[0])
  );


  direct_interc
  direct_interc_6_
  (
    .in(grid_clb_7_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_6_out[0])
  );


  direct_interc
  direct_interc_7_
  (
    .in(grid_clb_8_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_7_out[0])
  );


  direct_interc
  direct_interc_8_
  (
    .in(grid_clb_9_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_8_out[0])
  );


  direct_interc
  direct_interc_9_
  (
    .in(grid_clb_10_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_9_out[0])
  );


  direct_interc
  direct_interc_10_
  (
    .in(grid_clb_11_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_10_out[0])
  );


  direct_interc
  direct_interc_11_
  (
    .in(grid_clb_13_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_11_out[0])
  );


  direct_interc
  direct_interc_12_
  (
    .in(grid_clb_14_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_12_out[0])
  );


  direct_interc
  direct_interc_13_
  (
    .in(grid_clb_15_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_13_out[0])
  );


  direct_interc
  direct_interc_14_
  (
    .in(grid_clb_16_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_14_out[0])
  );


  direct_interc
  direct_interc_15_
  (
    .in(grid_clb_17_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_15_out[0])
  );


  direct_interc
  direct_interc_16_
  (
    .in(grid_clb_18_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_16_out[0])
  );


  direct_interc
  direct_interc_17_
  (
    .in(grid_clb_19_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_17_out[0])
  );


  direct_interc
  direct_interc_18_
  (
    .in(grid_clb_20_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_18_out[0])
  );


  direct_interc
  direct_interc_19_
  (
    .in(grid_clb_21_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_19_out[0])
  );


  direct_interc
  direct_interc_20_
  (
    .in(grid_clb_22_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_20_out[0])
  );


  direct_interc
  direct_interc_21_
  (
    .in(grid_clb_23_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_21_out[0])
  );


  direct_interc
  direct_interc_22_
  (
    .in(grid_clb_25_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_22_out[0])
  );


  direct_interc
  direct_interc_23_
  (
    .in(grid_clb_26_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_23_out[0])
  );


  direct_interc
  direct_interc_24_
  (
    .in(grid_clb_27_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_24_out[0])
  );


  direct_interc
  direct_interc_25_
  (
    .in(grid_clb_28_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_25_out[0])
  );


  direct_interc
  direct_interc_26_
  (
    .in(grid_clb_29_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_26_out[0])
  );


  direct_interc
  direct_interc_27_
  (
    .in(grid_clb_30_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_27_out[0])
  );


  direct_interc
  direct_interc_28_
  (
    .in(grid_clb_31_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_28_out[0])
  );


  direct_interc
  direct_interc_29_
  (
    .in(grid_clb_32_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_29_out[0])
  );


  direct_interc
  direct_interc_30_
  (
    .in(grid_clb_33_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_30_out[0])
  );


  direct_interc
  direct_interc_31_
  (
    .in(grid_clb_34_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_31_out[0])
  );


  direct_interc
  direct_interc_32_
  (
    .in(grid_clb_35_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_32_out[0])
  );


  direct_interc
  direct_interc_33_
  (
    .in(grid_clb_37_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_33_out[0])
  );


  direct_interc
  direct_interc_34_
  (
    .in(grid_clb_38_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_34_out[0])
  );


  direct_interc
  direct_interc_35_
  (
    .in(grid_clb_39_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_35_out[0])
  );


  direct_interc
  direct_interc_36_
  (
    .in(grid_clb_40_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_36_out[0])
  );


  direct_interc
  direct_interc_37_
  (
    .in(grid_clb_41_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_37_out[0])
  );


  direct_interc
  direct_interc_38_
  (
    .in(grid_clb_42_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_38_out[0])
  );


  direct_interc
  direct_interc_39_
  (
    .in(grid_clb_43_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_39_out[0])
  );


  direct_interc
  direct_interc_40_
  (
    .in(grid_clb_44_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_40_out[0])
  );


  direct_interc
  direct_interc_41_
  (
    .in(grid_clb_45_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_41_out[0])
  );


  direct_interc
  direct_interc_42_
  (
    .in(grid_clb_46_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_42_out[0])
  );


  direct_interc
  direct_interc_43_
  (
    .in(grid_clb_47_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_43_out[0])
  );


  direct_interc
  direct_interc_44_
  (
    .in(grid_clb_49_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_44_out[0])
  );


  direct_interc
  direct_interc_45_
  (
    .in(grid_clb_50_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_45_out[0])
  );


  direct_interc
  direct_interc_46_
  (
    .in(grid_clb_51_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_46_out[0])
  );


  direct_interc
  direct_interc_47_
  (
    .in(grid_clb_52_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_47_out[0])
  );


  direct_interc
  direct_interc_48_
  (
    .in(grid_clb_53_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_48_out[0])
  );


  direct_interc
  direct_interc_49_
  (
    .in(grid_clb_54_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_49_out[0])
  );


  direct_interc
  direct_interc_50_
  (
    .in(grid_clb_55_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_50_out[0])
  );


  direct_interc
  direct_interc_51_
  (
    .in(grid_clb_56_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_51_out[0])
  );


  direct_interc
  direct_interc_52_
  (
    .in(grid_clb_57_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_52_out[0])
  );


  direct_interc
  direct_interc_53_
  (
    .in(grid_clb_58_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_53_out[0])
  );


  direct_interc
  direct_interc_54_
  (
    .in(grid_clb_59_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_54_out[0])
  );


  direct_interc
  direct_interc_55_
  (
    .in(grid_clb_61_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_55_out[0])
  );


  direct_interc
  direct_interc_56_
  (
    .in(grid_clb_62_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_56_out[0])
  );


  direct_interc
  direct_interc_57_
  (
    .in(grid_clb_63_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_57_out[0])
  );


  direct_interc
  direct_interc_58_
  (
    .in(grid_clb_64_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_58_out[0])
  );


  direct_interc
  direct_interc_59_
  (
    .in(grid_clb_65_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_59_out[0])
  );


  direct_interc
  direct_interc_60_
  (
    .in(grid_clb_66_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_60_out[0])
  );


  direct_interc
  direct_interc_61_
  (
    .in(grid_clb_67_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_61_out[0])
  );


  direct_interc
  direct_interc_62_
  (
    .in(grid_clb_68_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_62_out[0])
  );


  direct_interc
  direct_interc_63_
  (
    .in(grid_clb_69_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_63_out[0])
  );


  direct_interc
  direct_interc_64_
  (
    .in(grid_clb_70_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_64_out[0])
  );


  direct_interc
  direct_interc_65_
  (
    .in(grid_clb_71_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_65_out[0])
  );


  direct_interc
  direct_interc_66_
  (
    .in(grid_clb_73_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_66_out[0])
  );


  direct_interc
  direct_interc_67_
  (
    .in(grid_clb_74_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_67_out[0])
  );


  direct_interc
  direct_interc_68_
  (
    .in(grid_clb_75_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_68_out[0])
  );


  direct_interc
  direct_interc_69_
  (
    .in(grid_clb_76_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_69_out[0])
  );


  direct_interc
  direct_interc_70_
  (
    .in(grid_clb_77_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_70_out[0])
  );


  direct_interc
  direct_interc_71_
  (
    .in(grid_clb_78_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_71_out[0])
  );


  direct_interc
  direct_interc_72_
  (
    .in(grid_clb_79_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_72_out[0])
  );


  direct_interc
  direct_interc_73_
  (
    .in(grid_clb_80_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_73_out[0])
  );


  direct_interc
  direct_interc_74_
  (
    .in(grid_clb_81_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_74_out[0])
  );


  direct_interc
  direct_interc_75_
  (
    .in(grid_clb_82_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_75_out[0])
  );


  direct_interc
  direct_interc_76_
  (
    .in(grid_clb_83_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_76_out[0])
  );


  direct_interc
  direct_interc_77_
  (
    .in(grid_clb_85_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_77_out[0])
  );


  direct_interc
  direct_interc_78_
  (
    .in(grid_clb_86_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_78_out[0])
  );


  direct_interc
  direct_interc_79_
  (
    .in(grid_clb_87_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_79_out[0])
  );


  direct_interc
  direct_interc_80_
  (
    .in(grid_clb_88_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_80_out[0])
  );


  direct_interc
  direct_interc_81_
  (
    .in(grid_clb_89_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_81_out[0])
  );


  direct_interc
  direct_interc_82_
  (
    .in(grid_clb_90_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_82_out[0])
  );


  direct_interc
  direct_interc_83_
  (
    .in(grid_clb_91_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_83_out[0])
  );


  direct_interc
  direct_interc_84_
  (
    .in(grid_clb_92_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_84_out[0])
  );


  direct_interc
  direct_interc_85_
  (
    .in(grid_clb_93_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_85_out[0])
  );


  direct_interc
  direct_interc_86_
  (
    .in(grid_clb_94_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_86_out[0])
  );


  direct_interc
  direct_interc_87_
  (
    .in(grid_clb_95_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_87_out[0])
  );


  direct_interc
  direct_interc_88_
  (
    .in(grid_clb_97_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_88_out[0])
  );


  direct_interc
  direct_interc_89_
  (
    .in(grid_clb_98_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_89_out[0])
  );


  direct_interc
  direct_interc_90_
  (
    .in(grid_clb_99_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_90_out[0])
  );


  direct_interc
  direct_interc_91_
  (
    .in(grid_clb_100_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_91_out[0])
  );


  direct_interc
  direct_interc_92_
  (
    .in(grid_clb_101_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_92_out[0])
  );


  direct_interc
  direct_interc_93_
  (
    .in(grid_clb_102_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_93_out[0])
  );


  direct_interc
  direct_interc_94_
  (
    .in(grid_clb_103_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_94_out[0])
  );


  direct_interc
  direct_interc_95_
  (
    .in(grid_clb_104_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_95_out[0])
  );


  direct_interc
  direct_interc_96_
  (
    .in(grid_clb_105_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_96_out[0])
  );


  direct_interc
  direct_interc_97_
  (
    .in(grid_clb_106_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_97_out[0])
  );


  direct_interc
  direct_interc_98_
  (
    .in(grid_clb_107_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_98_out[0])
  );


  direct_interc
  direct_interc_99_
  (
    .in(grid_clb_109_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_99_out[0])
  );


  direct_interc
  direct_interc_100_
  (
    .in(grid_clb_110_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_100_out[0])
  );


  direct_interc
  direct_interc_101_
  (
    .in(grid_clb_111_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_101_out[0])
  );


  direct_interc
  direct_interc_102_
  (
    .in(grid_clb_112_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_102_out[0])
  );


  direct_interc
  direct_interc_103_
  (
    .in(grid_clb_113_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_103_out[0])
  );


  direct_interc
  direct_interc_104_
  (
    .in(grid_clb_114_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_104_out[0])
  );


  direct_interc
  direct_interc_105_
  (
    .in(grid_clb_115_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_105_out[0])
  );


  direct_interc
  direct_interc_106_
  (
    .in(grid_clb_116_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_106_out[0])
  );


  direct_interc
  direct_interc_107_
  (
    .in(grid_clb_117_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_107_out[0])
  );


  direct_interc
  direct_interc_108_
  (
    .in(grid_clb_118_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_108_out[0])
  );


  direct_interc
  direct_interc_109_
  (
    .in(grid_clb_119_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_109_out[0])
  );


  direct_interc
  direct_interc_110_
  (
    .in(grid_clb_121_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_110_out[0])
  );


  direct_interc
  direct_interc_111_
  (
    .in(grid_clb_122_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_111_out[0])
  );


  direct_interc
  direct_interc_112_
  (
    .in(grid_clb_123_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_112_out[0])
  );


  direct_interc
  direct_interc_113_
  (
    .in(grid_clb_124_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_113_out[0])
  );


  direct_interc
  direct_interc_114_
  (
    .in(grid_clb_125_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_114_out[0])
  );


  direct_interc
  direct_interc_115_
  (
    .in(grid_clb_126_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_115_out[0])
  );


  direct_interc
  direct_interc_116_
  (
    .in(grid_clb_127_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_116_out[0])
  );


  direct_interc
  direct_interc_117_
  (
    .in(grid_clb_128_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_117_out[0])
  );


  direct_interc
  direct_interc_118_
  (
    .in(grid_clb_129_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_118_out[0])
  );


  direct_interc
  direct_interc_119_
  (
    .in(grid_clb_130_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_119_out[0])
  );


  direct_interc
  direct_interc_120_
  (
    .in(grid_clb_131_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_120_out[0])
  );


  direct_interc
  direct_interc_121_
  (
    .in(grid_clb_133_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_121_out[0])
  );


  direct_interc
  direct_interc_122_
  (
    .in(grid_clb_134_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_122_out[0])
  );


  direct_interc
  direct_interc_123_
  (
    .in(grid_clb_135_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_123_out[0])
  );


  direct_interc
  direct_interc_124_
  (
    .in(grid_clb_136_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_124_out[0])
  );


  direct_interc
  direct_interc_125_
  (
    .in(grid_clb_137_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_125_out[0])
  );


  direct_interc
  direct_interc_126_
  (
    .in(grid_clb_138_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_126_out[0])
  );


  direct_interc
  direct_interc_127_
  (
    .in(grid_clb_139_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_127_out[0])
  );


  direct_interc
  direct_interc_128_
  (
    .in(grid_clb_140_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_128_out[0])
  );


  direct_interc
  direct_interc_129_
  (
    .in(grid_clb_141_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_129_out[0])
  );


  direct_interc
  direct_interc_130_
  (
    .in(grid_clb_142_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_130_out[0])
  );


  direct_interc
  direct_interc_131_
  (
    .in(grid_clb_143_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_131_out[0])
  );


  direct_interc
  direct_interc_132_
  (
    .in(grid_clb_1_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_132_out[0])
  );


  direct_interc
  direct_interc_133_
  (
    .in(grid_clb_2_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_133_out[0])
  );


  direct_interc
  direct_interc_134_
  (
    .in(grid_clb_3_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_134_out[0])
  );


  direct_interc
  direct_interc_135_
  (
    .in(grid_clb_4_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_135_out[0])
  );


  direct_interc
  direct_interc_136_
  (
    .in(grid_clb_5_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_136_out[0])
  );


  direct_interc
  direct_interc_137_
  (
    .in(grid_clb_6_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_137_out[0])
  );


  direct_interc
  direct_interc_138_
  (
    .in(grid_clb_7_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_138_out[0])
  );


  direct_interc
  direct_interc_139_
  (
    .in(grid_clb_8_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_139_out[0])
  );


  direct_interc
  direct_interc_140_
  (
    .in(grid_clb_9_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_140_out[0])
  );


  direct_interc
  direct_interc_141_
  (
    .in(grid_clb_10_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_141_out[0])
  );


  direct_interc
  direct_interc_142_
  (
    .in(grid_clb_11_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_142_out[0])
  );


  direct_interc
  direct_interc_143_
  (
    .in(grid_clb_13_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_143_out[0])
  );


  direct_interc
  direct_interc_144_
  (
    .in(grid_clb_14_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_144_out[0])
  );


  direct_interc
  direct_interc_145_
  (
    .in(grid_clb_15_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_145_out[0])
  );


  direct_interc
  direct_interc_146_
  (
    .in(grid_clb_16_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_146_out[0])
  );


  direct_interc
  direct_interc_147_
  (
    .in(grid_clb_17_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_147_out[0])
  );


  direct_interc
  direct_interc_148_
  (
    .in(grid_clb_18_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_148_out[0])
  );


  direct_interc
  direct_interc_149_
  (
    .in(grid_clb_19_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_149_out[0])
  );


  direct_interc
  direct_interc_150_
  (
    .in(grid_clb_20_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_150_out[0])
  );


  direct_interc
  direct_interc_151_
  (
    .in(grid_clb_21_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_151_out[0])
  );


  direct_interc
  direct_interc_152_
  (
    .in(grid_clb_22_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_152_out[0])
  );


  direct_interc
  direct_interc_153_
  (
    .in(grid_clb_23_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_153_out[0])
  );


  direct_interc
  direct_interc_154_
  (
    .in(grid_clb_25_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_154_out[0])
  );


  direct_interc
  direct_interc_155_
  (
    .in(grid_clb_26_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_155_out[0])
  );


  direct_interc
  direct_interc_156_
  (
    .in(grid_clb_27_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_156_out[0])
  );


  direct_interc
  direct_interc_157_
  (
    .in(grid_clb_28_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_157_out[0])
  );


  direct_interc
  direct_interc_158_
  (
    .in(grid_clb_29_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_158_out[0])
  );


  direct_interc
  direct_interc_159_
  (
    .in(grid_clb_30_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_159_out[0])
  );


  direct_interc
  direct_interc_160_
  (
    .in(grid_clb_31_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_160_out[0])
  );


  direct_interc
  direct_interc_161_
  (
    .in(grid_clb_32_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_161_out[0])
  );


  direct_interc
  direct_interc_162_
  (
    .in(grid_clb_33_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_162_out[0])
  );


  direct_interc
  direct_interc_163_
  (
    .in(grid_clb_34_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_163_out[0])
  );


  direct_interc
  direct_interc_164_
  (
    .in(grid_clb_35_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_164_out[0])
  );


  direct_interc
  direct_interc_165_
  (
    .in(grid_clb_37_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_165_out[0])
  );


  direct_interc
  direct_interc_166_
  (
    .in(grid_clb_38_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_166_out[0])
  );


  direct_interc
  direct_interc_167_
  (
    .in(grid_clb_39_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_167_out[0])
  );


  direct_interc
  direct_interc_168_
  (
    .in(grid_clb_40_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_168_out[0])
  );


  direct_interc
  direct_interc_169_
  (
    .in(grid_clb_41_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_169_out[0])
  );


  direct_interc
  direct_interc_170_
  (
    .in(grid_clb_42_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_170_out[0])
  );


  direct_interc
  direct_interc_171_
  (
    .in(grid_clb_43_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_171_out[0])
  );


  direct_interc
  direct_interc_172_
  (
    .in(grid_clb_44_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_172_out[0])
  );


  direct_interc
  direct_interc_173_
  (
    .in(grid_clb_45_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_173_out[0])
  );


  direct_interc
  direct_interc_174_
  (
    .in(grid_clb_46_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_174_out[0])
  );


  direct_interc
  direct_interc_175_
  (
    .in(grid_clb_47_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_175_out[0])
  );


  direct_interc
  direct_interc_176_
  (
    .in(grid_clb_49_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_176_out[0])
  );


  direct_interc
  direct_interc_177_
  (
    .in(grid_clb_50_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_177_out[0])
  );


  direct_interc
  direct_interc_178_
  (
    .in(grid_clb_51_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_178_out[0])
  );


  direct_interc
  direct_interc_179_
  (
    .in(grid_clb_52_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_179_out[0])
  );


  direct_interc
  direct_interc_180_
  (
    .in(grid_clb_53_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_180_out[0])
  );


  direct_interc
  direct_interc_181_
  (
    .in(grid_clb_54_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_181_out[0])
  );


  direct_interc
  direct_interc_182_
  (
    .in(grid_clb_55_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_182_out[0])
  );


  direct_interc
  direct_interc_183_
  (
    .in(grid_clb_56_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_183_out[0])
  );


  direct_interc
  direct_interc_184_
  (
    .in(grid_clb_57_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_184_out[0])
  );


  direct_interc
  direct_interc_185_
  (
    .in(grid_clb_58_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_185_out[0])
  );


  direct_interc
  direct_interc_186_
  (
    .in(grid_clb_59_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_186_out[0])
  );


  direct_interc
  direct_interc_187_
  (
    .in(grid_clb_61_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_187_out[0])
  );


  direct_interc
  direct_interc_188_
  (
    .in(grid_clb_62_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_188_out[0])
  );


  direct_interc
  direct_interc_189_
  (
    .in(grid_clb_63_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_189_out[0])
  );


  direct_interc
  direct_interc_190_
  (
    .in(grid_clb_64_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_190_out[0])
  );


  direct_interc
  direct_interc_191_
  (
    .in(grid_clb_65_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_191_out[0])
  );


  direct_interc
  direct_interc_192_
  (
    .in(grid_clb_66_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_192_out[0])
  );


  direct_interc
  direct_interc_193_
  (
    .in(grid_clb_67_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_193_out[0])
  );


  direct_interc
  direct_interc_194_
  (
    .in(grid_clb_68_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_194_out[0])
  );


  direct_interc
  direct_interc_195_
  (
    .in(grid_clb_69_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_195_out[0])
  );


  direct_interc
  direct_interc_196_
  (
    .in(grid_clb_70_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_196_out[0])
  );


  direct_interc
  direct_interc_197_
  (
    .in(grid_clb_71_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_197_out[0])
  );


  direct_interc
  direct_interc_198_
  (
    .in(grid_clb_73_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_198_out[0])
  );


  direct_interc
  direct_interc_199_
  (
    .in(grid_clb_74_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_199_out[0])
  );


  direct_interc
  direct_interc_200_
  (
    .in(grid_clb_75_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_200_out[0])
  );


  direct_interc
  direct_interc_201_
  (
    .in(grid_clb_76_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_201_out[0])
  );


  direct_interc
  direct_interc_202_
  (
    .in(grid_clb_77_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_202_out[0])
  );


  direct_interc
  direct_interc_203_
  (
    .in(grid_clb_78_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_203_out[0])
  );


  direct_interc
  direct_interc_204_
  (
    .in(grid_clb_79_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_204_out[0])
  );


  direct_interc
  direct_interc_205_
  (
    .in(grid_clb_80_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_205_out[0])
  );


  direct_interc
  direct_interc_206_
  (
    .in(grid_clb_81_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_206_out[0])
  );


  direct_interc
  direct_interc_207_
  (
    .in(grid_clb_82_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_207_out[0])
  );


  direct_interc
  direct_interc_208_
  (
    .in(grid_clb_83_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_208_out[0])
  );


  direct_interc
  direct_interc_209_
  (
    .in(grid_clb_85_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_209_out[0])
  );


  direct_interc
  direct_interc_210_
  (
    .in(grid_clb_86_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_210_out[0])
  );


  direct_interc
  direct_interc_211_
  (
    .in(grid_clb_87_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_211_out[0])
  );


  direct_interc
  direct_interc_212_
  (
    .in(grid_clb_88_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_212_out[0])
  );


  direct_interc
  direct_interc_213_
  (
    .in(grid_clb_89_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_213_out[0])
  );


  direct_interc
  direct_interc_214_
  (
    .in(grid_clb_90_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_214_out[0])
  );


  direct_interc
  direct_interc_215_
  (
    .in(grid_clb_91_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_215_out[0])
  );


  direct_interc
  direct_interc_216_
  (
    .in(grid_clb_92_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_216_out[0])
  );


  direct_interc
  direct_interc_217_
  (
    .in(grid_clb_93_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_217_out[0])
  );


  direct_interc
  direct_interc_218_
  (
    .in(grid_clb_94_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_218_out[0])
  );


  direct_interc
  direct_interc_219_
  (
    .in(grid_clb_95_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_219_out[0])
  );


  direct_interc
  direct_interc_220_
  (
    .in(grid_clb_97_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_220_out[0])
  );


  direct_interc
  direct_interc_221_
  (
    .in(grid_clb_98_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_221_out[0])
  );


  direct_interc
  direct_interc_222_
  (
    .in(grid_clb_99_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_222_out[0])
  );


  direct_interc
  direct_interc_223_
  (
    .in(grid_clb_100_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_223_out[0])
  );


  direct_interc
  direct_interc_224_
  (
    .in(grid_clb_101_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_224_out[0])
  );


  direct_interc
  direct_interc_225_
  (
    .in(grid_clb_102_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_225_out[0])
  );


  direct_interc
  direct_interc_226_
  (
    .in(grid_clb_103_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_226_out[0])
  );


  direct_interc
  direct_interc_227_
  (
    .in(grid_clb_104_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_227_out[0])
  );


  direct_interc
  direct_interc_228_
  (
    .in(grid_clb_105_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_228_out[0])
  );


  direct_interc
  direct_interc_229_
  (
    .in(grid_clb_106_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_229_out[0])
  );


  direct_interc
  direct_interc_230_
  (
    .in(grid_clb_107_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_230_out[0])
  );


  direct_interc
  direct_interc_231_
  (
    .in(grid_clb_109_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_231_out[0])
  );


  direct_interc
  direct_interc_232_
  (
    .in(grid_clb_110_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_232_out[0])
  );


  direct_interc
  direct_interc_233_
  (
    .in(grid_clb_111_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_233_out[0])
  );


  direct_interc
  direct_interc_234_
  (
    .in(grid_clb_112_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_234_out[0])
  );


  direct_interc
  direct_interc_235_
  (
    .in(grid_clb_113_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_235_out[0])
  );


  direct_interc
  direct_interc_236_
  (
    .in(grid_clb_114_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_236_out[0])
  );


  direct_interc
  direct_interc_237_
  (
    .in(grid_clb_115_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_237_out[0])
  );


  direct_interc
  direct_interc_238_
  (
    .in(grid_clb_116_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_238_out[0])
  );


  direct_interc
  direct_interc_239_
  (
    .in(grid_clb_117_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_239_out[0])
  );


  direct_interc
  direct_interc_240_
  (
    .in(grid_clb_118_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_240_out[0])
  );


  direct_interc
  direct_interc_241_
  (
    .in(grid_clb_119_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_241_out[0])
  );


  direct_interc
  direct_interc_242_
  (
    .in(grid_clb_121_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_242_out[0])
  );


  direct_interc
  direct_interc_243_
  (
    .in(grid_clb_122_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_243_out[0])
  );


  direct_interc
  direct_interc_244_
  (
    .in(grid_clb_123_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_244_out[0])
  );


  direct_interc
  direct_interc_245_
  (
    .in(grid_clb_124_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_245_out[0])
  );


  direct_interc
  direct_interc_246_
  (
    .in(grid_clb_125_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_246_out[0])
  );


  direct_interc
  direct_interc_247_
  (
    .in(grid_clb_126_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_247_out[0])
  );


  direct_interc
  direct_interc_248_
  (
    .in(grid_clb_127_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_248_out[0])
  );


  direct_interc
  direct_interc_249_
  (
    .in(grid_clb_128_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_249_out[0])
  );


  direct_interc
  direct_interc_250_
  (
    .in(grid_clb_129_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_250_out[0])
  );


  direct_interc
  direct_interc_251_
  (
    .in(grid_clb_130_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_251_out[0])
  );


  direct_interc
  direct_interc_252_
  (
    .in(grid_clb_131_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_252_out[0])
  );


  direct_interc
  direct_interc_253_
  (
    .in(grid_clb_133_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_253_out[0])
  );


  direct_interc
  direct_interc_254_
  (
    .in(grid_clb_134_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_254_out[0])
  );


  direct_interc
  direct_interc_255_
  (
    .in(grid_clb_135_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_255_out[0])
  );


  direct_interc
  direct_interc_256_
  (
    .in(grid_clb_136_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_256_out[0])
  );


  direct_interc
  direct_interc_257_
  (
    .in(grid_clb_137_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_257_out[0])
  );


  direct_interc
  direct_interc_258_
  (
    .in(grid_clb_138_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_258_out[0])
  );


  direct_interc
  direct_interc_259_
  (
    .in(grid_clb_139_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_259_out[0])
  );


  direct_interc
  direct_interc_260_
  (
    .in(grid_clb_140_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_260_out[0])
  );


  direct_interc
  direct_interc_261_
  (
    .in(grid_clb_141_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_261_out[0])
  );


  direct_interc
  direct_interc_262_
  (
    .in(grid_clb_142_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_262_out[0])
  );


  direct_interc
  direct_interc_263_
  (
    .in(grid_clb_143_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_263_out[0])
  );


  direct_interc
  direct_interc_264_
  (
    .in(grid_clb_0_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_264_out[0])
  );


  direct_interc
  direct_interc_265_
  (
    .in(grid_clb_12_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_265_out[0])
  );


  direct_interc
  direct_interc_266_
  (
    .in(grid_clb_24_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_266_out[0])
  );


  direct_interc
  direct_interc_267_
  (
    .in(grid_clb_36_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_267_out[0])
  );


  direct_interc
  direct_interc_268_
  (
    .in(grid_clb_48_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_268_out[0])
  );


  direct_interc
  direct_interc_269_
  (
    .in(grid_clb_60_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_269_out[0])
  );


  direct_interc
  direct_interc_270_
  (
    .in(grid_clb_72_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_270_out[0])
  );


  direct_interc
  direct_interc_271_
  (
    .in(grid_clb_84_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_271_out[0])
  );


  direct_interc
  direct_interc_272_
  (
    .in(grid_clb_96_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_272_out[0])
  );


  direct_interc
  direct_interc_273_
  (
    .in(grid_clb_108_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_273_out[0])
  );


  direct_interc
  direct_interc_274_
  (
    .in(grid_clb_120_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_274_out[0])
  );


endmodule

