

module fpga_core
( pReset, prog_clk, Test_en, IO_ISOL_N, clk, Reset, gfpga_pad_EMBEDDED_IO_HD_SOC_IN, gfpga_pad_EMBEDDED_IO_HD_SOC_OUT, gfpga_pad_EMBEDDED_IO_HD_SOC_DIR, ccff_head, ccff_tail, sc_head, sc_tail ); 
  input [0:0] pReset;
  input [0:0] prog_clk;
  input [0:0] Test_en;
  input [0:0] IO_ISOL_N;
  input [0:0] clk;
  input [0:0] Reset;
  input [0:143] gfpga_pad_EMBEDDED_IO_HD_SOC_IN;
  output [0:143] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT;
  output [0:143] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR;
  input [0:0] ccff_head;
  output [0:0] ccff_tail;
  input sc_head;
  output sc_tail;

  wire [0:0] cbx_1__0__0_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__0_ccff_tail;
  wire [0:29] cbx_1__0__0_chanx_left_out;
  wire [0:29] cbx_1__0__0_chanx_right_out;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__10_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__10_ccff_tail;
  wire [0:29] cbx_1__0__10_chanx_left_out;
  wire [0:29] cbx_1__0__10_chanx_right_out;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__11_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__11_ccff_tail;
  wire [0:29] cbx_1__0__11_chanx_left_out;
  wire [0:29] cbx_1__0__11_chanx_right_out;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__1_ccff_tail;
  wire [0:29] cbx_1__0__1_chanx_left_out;
  wire [0:29] cbx_1__0__1_chanx_right_out;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__2_ccff_tail;
  wire [0:29] cbx_1__0__2_chanx_left_out;
  wire [0:29] cbx_1__0__2_chanx_right_out;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__3_ccff_tail;
  wire [0:29] cbx_1__0__3_chanx_left_out;
  wire [0:29] cbx_1__0__3_chanx_right_out;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__4_ccff_tail;
  wire [0:29] cbx_1__0__4_chanx_left_out;
  wire [0:29] cbx_1__0__4_chanx_right_out;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__5_ccff_tail;
  wire [0:29] cbx_1__0__5_chanx_left_out;
  wire [0:29] cbx_1__0__5_chanx_right_out;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__6_ccff_tail;
  wire [0:29] cbx_1__0__6_chanx_left_out;
  wire [0:29] cbx_1__0__6_chanx_right_out;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__7_ccff_tail;
  wire [0:29] cbx_1__0__7_chanx_left_out;
  wire [0:29] cbx_1__0__7_chanx_right_out;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__8_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__8_ccff_tail;
  wire [0:29] cbx_1__0__8_chanx_left_out;
  wire [0:29] cbx_1__0__8_chanx_right_out;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__9_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__9_ccff_tail;
  wire [0:29] cbx_1__0__9_chanx_left_out;
  wire [0:29] cbx_1__0__9_chanx_right_out;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__0_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__0_ccff_tail;
  wire [0:29] cbx_1__12__0_chanx_left_out;
  wire [0:29] cbx_1__12__0_chanx_right_out;
  wire [0:0] cbx_1__12__0_top_grid_pin_0_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__10_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__10_ccff_tail;
  wire [0:29] cbx_1__12__10_chanx_left_out;
  wire [0:29] cbx_1__12__10_chanx_right_out;
  wire [0:0] cbx_1__12__10_top_grid_pin_0_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__11_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__11_ccff_tail;
  wire [0:29] cbx_1__12__11_chanx_left_out;
  wire [0:29] cbx_1__12__11_chanx_right_out;
  wire [0:0] cbx_1__12__11_top_grid_pin_0_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__1_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__1_ccff_tail;
  wire [0:29] cbx_1__12__1_chanx_left_out;
  wire [0:29] cbx_1__12__1_chanx_right_out;
  wire [0:0] cbx_1__12__1_top_grid_pin_0_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__2_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__2_ccff_tail;
  wire [0:29] cbx_1__12__2_chanx_left_out;
  wire [0:29] cbx_1__12__2_chanx_right_out;
  wire [0:0] cbx_1__12__2_top_grid_pin_0_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__3_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__3_ccff_tail;
  wire [0:29] cbx_1__12__3_chanx_left_out;
  wire [0:29] cbx_1__12__3_chanx_right_out;
  wire [0:0] cbx_1__12__3_top_grid_pin_0_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__4_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__4_ccff_tail;
  wire [0:29] cbx_1__12__4_chanx_left_out;
  wire [0:29] cbx_1__12__4_chanx_right_out;
  wire [0:0] cbx_1__12__4_top_grid_pin_0_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__5_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__5_ccff_tail;
  wire [0:29] cbx_1__12__5_chanx_left_out;
  wire [0:29] cbx_1__12__5_chanx_right_out;
  wire [0:0] cbx_1__12__5_top_grid_pin_0_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__6_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__6_ccff_tail;
  wire [0:29] cbx_1__12__6_chanx_left_out;
  wire [0:29] cbx_1__12__6_chanx_right_out;
  wire [0:0] cbx_1__12__6_top_grid_pin_0_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__7_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__7_ccff_tail;
  wire [0:29] cbx_1__12__7_chanx_left_out;
  wire [0:29] cbx_1__12__7_chanx_right_out;
  wire [0:0] cbx_1__12__7_top_grid_pin_0_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__8_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__8_ccff_tail;
  wire [0:29] cbx_1__12__8_chanx_left_out;
  wire [0:29] cbx_1__12__8_chanx_right_out;
  wire [0:0] cbx_1__12__8_top_grid_pin_0_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_0_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_10_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_11_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_12_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_13_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_14_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_15_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_1_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_2_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_3_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_4_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_5_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_6_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_7_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_8_;
  wire [0:0] cbx_1__12__9_bottom_grid_pin_9_;
  wire [0:0] cbx_1__12__9_ccff_tail;
  wire [0:29] cbx_1__12__9_chanx_left_out;
  wire [0:29] cbx_1__12__9_chanx_right_out;
  wire [0:0] cbx_1__12__9_top_grid_pin_0_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__0_ccff_tail;
  wire [0:29] cbx_1__1__0_chanx_left_out;
  wire [0:29] cbx_1__1__0_chanx_right_out;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__100_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__100_ccff_tail;
  wire [0:29] cbx_1__1__100_chanx_left_out;
  wire [0:29] cbx_1__1__100_chanx_right_out;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__101_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__101_ccff_tail;
  wire [0:29] cbx_1__1__101_chanx_left_out;
  wire [0:29] cbx_1__1__101_chanx_right_out;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__102_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__102_ccff_tail;
  wire [0:29] cbx_1__1__102_chanx_left_out;
  wire [0:29] cbx_1__1__102_chanx_right_out;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__103_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__103_ccff_tail;
  wire [0:29] cbx_1__1__103_chanx_left_out;
  wire [0:29] cbx_1__1__103_chanx_right_out;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__104_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__104_ccff_tail;
  wire [0:29] cbx_1__1__104_chanx_left_out;
  wire [0:29] cbx_1__1__104_chanx_right_out;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__105_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__105_ccff_tail;
  wire [0:29] cbx_1__1__105_chanx_left_out;
  wire [0:29] cbx_1__1__105_chanx_right_out;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__106_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__106_ccff_tail;
  wire [0:29] cbx_1__1__106_chanx_left_out;
  wire [0:29] cbx_1__1__106_chanx_right_out;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__107_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__107_ccff_tail;
  wire [0:29] cbx_1__1__107_chanx_left_out;
  wire [0:29] cbx_1__1__107_chanx_right_out;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__108_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__108_ccff_tail;
  wire [0:29] cbx_1__1__108_chanx_left_out;
  wire [0:29] cbx_1__1__108_chanx_right_out;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__109_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__109_ccff_tail;
  wire [0:29] cbx_1__1__109_chanx_left_out;
  wire [0:29] cbx_1__1__109_chanx_right_out;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__10_ccff_tail;
  wire [0:29] cbx_1__1__10_chanx_left_out;
  wire [0:29] cbx_1__1__10_chanx_right_out;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__110_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__110_ccff_tail;
  wire [0:29] cbx_1__1__110_chanx_left_out;
  wire [0:29] cbx_1__1__110_chanx_right_out;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__111_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__111_ccff_tail;
  wire [0:29] cbx_1__1__111_chanx_left_out;
  wire [0:29] cbx_1__1__111_chanx_right_out;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__112_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__112_ccff_tail;
  wire [0:29] cbx_1__1__112_chanx_left_out;
  wire [0:29] cbx_1__1__112_chanx_right_out;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__113_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__113_ccff_tail;
  wire [0:29] cbx_1__1__113_chanx_left_out;
  wire [0:29] cbx_1__1__113_chanx_right_out;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__114_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__114_ccff_tail;
  wire [0:29] cbx_1__1__114_chanx_left_out;
  wire [0:29] cbx_1__1__114_chanx_right_out;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__115_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__115_ccff_tail;
  wire [0:29] cbx_1__1__115_chanx_left_out;
  wire [0:29] cbx_1__1__115_chanx_right_out;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__116_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__116_ccff_tail;
  wire [0:29] cbx_1__1__116_chanx_left_out;
  wire [0:29] cbx_1__1__116_chanx_right_out;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__117_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__117_ccff_tail;
  wire [0:29] cbx_1__1__117_chanx_left_out;
  wire [0:29] cbx_1__1__117_chanx_right_out;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__118_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__118_ccff_tail;
  wire [0:29] cbx_1__1__118_chanx_left_out;
  wire [0:29] cbx_1__1__118_chanx_right_out;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__119_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__119_ccff_tail;
  wire [0:29] cbx_1__1__119_chanx_left_out;
  wire [0:29] cbx_1__1__119_chanx_right_out;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__11_ccff_tail;
  wire [0:29] cbx_1__1__11_chanx_left_out;
  wire [0:29] cbx_1__1__11_chanx_right_out;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__120_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__120_ccff_tail;
  wire [0:29] cbx_1__1__120_chanx_left_out;
  wire [0:29] cbx_1__1__120_chanx_right_out;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__121_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__121_ccff_tail;
  wire [0:29] cbx_1__1__121_chanx_left_out;
  wire [0:29] cbx_1__1__121_chanx_right_out;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__122_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__122_ccff_tail;
  wire [0:29] cbx_1__1__122_chanx_left_out;
  wire [0:29] cbx_1__1__122_chanx_right_out;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__123_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__123_ccff_tail;
  wire [0:29] cbx_1__1__123_chanx_left_out;
  wire [0:29] cbx_1__1__123_chanx_right_out;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__124_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__124_ccff_tail;
  wire [0:29] cbx_1__1__124_chanx_left_out;
  wire [0:29] cbx_1__1__124_chanx_right_out;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__125_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__125_ccff_tail;
  wire [0:29] cbx_1__1__125_chanx_left_out;
  wire [0:29] cbx_1__1__125_chanx_right_out;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__126_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__126_ccff_tail;
  wire [0:29] cbx_1__1__126_chanx_left_out;
  wire [0:29] cbx_1__1__126_chanx_right_out;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__127_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__127_ccff_tail;
  wire [0:29] cbx_1__1__127_chanx_left_out;
  wire [0:29] cbx_1__1__127_chanx_right_out;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__128_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__128_ccff_tail;
  wire [0:29] cbx_1__1__128_chanx_left_out;
  wire [0:29] cbx_1__1__128_chanx_right_out;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__129_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__129_ccff_tail;
  wire [0:29] cbx_1__1__129_chanx_left_out;
  wire [0:29] cbx_1__1__129_chanx_right_out;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__12_ccff_tail;
  wire [0:29] cbx_1__1__12_chanx_left_out;
  wire [0:29] cbx_1__1__12_chanx_right_out;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__130_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__130_ccff_tail;
  wire [0:29] cbx_1__1__130_chanx_left_out;
  wire [0:29] cbx_1__1__130_chanx_right_out;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__131_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__131_ccff_tail;
  wire [0:29] cbx_1__1__131_chanx_left_out;
  wire [0:29] cbx_1__1__131_chanx_right_out;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__13_ccff_tail;
  wire [0:29] cbx_1__1__13_chanx_left_out;
  wire [0:29] cbx_1__1__13_chanx_right_out;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__14_ccff_tail;
  wire [0:29] cbx_1__1__14_chanx_left_out;
  wire [0:29] cbx_1__1__14_chanx_right_out;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__15_ccff_tail;
  wire [0:29] cbx_1__1__15_chanx_left_out;
  wire [0:29] cbx_1__1__15_chanx_right_out;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__16_ccff_tail;
  wire [0:29] cbx_1__1__16_chanx_left_out;
  wire [0:29] cbx_1__1__16_chanx_right_out;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__17_ccff_tail;
  wire [0:29] cbx_1__1__17_chanx_left_out;
  wire [0:29] cbx_1__1__17_chanx_right_out;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__18_ccff_tail;
  wire [0:29] cbx_1__1__18_chanx_left_out;
  wire [0:29] cbx_1__1__18_chanx_right_out;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__19_ccff_tail;
  wire [0:29] cbx_1__1__19_chanx_left_out;
  wire [0:29] cbx_1__1__19_chanx_right_out;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__1_ccff_tail;
  wire [0:29] cbx_1__1__1_chanx_left_out;
  wire [0:29] cbx_1__1__1_chanx_right_out;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__20_ccff_tail;
  wire [0:29] cbx_1__1__20_chanx_left_out;
  wire [0:29] cbx_1__1__20_chanx_right_out;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__21_ccff_tail;
  wire [0:29] cbx_1__1__21_chanx_left_out;
  wire [0:29] cbx_1__1__21_chanx_right_out;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__22_ccff_tail;
  wire [0:29] cbx_1__1__22_chanx_left_out;
  wire [0:29] cbx_1__1__22_chanx_right_out;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__23_ccff_tail;
  wire [0:29] cbx_1__1__23_chanx_left_out;
  wire [0:29] cbx_1__1__23_chanx_right_out;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__24_ccff_tail;
  wire [0:29] cbx_1__1__24_chanx_left_out;
  wire [0:29] cbx_1__1__24_chanx_right_out;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__25_ccff_tail;
  wire [0:29] cbx_1__1__25_chanx_left_out;
  wire [0:29] cbx_1__1__25_chanx_right_out;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__26_ccff_tail;
  wire [0:29] cbx_1__1__26_chanx_left_out;
  wire [0:29] cbx_1__1__26_chanx_right_out;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__27_ccff_tail;
  wire [0:29] cbx_1__1__27_chanx_left_out;
  wire [0:29] cbx_1__1__27_chanx_right_out;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__28_ccff_tail;
  wire [0:29] cbx_1__1__28_chanx_left_out;
  wire [0:29] cbx_1__1__28_chanx_right_out;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__29_ccff_tail;
  wire [0:29] cbx_1__1__29_chanx_left_out;
  wire [0:29] cbx_1__1__29_chanx_right_out;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__2_ccff_tail;
  wire [0:29] cbx_1__1__2_chanx_left_out;
  wire [0:29] cbx_1__1__2_chanx_right_out;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__30_ccff_tail;
  wire [0:29] cbx_1__1__30_chanx_left_out;
  wire [0:29] cbx_1__1__30_chanx_right_out;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__31_ccff_tail;
  wire [0:29] cbx_1__1__31_chanx_left_out;
  wire [0:29] cbx_1__1__31_chanx_right_out;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__32_ccff_tail;
  wire [0:29] cbx_1__1__32_chanx_left_out;
  wire [0:29] cbx_1__1__32_chanx_right_out;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__33_ccff_tail;
  wire [0:29] cbx_1__1__33_chanx_left_out;
  wire [0:29] cbx_1__1__33_chanx_right_out;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__34_ccff_tail;
  wire [0:29] cbx_1__1__34_chanx_left_out;
  wire [0:29] cbx_1__1__34_chanx_right_out;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__35_ccff_tail;
  wire [0:29] cbx_1__1__35_chanx_left_out;
  wire [0:29] cbx_1__1__35_chanx_right_out;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__36_ccff_tail;
  wire [0:29] cbx_1__1__36_chanx_left_out;
  wire [0:29] cbx_1__1__36_chanx_right_out;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__37_ccff_tail;
  wire [0:29] cbx_1__1__37_chanx_left_out;
  wire [0:29] cbx_1__1__37_chanx_right_out;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__38_ccff_tail;
  wire [0:29] cbx_1__1__38_chanx_left_out;
  wire [0:29] cbx_1__1__38_chanx_right_out;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__39_ccff_tail;
  wire [0:29] cbx_1__1__39_chanx_left_out;
  wire [0:29] cbx_1__1__39_chanx_right_out;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__3_ccff_tail;
  wire [0:29] cbx_1__1__3_chanx_left_out;
  wire [0:29] cbx_1__1__3_chanx_right_out;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__40_ccff_tail;
  wire [0:29] cbx_1__1__40_chanx_left_out;
  wire [0:29] cbx_1__1__40_chanx_right_out;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__41_ccff_tail;
  wire [0:29] cbx_1__1__41_chanx_left_out;
  wire [0:29] cbx_1__1__41_chanx_right_out;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__42_ccff_tail;
  wire [0:29] cbx_1__1__42_chanx_left_out;
  wire [0:29] cbx_1__1__42_chanx_right_out;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__43_ccff_tail;
  wire [0:29] cbx_1__1__43_chanx_left_out;
  wire [0:29] cbx_1__1__43_chanx_right_out;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__44_ccff_tail;
  wire [0:29] cbx_1__1__44_chanx_left_out;
  wire [0:29] cbx_1__1__44_chanx_right_out;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__45_ccff_tail;
  wire [0:29] cbx_1__1__45_chanx_left_out;
  wire [0:29] cbx_1__1__45_chanx_right_out;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__46_ccff_tail;
  wire [0:29] cbx_1__1__46_chanx_left_out;
  wire [0:29] cbx_1__1__46_chanx_right_out;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__47_ccff_tail;
  wire [0:29] cbx_1__1__47_chanx_left_out;
  wire [0:29] cbx_1__1__47_chanx_right_out;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__48_ccff_tail;
  wire [0:29] cbx_1__1__48_chanx_left_out;
  wire [0:29] cbx_1__1__48_chanx_right_out;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__49_ccff_tail;
  wire [0:29] cbx_1__1__49_chanx_left_out;
  wire [0:29] cbx_1__1__49_chanx_right_out;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__4_ccff_tail;
  wire [0:29] cbx_1__1__4_chanx_left_out;
  wire [0:29] cbx_1__1__4_chanx_right_out;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__50_ccff_tail;
  wire [0:29] cbx_1__1__50_chanx_left_out;
  wire [0:29] cbx_1__1__50_chanx_right_out;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__51_ccff_tail;
  wire [0:29] cbx_1__1__51_chanx_left_out;
  wire [0:29] cbx_1__1__51_chanx_right_out;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__52_ccff_tail;
  wire [0:29] cbx_1__1__52_chanx_left_out;
  wire [0:29] cbx_1__1__52_chanx_right_out;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__53_ccff_tail;
  wire [0:29] cbx_1__1__53_chanx_left_out;
  wire [0:29] cbx_1__1__53_chanx_right_out;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__54_ccff_tail;
  wire [0:29] cbx_1__1__54_chanx_left_out;
  wire [0:29] cbx_1__1__54_chanx_right_out;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__55_ccff_tail;
  wire [0:29] cbx_1__1__55_chanx_left_out;
  wire [0:29] cbx_1__1__55_chanx_right_out;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__56_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__56_ccff_tail;
  wire [0:29] cbx_1__1__56_chanx_left_out;
  wire [0:29] cbx_1__1__56_chanx_right_out;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__57_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__57_ccff_tail;
  wire [0:29] cbx_1__1__57_chanx_left_out;
  wire [0:29] cbx_1__1__57_chanx_right_out;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__58_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__58_ccff_tail;
  wire [0:29] cbx_1__1__58_chanx_left_out;
  wire [0:29] cbx_1__1__58_chanx_right_out;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__59_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__59_ccff_tail;
  wire [0:29] cbx_1__1__59_chanx_left_out;
  wire [0:29] cbx_1__1__59_chanx_right_out;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__5_ccff_tail;
  wire [0:29] cbx_1__1__5_chanx_left_out;
  wire [0:29] cbx_1__1__5_chanx_right_out;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__60_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__60_ccff_tail;
  wire [0:29] cbx_1__1__60_chanx_left_out;
  wire [0:29] cbx_1__1__60_chanx_right_out;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__61_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__61_ccff_tail;
  wire [0:29] cbx_1__1__61_chanx_left_out;
  wire [0:29] cbx_1__1__61_chanx_right_out;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__62_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__62_ccff_tail;
  wire [0:29] cbx_1__1__62_chanx_left_out;
  wire [0:29] cbx_1__1__62_chanx_right_out;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__63_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__63_ccff_tail;
  wire [0:29] cbx_1__1__63_chanx_left_out;
  wire [0:29] cbx_1__1__63_chanx_right_out;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__64_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__64_ccff_tail;
  wire [0:29] cbx_1__1__64_chanx_left_out;
  wire [0:29] cbx_1__1__64_chanx_right_out;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__65_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__65_ccff_tail;
  wire [0:29] cbx_1__1__65_chanx_left_out;
  wire [0:29] cbx_1__1__65_chanx_right_out;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__66_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__66_ccff_tail;
  wire [0:29] cbx_1__1__66_chanx_left_out;
  wire [0:29] cbx_1__1__66_chanx_right_out;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__67_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__67_ccff_tail;
  wire [0:29] cbx_1__1__67_chanx_left_out;
  wire [0:29] cbx_1__1__67_chanx_right_out;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__68_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__68_ccff_tail;
  wire [0:29] cbx_1__1__68_chanx_left_out;
  wire [0:29] cbx_1__1__68_chanx_right_out;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__69_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__69_ccff_tail;
  wire [0:29] cbx_1__1__69_chanx_left_out;
  wire [0:29] cbx_1__1__69_chanx_right_out;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__6_ccff_tail;
  wire [0:29] cbx_1__1__6_chanx_left_out;
  wire [0:29] cbx_1__1__6_chanx_right_out;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__70_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__70_ccff_tail;
  wire [0:29] cbx_1__1__70_chanx_left_out;
  wire [0:29] cbx_1__1__70_chanx_right_out;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__71_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__71_ccff_tail;
  wire [0:29] cbx_1__1__71_chanx_left_out;
  wire [0:29] cbx_1__1__71_chanx_right_out;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__72_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__72_ccff_tail;
  wire [0:29] cbx_1__1__72_chanx_left_out;
  wire [0:29] cbx_1__1__72_chanx_right_out;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__73_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__73_ccff_tail;
  wire [0:29] cbx_1__1__73_chanx_left_out;
  wire [0:29] cbx_1__1__73_chanx_right_out;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__74_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__74_ccff_tail;
  wire [0:29] cbx_1__1__74_chanx_left_out;
  wire [0:29] cbx_1__1__74_chanx_right_out;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__75_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__75_ccff_tail;
  wire [0:29] cbx_1__1__75_chanx_left_out;
  wire [0:29] cbx_1__1__75_chanx_right_out;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__76_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__76_ccff_tail;
  wire [0:29] cbx_1__1__76_chanx_left_out;
  wire [0:29] cbx_1__1__76_chanx_right_out;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__77_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__77_ccff_tail;
  wire [0:29] cbx_1__1__77_chanx_left_out;
  wire [0:29] cbx_1__1__77_chanx_right_out;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__78_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__78_ccff_tail;
  wire [0:29] cbx_1__1__78_chanx_left_out;
  wire [0:29] cbx_1__1__78_chanx_right_out;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__79_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__79_ccff_tail;
  wire [0:29] cbx_1__1__79_chanx_left_out;
  wire [0:29] cbx_1__1__79_chanx_right_out;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__7_ccff_tail;
  wire [0:29] cbx_1__1__7_chanx_left_out;
  wire [0:29] cbx_1__1__7_chanx_right_out;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__80_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__80_ccff_tail;
  wire [0:29] cbx_1__1__80_chanx_left_out;
  wire [0:29] cbx_1__1__80_chanx_right_out;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__81_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__81_ccff_tail;
  wire [0:29] cbx_1__1__81_chanx_left_out;
  wire [0:29] cbx_1__1__81_chanx_right_out;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__82_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__82_ccff_tail;
  wire [0:29] cbx_1__1__82_chanx_left_out;
  wire [0:29] cbx_1__1__82_chanx_right_out;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__83_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__83_ccff_tail;
  wire [0:29] cbx_1__1__83_chanx_left_out;
  wire [0:29] cbx_1__1__83_chanx_right_out;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__84_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__84_ccff_tail;
  wire [0:29] cbx_1__1__84_chanx_left_out;
  wire [0:29] cbx_1__1__84_chanx_right_out;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__85_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__85_ccff_tail;
  wire [0:29] cbx_1__1__85_chanx_left_out;
  wire [0:29] cbx_1__1__85_chanx_right_out;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__86_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__86_ccff_tail;
  wire [0:29] cbx_1__1__86_chanx_left_out;
  wire [0:29] cbx_1__1__86_chanx_right_out;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__87_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__87_ccff_tail;
  wire [0:29] cbx_1__1__87_chanx_left_out;
  wire [0:29] cbx_1__1__87_chanx_right_out;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__88_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__88_ccff_tail;
  wire [0:29] cbx_1__1__88_chanx_left_out;
  wire [0:29] cbx_1__1__88_chanx_right_out;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__89_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__89_ccff_tail;
  wire [0:29] cbx_1__1__89_chanx_left_out;
  wire [0:29] cbx_1__1__89_chanx_right_out;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__8_ccff_tail;
  wire [0:29] cbx_1__1__8_chanx_left_out;
  wire [0:29] cbx_1__1__8_chanx_right_out;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__90_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__90_ccff_tail;
  wire [0:29] cbx_1__1__90_chanx_left_out;
  wire [0:29] cbx_1__1__90_chanx_right_out;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__91_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__91_ccff_tail;
  wire [0:29] cbx_1__1__91_chanx_left_out;
  wire [0:29] cbx_1__1__91_chanx_right_out;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__92_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__92_ccff_tail;
  wire [0:29] cbx_1__1__92_chanx_left_out;
  wire [0:29] cbx_1__1__92_chanx_right_out;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__93_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__93_ccff_tail;
  wire [0:29] cbx_1__1__93_chanx_left_out;
  wire [0:29] cbx_1__1__93_chanx_right_out;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__94_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__94_ccff_tail;
  wire [0:29] cbx_1__1__94_chanx_left_out;
  wire [0:29] cbx_1__1__94_chanx_right_out;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__95_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__95_ccff_tail;
  wire [0:29] cbx_1__1__95_chanx_left_out;
  wire [0:29] cbx_1__1__95_chanx_right_out;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__96_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__96_ccff_tail;
  wire [0:29] cbx_1__1__96_chanx_left_out;
  wire [0:29] cbx_1__1__96_chanx_right_out;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__97_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__97_ccff_tail;
  wire [0:29] cbx_1__1__97_chanx_left_out;
  wire [0:29] cbx_1__1__97_chanx_right_out;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__98_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__98_ccff_tail;
  wire [0:29] cbx_1__1__98_chanx_left_out;
  wire [0:29] cbx_1__1__98_chanx_right_out;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__99_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__99_ccff_tail;
  wire [0:29] cbx_1__1__99_chanx_left_out;
  wire [0:29] cbx_1__1__99_chanx_right_out;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__9_ccff_tail;
  wire [0:29] cbx_1__1__9_chanx_left_out;
  wire [0:29] cbx_1__1__9_chanx_right_out;
  wire [0:0] cby_0__1__0_ccff_tail;
  wire [0:29] cby_0__1__0_chany_bottom_out;
  wire [0:29] cby_0__1__0_chany_top_out;
  wire [0:0] cby_0__1__0_left_grid_pin_0_;
  wire [0:0] cby_0__1__10_ccff_tail;
  wire [0:29] cby_0__1__10_chany_bottom_out;
  wire [0:29] cby_0__1__10_chany_top_out;
  wire [0:0] cby_0__1__10_left_grid_pin_0_;
  wire [0:0] cby_0__1__11_ccff_tail;
  wire [0:29] cby_0__1__11_chany_bottom_out;
  wire [0:29] cby_0__1__11_chany_top_out;
  wire [0:0] cby_0__1__11_left_grid_pin_0_;
  wire [0:0] cby_0__1__1_ccff_tail;
  wire [0:29] cby_0__1__1_chany_bottom_out;
  wire [0:29] cby_0__1__1_chany_top_out;
  wire [0:0] cby_0__1__1_left_grid_pin_0_;
  wire [0:0] cby_0__1__2_ccff_tail;
  wire [0:29] cby_0__1__2_chany_bottom_out;
  wire [0:29] cby_0__1__2_chany_top_out;
  wire [0:0] cby_0__1__2_left_grid_pin_0_;
  wire [0:0] cby_0__1__3_ccff_tail;
  wire [0:29] cby_0__1__3_chany_bottom_out;
  wire [0:29] cby_0__1__3_chany_top_out;
  wire [0:0] cby_0__1__3_left_grid_pin_0_;
  wire [0:0] cby_0__1__4_ccff_tail;
  wire [0:29] cby_0__1__4_chany_bottom_out;
  wire [0:29] cby_0__1__4_chany_top_out;
  wire [0:0] cby_0__1__4_left_grid_pin_0_;
  wire [0:0] cby_0__1__5_ccff_tail;
  wire [0:29] cby_0__1__5_chany_bottom_out;
  wire [0:29] cby_0__1__5_chany_top_out;
  wire [0:0] cby_0__1__5_left_grid_pin_0_;
  wire [0:0] cby_0__1__6_ccff_tail;
  wire [0:29] cby_0__1__6_chany_bottom_out;
  wire [0:29] cby_0__1__6_chany_top_out;
  wire [0:0] cby_0__1__6_left_grid_pin_0_;
  wire [0:0] cby_0__1__7_ccff_tail;
  wire [0:29] cby_0__1__7_chany_bottom_out;
  wire [0:29] cby_0__1__7_chany_top_out;
  wire [0:0] cby_0__1__7_left_grid_pin_0_;
  wire [0:0] cby_0__1__8_ccff_tail;
  wire [0:29] cby_0__1__8_chany_bottom_out;
  wire [0:29] cby_0__1__8_chany_top_out;
  wire [0:0] cby_0__1__8_left_grid_pin_0_;
  wire [0:0] cby_0__1__9_ccff_tail;
  wire [0:29] cby_0__1__9_chany_bottom_out;
  wire [0:29] cby_0__1__9_chany_top_out;
  wire [0:0] cby_0__1__9_left_grid_pin_0_;
  wire [0:0] cby_12__1__0_ccff_tail;
  wire [0:29] cby_12__1__0_chany_bottom_out;
  wire [0:29] cby_12__1__0_chany_top_out;
  wire [0:0] cby_12__1__0_left_grid_pin_16_;
  wire [0:0] cby_12__1__0_left_grid_pin_17_;
  wire [0:0] cby_12__1__0_left_grid_pin_18_;
  wire [0:0] cby_12__1__0_left_grid_pin_19_;
  wire [0:0] cby_12__1__0_left_grid_pin_20_;
  wire [0:0] cby_12__1__0_left_grid_pin_21_;
  wire [0:0] cby_12__1__0_left_grid_pin_22_;
  wire [0:0] cby_12__1__0_left_grid_pin_23_;
  wire [0:0] cby_12__1__0_left_grid_pin_24_;
  wire [0:0] cby_12__1__0_left_grid_pin_25_;
  wire [0:0] cby_12__1__0_left_grid_pin_26_;
  wire [0:0] cby_12__1__0_left_grid_pin_27_;
  wire [0:0] cby_12__1__0_left_grid_pin_28_;
  wire [0:0] cby_12__1__0_left_grid_pin_29_;
  wire [0:0] cby_12__1__0_left_grid_pin_30_;
  wire [0:0] cby_12__1__0_left_grid_pin_31_;
  wire [0:0] cby_12__1__0_right_grid_pin_0_;
  wire [0:0] cby_12__1__10_ccff_tail;
  wire [0:29] cby_12__1__10_chany_bottom_out;
  wire [0:29] cby_12__1__10_chany_top_out;
  wire [0:0] cby_12__1__10_left_grid_pin_16_;
  wire [0:0] cby_12__1__10_left_grid_pin_17_;
  wire [0:0] cby_12__1__10_left_grid_pin_18_;
  wire [0:0] cby_12__1__10_left_grid_pin_19_;
  wire [0:0] cby_12__1__10_left_grid_pin_20_;
  wire [0:0] cby_12__1__10_left_grid_pin_21_;
  wire [0:0] cby_12__1__10_left_grid_pin_22_;
  wire [0:0] cby_12__1__10_left_grid_pin_23_;
  wire [0:0] cby_12__1__10_left_grid_pin_24_;
  wire [0:0] cby_12__1__10_left_grid_pin_25_;
  wire [0:0] cby_12__1__10_left_grid_pin_26_;
  wire [0:0] cby_12__1__10_left_grid_pin_27_;
  wire [0:0] cby_12__1__10_left_grid_pin_28_;
  wire [0:0] cby_12__1__10_left_grid_pin_29_;
  wire [0:0] cby_12__1__10_left_grid_pin_30_;
  wire [0:0] cby_12__1__10_left_grid_pin_31_;
  wire [0:0] cby_12__1__10_right_grid_pin_0_;
  wire [0:0] cby_12__1__11_ccff_tail;
  wire [0:29] cby_12__1__11_chany_bottom_out;
  wire [0:29] cby_12__1__11_chany_top_out;
  wire [0:0] cby_12__1__11_left_grid_pin_16_;
  wire [0:0] cby_12__1__11_left_grid_pin_17_;
  wire [0:0] cby_12__1__11_left_grid_pin_18_;
  wire [0:0] cby_12__1__11_left_grid_pin_19_;
  wire [0:0] cby_12__1__11_left_grid_pin_20_;
  wire [0:0] cby_12__1__11_left_grid_pin_21_;
  wire [0:0] cby_12__1__11_left_grid_pin_22_;
  wire [0:0] cby_12__1__11_left_grid_pin_23_;
  wire [0:0] cby_12__1__11_left_grid_pin_24_;
  wire [0:0] cby_12__1__11_left_grid_pin_25_;
  wire [0:0] cby_12__1__11_left_grid_pin_26_;
  wire [0:0] cby_12__1__11_left_grid_pin_27_;
  wire [0:0] cby_12__1__11_left_grid_pin_28_;
  wire [0:0] cby_12__1__11_left_grid_pin_29_;
  wire [0:0] cby_12__1__11_left_grid_pin_30_;
  wire [0:0] cby_12__1__11_left_grid_pin_31_;
  wire [0:0] cby_12__1__11_right_grid_pin_0_;
  wire [0:0] cby_12__1__1_ccff_tail;
  wire [0:29] cby_12__1__1_chany_bottom_out;
  wire [0:29] cby_12__1__1_chany_top_out;
  wire [0:0] cby_12__1__1_left_grid_pin_16_;
  wire [0:0] cby_12__1__1_left_grid_pin_17_;
  wire [0:0] cby_12__1__1_left_grid_pin_18_;
  wire [0:0] cby_12__1__1_left_grid_pin_19_;
  wire [0:0] cby_12__1__1_left_grid_pin_20_;
  wire [0:0] cby_12__1__1_left_grid_pin_21_;
  wire [0:0] cby_12__1__1_left_grid_pin_22_;
  wire [0:0] cby_12__1__1_left_grid_pin_23_;
  wire [0:0] cby_12__1__1_left_grid_pin_24_;
  wire [0:0] cby_12__1__1_left_grid_pin_25_;
  wire [0:0] cby_12__1__1_left_grid_pin_26_;
  wire [0:0] cby_12__1__1_left_grid_pin_27_;
  wire [0:0] cby_12__1__1_left_grid_pin_28_;
  wire [0:0] cby_12__1__1_left_grid_pin_29_;
  wire [0:0] cby_12__1__1_left_grid_pin_30_;
  wire [0:0] cby_12__1__1_left_grid_pin_31_;
  wire [0:0] cby_12__1__1_right_grid_pin_0_;
  wire [0:0] cby_12__1__2_ccff_tail;
  wire [0:29] cby_12__1__2_chany_bottom_out;
  wire [0:29] cby_12__1__2_chany_top_out;
  wire [0:0] cby_12__1__2_left_grid_pin_16_;
  wire [0:0] cby_12__1__2_left_grid_pin_17_;
  wire [0:0] cby_12__1__2_left_grid_pin_18_;
  wire [0:0] cby_12__1__2_left_grid_pin_19_;
  wire [0:0] cby_12__1__2_left_grid_pin_20_;
  wire [0:0] cby_12__1__2_left_grid_pin_21_;
  wire [0:0] cby_12__1__2_left_grid_pin_22_;
  wire [0:0] cby_12__1__2_left_grid_pin_23_;
  wire [0:0] cby_12__1__2_left_grid_pin_24_;
  wire [0:0] cby_12__1__2_left_grid_pin_25_;
  wire [0:0] cby_12__1__2_left_grid_pin_26_;
  wire [0:0] cby_12__1__2_left_grid_pin_27_;
  wire [0:0] cby_12__1__2_left_grid_pin_28_;
  wire [0:0] cby_12__1__2_left_grid_pin_29_;
  wire [0:0] cby_12__1__2_left_grid_pin_30_;
  wire [0:0] cby_12__1__2_left_grid_pin_31_;
  wire [0:0] cby_12__1__2_right_grid_pin_0_;
  wire [0:0] cby_12__1__3_ccff_tail;
  wire [0:29] cby_12__1__3_chany_bottom_out;
  wire [0:29] cby_12__1__3_chany_top_out;
  wire [0:0] cby_12__1__3_left_grid_pin_16_;
  wire [0:0] cby_12__1__3_left_grid_pin_17_;
  wire [0:0] cby_12__1__3_left_grid_pin_18_;
  wire [0:0] cby_12__1__3_left_grid_pin_19_;
  wire [0:0] cby_12__1__3_left_grid_pin_20_;
  wire [0:0] cby_12__1__3_left_grid_pin_21_;
  wire [0:0] cby_12__1__3_left_grid_pin_22_;
  wire [0:0] cby_12__1__3_left_grid_pin_23_;
  wire [0:0] cby_12__1__3_left_grid_pin_24_;
  wire [0:0] cby_12__1__3_left_grid_pin_25_;
  wire [0:0] cby_12__1__3_left_grid_pin_26_;
  wire [0:0] cby_12__1__3_left_grid_pin_27_;
  wire [0:0] cby_12__1__3_left_grid_pin_28_;
  wire [0:0] cby_12__1__3_left_grid_pin_29_;
  wire [0:0] cby_12__1__3_left_grid_pin_30_;
  wire [0:0] cby_12__1__3_left_grid_pin_31_;
  wire [0:0] cby_12__1__3_right_grid_pin_0_;
  wire [0:0] cby_12__1__4_ccff_tail;
  wire [0:29] cby_12__1__4_chany_bottom_out;
  wire [0:29] cby_12__1__4_chany_top_out;
  wire [0:0] cby_12__1__4_left_grid_pin_16_;
  wire [0:0] cby_12__1__4_left_grid_pin_17_;
  wire [0:0] cby_12__1__4_left_grid_pin_18_;
  wire [0:0] cby_12__1__4_left_grid_pin_19_;
  wire [0:0] cby_12__1__4_left_grid_pin_20_;
  wire [0:0] cby_12__1__4_left_grid_pin_21_;
  wire [0:0] cby_12__1__4_left_grid_pin_22_;
  wire [0:0] cby_12__1__4_left_grid_pin_23_;
  wire [0:0] cby_12__1__4_left_grid_pin_24_;
  wire [0:0] cby_12__1__4_left_grid_pin_25_;
  wire [0:0] cby_12__1__4_left_grid_pin_26_;
  wire [0:0] cby_12__1__4_left_grid_pin_27_;
  wire [0:0] cby_12__1__4_left_grid_pin_28_;
  wire [0:0] cby_12__1__4_left_grid_pin_29_;
  wire [0:0] cby_12__1__4_left_grid_pin_30_;
  wire [0:0] cby_12__1__4_left_grid_pin_31_;
  wire [0:0] cby_12__1__4_right_grid_pin_0_;
  wire [0:0] cby_12__1__5_ccff_tail;
  wire [0:29] cby_12__1__5_chany_bottom_out;
  wire [0:29] cby_12__1__5_chany_top_out;
  wire [0:0] cby_12__1__5_left_grid_pin_16_;
  wire [0:0] cby_12__1__5_left_grid_pin_17_;
  wire [0:0] cby_12__1__5_left_grid_pin_18_;
  wire [0:0] cby_12__1__5_left_grid_pin_19_;
  wire [0:0] cby_12__1__5_left_grid_pin_20_;
  wire [0:0] cby_12__1__5_left_grid_pin_21_;
  wire [0:0] cby_12__1__5_left_grid_pin_22_;
  wire [0:0] cby_12__1__5_left_grid_pin_23_;
  wire [0:0] cby_12__1__5_left_grid_pin_24_;
  wire [0:0] cby_12__1__5_left_grid_pin_25_;
  wire [0:0] cby_12__1__5_left_grid_pin_26_;
  wire [0:0] cby_12__1__5_left_grid_pin_27_;
  wire [0:0] cby_12__1__5_left_grid_pin_28_;
  wire [0:0] cby_12__1__5_left_grid_pin_29_;
  wire [0:0] cby_12__1__5_left_grid_pin_30_;
  wire [0:0] cby_12__1__5_left_grid_pin_31_;
  wire [0:0] cby_12__1__5_right_grid_pin_0_;
  wire [0:0] cby_12__1__6_ccff_tail;
  wire [0:29] cby_12__1__6_chany_bottom_out;
  wire [0:29] cby_12__1__6_chany_top_out;
  wire [0:0] cby_12__1__6_left_grid_pin_16_;
  wire [0:0] cby_12__1__6_left_grid_pin_17_;
  wire [0:0] cby_12__1__6_left_grid_pin_18_;
  wire [0:0] cby_12__1__6_left_grid_pin_19_;
  wire [0:0] cby_12__1__6_left_grid_pin_20_;
  wire [0:0] cby_12__1__6_left_grid_pin_21_;
  wire [0:0] cby_12__1__6_left_grid_pin_22_;
  wire [0:0] cby_12__1__6_left_grid_pin_23_;
  wire [0:0] cby_12__1__6_left_grid_pin_24_;
  wire [0:0] cby_12__1__6_left_grid_pin_25_;
  wire [0:0] cby_12__1__6_left_grid_pin_26_;
  wire [0:0] cby_12__1__6_left_grid_pin_27_;
  wire [0:0] cby_12__1__6_left_grid_pin_28_;
  wire [0:0] cby_12__1__6_left_grid_pin_29_;
  wire [0:0] cby_12__1__6_left_grid_pin_30_;
  wire [0:0] cby_12__1__6_left_grid_pin_31_;
  wire [0:0] cby_12__1__6_right_grid_pin_0_;
  wire [0:0] cby_12__1__7_ccff_tail;
  wire [0:29] cby_12__1__7_chany_bottom_out;
  wire [0:29] cby_12__1__7_chany_top_out;
  wire [0:0] cby_12__1__7_left_grid_pin_16_;
  wire [0:0] cby_12__1__7_left_grid_pin_17_;
  wire [0:0] cby_12__1__7_left_grid_pin_18_;
  wire [0:0] cby_12__1__7_left_grid_pin_19_;
  wire [0:0] cby_12__1__7_left_grid_pin_20_;
  wire [0:0] cby_12__1__7_left_grid_pin_21_;
  wire [0:0] cby_12__1__7_left_grid_pin_22_;
  wire [0:0] cby_12__1__7_left_grid_pin_23_;
  wire [0:0] cby_12__1__7_left_grid_pin_24_;
  wire [0:0] cby_12__1__7_left_grid_pin_25_;
  wire [0:0] cby_12__1__7_left_grid_pin_26_;
  wire [0:0] cby_12__1__7_left_grid_pin_27_;
  wire [0:0] cby_12__1__7_left_grid_pin_28_;
  wire [0:0] cby_12__1__7_left_grid_pin_29_;
  wire [0:0] cby_12__1__7_left_grid_pin_30_;
  wire [0:0] cby_12__1__7_left_grid_pin_31_;
  wire [0:0] cby_12__1__7_right_grid_pin_0_;
  wire [0:0] cby_12__1__8_ccff_tail;
  wire [0:29] cby_12__1__8_chany_bottom_out;
  wire [0:29] cby_12__1__8_chany_top_out;
  wire [0:0] cby_12__1__8_left_grid_pin_16_;
  wire [0:0] cby_12__1__8_left_grid_pin_17_;
  wire [0:0] cby_12__1__8_left_grid_pin_18_;
  wire [0:0] cby_12__1__8_left_grid_pin_19_;
  wire [0:0] cby_12__1__8_left_grid_pin_20_;
  wire [0:0] cby_12__1__8_left_grid_pin_21_;
  wire [0:0] cby_12__1__8_left_grid_pin_22_;
  wire [0:0] cby_12__1__8_left_grid_pin_23_;
  wire [0:0] cby_12__1__8_left_grid_pin_24_;
  wire [0:0] cby_12__1__8_left_grid_pin_25_;
  wire [0:0] cby_12__1__8_left_grid_pin_26_;
  wire [0:0] cby_12__1__8_left_grid_pin_27_;
  wire [0:0] cby_12__1__8_left_grid_pin_28_;
  wire [0:0] cby_12__1__8_left_grid_pin_29_;
  wire [0:0] cby_12__1__8_left_grid_pin_30_;
  wire [0:0] cby_12__1__8_left_grid_pin_31_;
  wire [0:0] cby_12__1__8_right_grid_pin_0_;
  wire [0:0] cby_12__1__9_ccff_tail;
  wire [0:29] cby_12__1__9_chany_bottom_out;
  wire [0:29] cby_12__1__9_chany_top_out;
  wire [0:0] cby_12__1__9_left_grid_pin_16_;
  wire [0:0] cby_12__1__9_left_grid_pin_17_;
  wire [0:0] cby_12__1__9_left_grid_pin_18_;
  wire [0:0] cby_12__1__9_left_grid_pin_19_;
  wire [0:0] cby_12__1__9_left_grid_pin_20_;
  wire [0:0] cby_12__1__9_left_grid_pin_21_;
  wire [0:0] cby_12__1__9_left_grid_pin_22_;
  wire [0:0] cby_12__1__9_left_grid_pin_23_;
  wire [0:0] cby_12__1__9_left_grid_pin_24_;
  wire [0:0] cby_12__1__9_left_grid_pin_25_;
  wire [0:0] cby_12__1__9_left_grid_pin_26_;
  wire [0:0] cby_12__1__9_left_grid_pin_27_;
  wire [0:0] cby_12__1__9_left_grid_pin_28_;
  wire [0:0] cby_12__1__9_left_grid_pin_29_;
  wire [0:0] cby_12__1__9_left_grid_pin_30_;
  wire [0:0] cby_12__1__9_left_grid_pin_31_;
  wire [0:0] cby_12__1__9_right_grid_pin_0_;
  wire [0:0] cby_1__1__0_ccff_tail;
  wire [0:29] cby_1__1__0_chany_bottom_out;
  wire [0:29] cby_1__1__0_chany_top_out;
  wire [0:0] cby_1__1__0_left_grid_pin_16_;
  wire [0:0] cby_1__1__0_left_grid_pin_17_;
  wire [0:0] cby_1__1__0_left_grid_pin_18_;
  wire [0:0] cby_1__1__0_left_grid_pin_19_;
  wire [0:0] cby_1__1__0_left_grid_pin_20_;
  wire [0:0] cby_1__1__0_left_grid_pin_21_;
  wire [0:0] cby_1__1__0_left_grid_pin_22_;
  wire [0:0] cby_1__1__0_left_grid_pin_23_;
  wire [0:0] cby_1__1__0_left_grid_pin_24_;
  wire [0:0] cby_1__1__0_left_grid_pin_25_;
  wire [0:0] cby_1__1__0_left_grid_pin_26_;
  wire [0:0] cby_1__1__0_left_grid_pin_27_;
  wire [0:0] cby_1__1__0_left_grid_pin_28_;
  wire [0:0] cby_1__1__0_left_grid_pin_29_;
  wire [0:0] cby_1__1__0_left_grid_pin_30_;
  wire [0:0] cby_1__1__0_left_grid_pin_31_;
  wire [0:0] cby_1__1__100_ccff_tail;
  wire [0:29] cby_1__1__100_chany_bottom_out;
  wire [0:29] cby_1__1__100_chany_top_out;
  wire [0:0] cby_1__1__100_left_grid_pin_16_;
  wire [0:0] cby_1__1__100_left_grid_pin_17_;
  wire [0:0] cby_1__1__100_left_grid_pin_18_;
  wire [0:0] cby_1__1__100_left_grid_pin_19_;
  wire [0:0] cby_1__1__100_left_grid_pin_20_;
  wire [0:0] cby_1__1__100_left_grid_pin_21_;
  wire [0:0] cby_1__1__100_left_grid_pin_22_;
  wire [0:0] cby_1__1__100_left_grid_pin_23_;
  wire [0:0] cby_1__1__100_left_grid_pin_24_;
  wire [0:0] cby_1__1__100_left_grid_pin_25_;
  wire [0:0] cby_1__1__100_left_grid_pin_26_;
  wire [0:0] cby_1__1__100_left_grid_pin_27_;
  wire [0:0] cby_1__1__100_left_grid_pin_28_;
  wire [0:0] cby_1__1__100_left_grid_pin_29_;
  wire [0:0] cby_1__1__100_left_grid_pin_30_;
  wire [0:0] cby_1__1__100_left_grid_pin_31_;
  wire [0:0] cby_1__1__101_ccff_tail;
  wire [0:29] cby_1__1__101_chany_bottom_out;
  wire [0:29] cby_1__1__101_chany_top_out;
  wire [0:0] cby_1__1__101_left_grid_pin_16_;
  wire [0:0] cby_1__1__101_left_grid_pin_17_;
  wire [0:0] cby_1__1__101_left_grid_pin_18_;
  wire [0:0] cby_1__1__101_left_grid_pin_19_;
  wire [0:0] cby_1__1__101_left_grid_pin_20_;
  wire [0:0] cby_1__1__101_left_grid_pin_21_;
  wire [0:0] cby_1__1__101_left_grid_pin_22_;
  wire [0:0] cby_1__1__101_left_grid_pin_23_;
  wire [0:0] cby_1__1__101_left_grid_pin_24_;
  wire [0:0] cby_1__1__101_left_grid_pin_25_;
  wire [0:0] cby_1__1__101_left_grid_pin_26_;
  wire [0:0] cby_1__1__101_left_grid_pin_27_;
  wire [0:0] cby_1__1__101_left_grid_pin_28_;
  wire [0:0] cby_1__1__101_left_grid_pin_29_;
  wire [0:0] cby_1__1__101_left_grid_pin_30_;
  wire [0:0] cby_1__1__101_left_grid_pin_31_;
  wire [0:0] cby_1__1__102_ccff_tail;
  wire [0:29] cby_1__1__102_chany_bottom_out;
  wire [0:29] cby_1__1__102_chany_top_out;
  wire [0:0] cby_1__1__102_left_grid_pin_16_;
  wire [0:0] cby_1__1__102_left_grid_pin_17_;
  wire [0:0] cby_1__1__102_left_grid_pin_18_;
  wire [0:0] cby_1__1__102_left_grid_pin_19_;
  wire [0:0] cby_1__1__102_left_grid_pin_20_;
  wire [0:0] cby_1__1__102_left_grid_pin_21_;
  wire [0:0] cby_1__1__102_left_grid_pin_22_;
  wire [0:0] cby_1__1__102_left_grid_pin_23_;
  wire [0:0] cby_1__1__102_left_grid_pin_24_;
  wire [0:0] cby_1__1__102_left_grid_pin_25_;
  wire [0:0] cby_1__1__102_left_grid_pin_26_;
  wire [0:0] cby_1__1__102_left_grid_pin_27_;
  wire [0:0] cby_1__1__102_left_grid_pin_28_;
  wire [0:0] cby_1__1__102_left_grid_pin_29_;
  wire [0:0] cby_1__1__102_left_grid_pin_30_;
  wire [0:0] cby_1__1__102_left_grid_pin_31_;
  wire [0:0] cby_1__1__103_ccff_tail;
  wire [0:29] cby_1__1__103_chany_bottom_out;
  wire [0:29] cby_1__1__103_chany_top_out;
  wire [0:0] cby_1__1__103_left_grid_pin_16_;
  wire [0:0] cby_1__1__103_left_grid_pin_17_;
  wire [0:0] cby_1__1__103_left_grid_pin_18_;
  wire [0:0] cby_1__1__103_left_grid_pin_19_;
  wire [0:0] cby_1__1__103_left_grid_pin_20_;
  wire [0:0] cby_1__1__103_left_grid_pin_21_;
  wire [0:0] cby_1__1__103_left_grid_pin_22_;
  wire [0:0] cby_1__1__103_left_grid_pin_23_;
  wire [0:0] cby_1__1__103_left_grid_pin_24_;
  wire [0:0] cby_1__1__103_left_grid_pin_25_;
  wire [0:0] cby_1__1__103_left_grid_pin_26_;
  wire [0:0] cby_1__1__103_left_grid_pin_27_;
  wire [0:0] cby_1__1__103_left_grid_pin_28_;
  wire [0:0] cby_1__1__103_left_grid_pin_29_;
  wire [0:0] cby_1__1__103_left_grid_pin_30_;
  wire [0:0] cby_1__1__103_left_grid_pin_31_;
  wire [0:0] cby_1__1__104_ccff_tail;
  wire [0:29] cby_1__1__104_chany_bottom_out;
  wire [0:29] cby_1__1__104_chany_top_out;
  wire [0:0] cby_1__1__104_left_grid_pin_16_;
  wire [0:0] cby_1__1__104_left_grid_pin_17_;
  wire [0:0] cby_1__1__104_left_grid_pin_18_;
  wire [0:0] cby_1__1__104_left_grid_pin_19_;
  wire [0:0] cby_1__1__104_left_grid_pin_20_;
  wire [0:0] cby_1__1__104_left_grid_pin_21_;
  wire [0:0] cby_1__1__104_left_grid_pin_22_;
  wire [0:0] cby_1__1__104_left_grid_pin_23_;
  wire [0:0] cby_1__1__104_left_grid_pin_24_;
  wire [0:0] cby_1__1__104_left_grid_pin_25_;
  wire [0:0] cby_1__1__104_left_grid_pin_26_;
  wire [0:0] cby_1__1__104_left_grid_pin_27_;
  wire [0:0] cby_1__1__104_left_grid_pin_28_;
  wire [0:0] cby_1__1__104_left_grid_pin_29_;
  wire [0:0] cby_1__1__104_left_grid_pin_30_;
  wire [0:0] cby_1__1__104_left_grid_pin_31_;
  wire [0:0] cby_1__1__105_ccff_tail;
  wire [0:29] cby_1__1__105_chany_bottom_out;
  wire [0:29] cby_1__1__105_chany_top_out;
  wire [0:0] cby_1__1__105_left_grid_pin_16_;
  wire [0:0] cby_1__1__105_left_grid_pin_17_;
  wire [0:0] cby_1__1__105_left_grid_pin_18_;
  wire [0:0] cby_1__1__105_left_grid_pin_19_;
  wire [0:0] cby_1__1__105_left_grid_pin_20_;
  wire [0:0] cby_1__1__105_left_grid_pin_21_;
  wire [0:0] cby_1__1__105_left_grid_pin_22_;
  wire [0:0] cby_1__1__105_left_grid_pin_23_;
  wire [0:0] cby_1__1__105_left_grid_pin_24_;
  wire [0:0] cby_1__1__105_left_grid_pin_25_;
  wire [0:0] cby_1__1__105_left_grid_pin_26_;
  wire [0:0] cby_1__1__105_left_grid_pin_27_;
  wire [0:0] cby_1__1__105_left_grid_pin_28_;
  wire [0:0] cby_1__1__105_left_grid_pin_29_;
  wire [0:0] cby_1__1__105_left_grid_pin_30_;
  wire [0:0] cby_1__1__105_left_grid_pin_31_;
  wire [0:0] cby_1__1__106_ccff_tail;
  wire [0:29] cby_1__1__106_chany_bottom_out;
  wire [0:29] cby_1__1__106_chany_top_out;
  wire [0:0] cby_1__1__106_left_grid_pin_16_;
  wire [0:0] cby_1__1__106_left_grid_pin_17_;
  wire [0:0] cby_1__1__106_left_grid_pin_18_;
  wire [0:0] cby_1__1__106_left_grid_pin_19_;
  wire [0:0] cby_1__1__106_left_grid_pin_20_;
  wire [0:0] cby_1__1__106_left_grid_pin_21_;
  wire [0:0] cby_1__1__106_left_grid_pin_22_;
  wire [0:0] cby_1__1__106_left_grid_pin_23_;
  wire [0:0] cby_1__1__106_left_grid_pin_24_;
  wire [0:0] cby_1__1__106_left_grid_pin_25_;
  wire [0:0] cby_1__1__106_left_grid_pin_26_;
  wire [0:0] cby_1__1__106_left_grid_pin_27_;
  wire [0:0] cby_1__1__106_left_grid_pin_28_;
  wire [0:0] cby_1__1__106_left_grid_pin_29_;
  wire [0:0] cby_1__1__106_left_grid_pin_30_;
  wire [0:0] cby_1__1__106_left_grid_pin_31_;
  wire [0:0] cby_1__1__107_ccff_tail;
  wire [0:29] cby_1__1__107_chany_bottom_out;
  wire [0:29] cby_1__1__107_chany_top_out;
  wire [0:0] cby_1__1__107_left_grid_pin_16_;
  wire [0:0] cby_1__1__107_left_grid_pin_17_;
  wire [0:0] cby_1__1__107_left_grid_pin_18_;
  wire [0:0] cby_1__1__107_left_grid_pin_19_;
  wire [0:0] cby_1__1__107_left_grid_pin_20_;
  wire [0:0] cby_1__1__107_left_grid_pin_21_;
  wire [0:0] cby_1__1__107_left_grid_pin_22_;
  wire [0:0] cby_1__1__107_left_grid_pin_23_;
  wire [0:0] cby_1__1__107_left_grid_pin_24_;
  wire [0:0] cby_1__1__107_left_grid_pin_25_;
  wire [0:0] cby_1__1__107_left_grid_pin_26_;
  wire [0:0] cby_1__1__107_left_grid_pin_27_;
  wire [0:0] cby_1__1__107_left_grid_pin_28_;
  wire [0:0] cby_1__1__107_left_grid_pin_29_;
  wire [0:0] cby_1__1__107_left_grid_pin_30_;
  wire [0:0] cby_1__1__107_left_grid_pin_31_;
  wire [0:0] cby_1__1__108_ccff_tail;
  wire [0:29] cby_1__1__108_chany_bottom_out;
  wire [0:29] cby_1__1__108_chany_top_out;
  wire [0:0] cby_1__1__108_left_grid_pin_16_;
  wire [0:0] cby_1__1__108_left_grid_pin_17_;
  wire [0:0] cby_1__1__108_left_grid_pin_18_;
  wire [0:0] cby_1__1__108_left_grid_pin_19_;
  wire [0:0] cby_1__1__108_left_grid_pin_20_;
  wire [0:0] cby_1__1__108_left_grid_pin_21_;
  wire [0:0] cby_1__1__108_left_grid_pin_22_;
  wire [0:0] cby_1__1__108_left_grid_pin_23_;
  wire [0:0] cby_1__1__108_left_grid_pin_24_;
  wire [0:0] cby_1__1__108_left_grid_pin_25_;
  wire [0:0] cby_1__1__108_left_grid_pin_26_;
  wire [0:0] cby_1__1__108_left_grid_pin_27_;
  wire [0:0] cby_1__1__108_left_grid_pin_28_;
  wire [0:0] cby_1__1__108_left_grid_pin_29_;
  wire [0:0] cby_1__1__108_left_grid_pin_30_;
  wire [0:0] cby_1__1__108_left_grid_pin_31_;
  wire [0:0] cby_1__1__109_ccff_tail;
  wire [0:29] cby_1__1__109_chany_bottom_out;
  wire [0:29] cby_1__1__109_chany_top_out;
  wire [0:0] cby_1__1__109_left_grid_pin_16_;
  wire [0:0] cby_1__1__109_left_grid_pin_17_;
  wire [0:0] cby_1__1__109_left_grid_pin_18_;
  wire [0:0] cby_1__1__109_left_grid_pin_19_;
  wire [0:0] cby_1__1__109_left_grid_pin_20_;
  wire [0:0] cby_1__1__109_left_grid_pin_21_;
  wire [0:0] cby_1__1__109_left_grid_pin_22_;
  wire [0:0] cby_1__1__109_left_grid_pin_23_;
  wire [0:0] cby_1__1__109_left_grid_pin_24_;
  wire [0:0] cby_1__1__109_left_grid_pin_25_;
  wire [0:0] cby_1__1__109_left_grid_pin_26_;
  wire [0:0] cby_1__1__109_left_grid_pin_27_;
  wire [0:0] cby_1__1__109_left_grid_pin_28_;
  wire [0:0] cby_1__1__109_left_grid_pin_29_;
  wire [0:0] cby_1__1__109_left_grid_pin_30_;
  wire [0:0] cby_1__1__109_left_grid_pin_31_;
  wire [0:0] cby_1__1__10_ccff_tail;
  wire [0:29] cby_1__1__10_chany_bottom_out;
  wire [0:29] cby_1__1__10_chany_top_out;
  wire [0:0] cby_1__1__10_left_grid_pin_16_;
  wire [0:0] cby_1__1__10_left_grid_pin_17_;
  wire [0:0] cby_1__1__10_left_grid_pin_18_;
  wire [0:0] cby_1__1__10_left_grid_pin_19_;
  wire [0:0] cby_1__1__10_left_grid_pin_20_;
  wire [0:0] cby_1__1__10_left_grid_pin_21_;
  wire [0:0] cby_1__1__10_left_grid_pin_22_;
  wire [0:0] cby_1__1__10_left_grid_pin_23_;
  wire [0:0] cby_1__1__10_left_grid_pin_24_;
  wire [0:0] cby_1__1__10_left_grid_pin_25_;
  wire [0:0] cby_1__1__10_left_grid_pin_26_;
  wire [0:0] cby_1__1__10_left_grid_pin_27_;
  wire [0:0] cby_1__1__10_left_grid_pin_28_;
  wire [0:0] cby_1__1__10_left_grid_pin_29_;
  wire [0:0] cby_1__1__10_left_grid_pin_30_;
  wire [0:0] cby_1__1__10_left_grid_pin_31_;
  wire [0:0] cby_1__1__110_ccff_tail;
  wire [0:29] cby_1__1__110_chany_bottom_out;
  wire [0:29] cby_1__1__110_chany_top_out;
  wire [0:0] cby_1__1__110_left_grid_pin_16_;
  wire [0:0] cby_1__1__110_left_grid_pin_17_;
  wire [0:0] cby_1__1__110_left_grid_pin_18_;
  wire [0:0] cby_1__1__110_left_grid_pin_19_;
  wire [0:0] cby_1__1__110_left_grid_pin_20_;
  wire [0:0] cby_1__1__110_left_grid_pin_21_;
  wire [0:0] cby_1__1__110_left_grid_pin_22_;
  wire [0:0] cby_1__1__110_left_grid_pin_23_;
  wire [0:0] cby_1__1__110_left_grid_pin_24_;
  wire [0:0] cby_1__1__110_left_grid_pin_25_;
  wire [0:0] cby_1__1__110_left_grid_pin_26_;
  wire [0:0] cby_1__1__110_left_grid_pin_27_;
  wire [0:0] cby_1__1__110_left_grid_pin_28_;
  wire [0:0] cby_1__1__110_left_grid_pin_29_;
  wire [0:0] cby_1__1__110_left_grid_pin_30_;
  wire [0:0] cby_1__1__110_left_grid_pin_31_;
  wire [0:0] cby_1__1__111_ccff_tail;
  wire [0:29] cby_1__1__111_chany_bottom_out;
  wire [0:29] cby_1__1__111_chany_top_out;
  wire [0:0] cby_1__1__111_left_grid_pin_16_;
  wire [0:0] cby_1__1__111_left_grid_pin_17_;
  wire [0:0] cby_1__1__111_left_grid_pin_18_;
  wire [0:0] cby_1__1__111_left_grid_pin_19_;
  wire [0:0] cby_1__1__111_left_grid_pin_20_;
  wire [0:0] cby_1__1__111_left_grid_pin_21_;
  wire [0:0] cby_1__1__111_left_grid_pin_22_;
  wire [0:0] cby_1__1__111_left_grid_pin_23_;
  wire [0:0] cby_1__1__111_left_grid_pin_24_;
  wire [0:0] cby_1__1__111_left_grid_pin_25_;
  wire [0:0] cby_1__1__111_left_grid_pin_26_;
  wire [0:0] cby_1__1__111_left_grid_pin_27_;
  wire [0:0] cby_1__1__111_left_grid_pin_28_;
  wire [0:0] cby_1__1__111_left_grid_pin_29_;
  wire [0:0] cby_1__1__111_left_grid_pin_30_;
  wire [0:0] cby_1__1__111_left_grid_pin_31_;
  wire [0:0] cby_1__1__112_ccff_tail;
  wire [0:29] cby_1__1__112_chany_bottom_out;
  wire [0:29] cby_1__1__112_chany_top_out;
  wire [0:0] cby_1__1__112_left_grid_pin_16_;
  wire [0:0] cby_1__1__112_left_grid_pin_17_;
  wire [0:0] cby_1__1__112_left_grid_pin_18_;
  wire [0:0] cby_1__1__112_left_grid_pin_19_;
  wire [0:0] cby_1__1__112_left_grid_pin_20_;
  wire [0:0] cby_1__1__112_left_grid_pin_21_;
  wire [0:0] cby_1__1__112_left_grid_pin_22_;
  wire [0:0] cby_1__1__112_left_grid_pin_23_;
  wire [0:0] cby_1__1__112_left_grid_pin_24_;
  wire [0:0] cby_1__1__112_left_grid_pin_25_;
  wire [0:0] cby_1__1__112_left_grid_pin_26_;
  wire [0:0] cby_1__1__112_left_grid_pin_27_;
  wire [0:0] cby_1__1__112_left_grid_pin_28_;
  wire [0:0] cby_1__1__112_left_grid_pin_29_;
  wire [0:0] cby_1__1__112_left_grid_pin_30_;
  wire [0:0] cby_1__1__112_left_grid_pin_31_;
  wire [0:0] cby_1__1__113_ccff_tail;
  wire [0:29] cby_1__1__113_chany_bottom_out;
  wire [0:29] cby_1__1__113_chany_top_out;
  wire [0:0] cby_1__1__113_left_grid_pin_16_;
  wire [0:0] cby_1__1__113_left_grid_pin_17_;
  wire [0:0] cby_1__1__113_left_grid_pin_18_;
  wire [0:0] cby_1__1__113_left_grid_pin_19_;
  wire [0:0] cby_1__1__113_left_grid_pin_20_;
  wire [0:0] cby_1__1__113_left_grid_pin_21_;
  wire [0:0] cby_1__1__113_left_grid_pin_22_;
  wire [0:0] cby_1__1__113_left_grid_pin_23_;
  wire [0:0] cby_1__1__113_left_grid_pin_24_;
  wire [0:0] cby_1__1__113_left_grid_pin_25_;
  wire [0:0] cby_1__1__113_left_grid_pin_26_;
  wire [0:0] cby_1__1__113_left_grid_pin_27_;
  wire [0:0] cby_1__1__113_left_grid_pin_28_;
  wire [0:0] cby_1__1__113_left_grid_pin_29_;
  wire [0:0] cby_1__1__113_left_grid_pin_30_;
  wire [0:0] cby_1__1__113_left_grid_pin_31_;
  wire [0:0] cby_1__1__114_ccff_tail;
  wire [0:29] cby_1__1__114_chany_bottom_out;
  wire [0:29] cby_1__1__114_chany_top_out;
  wire [0:0] cby_1__1__114_left_grid_pin_16_;
  wire [0:0] cby_1__1__114_left_grid_pin_17_;
  wire [0:0] cby_1__1__114_left_grid_pin_18_;
  wire [0:0] cby_1__1__114_left_grid_pin_19_;
  wire [0:0] cby_1__1__114_left_grid_pin_20_;
  wire [0:0] cby_1__1__114_left_grid_pin_21_;
  wire [0:0] cby_1__1__114_left_grid_pin_22_;
  wire [0:0] cby_1__1__114_left_grid_pin_23_;
  wire [0:0] cby_1__1__114_left_grid_pin_24_;
  wire [0:0] cby_1__1__114_left_grid_pin_25_;
  wire [0:0] cby_1__1__114_left_grid_pin_26_;
  wire [0:0] cby_1__1__114_left_grid_pin_27_;
  wire [0:0] cby_1__1__114_left_grid_pin_28_;
  wire [0:0] cby_1__1__114_left_grid_pin_29_;
  wire [0:0] cby_1__1__114_left_grid_pin_30_;
  wire [0:0] cby_1__1__114_left_grid_pin_31_;
  wire [0:0] cby_1__1__115_ccff_tail;
  wire [0:29] cby_1__1__115_chany_bottom_out;
  wire [0:29] cby_1__1__115_chany_top_out;
  wire [0:0] cby_1__1__115_left_grid_pin_16_;
  wire [0:0] cby_1__1__115_left_grid_pin_17_;
  wire [0:0] cby_1__1__115_left_grid_pin_18_;
  wire [0:0] cby_1__1__115_left_grid_pin_19_;
  wire [0:0] cby_1__1__115_left_grid_pin_20_;
  wire [0:0] cby_1__1__115_left_grid_pin_21_;
  wire [0:0] cby_1__1__115_left_grid_pin_22_;
  wire [0:0] cby_1__1__115_left_grid_pin_23_;
  wire [0:0] cby_1__1__115_left_grid_pin_24_;
  wire [0:0] cby_1__1__115_left_grid_pin_25_;
  wire [0:0] cby_1__1__115_left_grid_pin_26_;
  wire [0:0] cby_1__1__115_left_grid_pin_27_;
  wire [0:0] cby_1__1__115_left_grid_pin_28_;
  wire [0:0] cby_1__1__115_left_grid_pin_29_;
  wire [0:0] cby_1__1__115_left_grid_pin_30_;
  wire [0:0] cby_1__1__115_left_grid_pin_31_;
  wire [0:0] cby_1__1__116_ccff_tail;
  wire [0:29] cby_1__1__116_chany_bottom_out;
  wire [0:29] cby_1__1__116_chany_top_out;
  wire [0:0] cby_1__1__116_left_grid_pin_16_;
  wire [0:0] cby_1__1__116_left_grid_pin_17_;
  wire [0:0] cby_1__1__116_left_grid_pin_18_;
  wire [0:0] cby_1__1__116_left_grid_pin_19_;
  wire [0:0] cby_1__1__116_left_grid_pin_20_;
  wire [0:0] cby_1__1__116_left_grid_pin_21_;
  wire [0:0] cby_1__1__116_left_grid_pin_22_;
  wire [0:0] cby_1__1__116_left_grid_pin_23_;
  wire [0:0] cby_1__1__116_left_grid_pin_24_;
  wire [0:0] cby_1__1__116_left_grid_pin_25_;
  wire [0:0] cby_1__1__116_left_grid_pin_26_;
  wire [0:0] cby_1__1__116_left_grid_pin_27_;
  wire [0:0] cby_1__1__116_left_grid_pin_28_;
  wire [0:0] cby_1__1__116_left_grid_pin_29_;
  wire [0:0] cby_1__1__116_left_grid_pin_30_;
  wire [0:0] cby_1__1__116_left_grid_pin_31_;
  wire [0:0] cby_1__1__117_ccff_tail;
  wire [0:29] cby_1__1__117_chany_bottom_out;
  wire [0:29] cby_1__1__117_chany_top_out;
  wire [0:0] cby_1__1__117_left_grid_pin_16_;
  wire [0:0] cby_1__1__117_left_grid_pin_17_;
  wire [0:0] cby_1__1__117_left_grid_pin_18_;
  wire [0:0] cby_1__1__117_left_grid_pin_19_;
  wire [0:0] cby_1__1__117_left_grid_pin_20_;
  wire [0:0] cby_1__1__117_left_grid_pin_21_;
  wire [0:0] cby_1__1__117_left_grid_pin_22_;
  wire [0:0] cby_1__1__117_left_grid_pin_23_;
  wire [0:0] cby_1__1__117_left_grid_pin_24_;
  wire [0:0] cby_1__1__117_left_grid_pin_25_;
  wire [0:0] cby_1__1__117_left_grid_pin_26_;
  wire [0:0] cby_1__1__117_left_grid_pin_27_;
  wire [0:0] cby_1__1__117_left_grid_pin_28_;
  wire [0:0] cby_1__1__117_left_grid_pin_29_;
  wire [0:0] cby_1__1__117_left_grid_pin_30_;
  wire [0:0] cby_1__1__117_left_grid_pin_31_;
  wire [0:0] cby_1__1__118_ccff_tail;
  wire [0:29] cby_1__1__118_chany_bottom_out;
  wire [0:29] cby_1__1__118_chany_top_out;
  wire [0:0] cby_1__1__118_left_grid_pin_16_;
  wire [0:0] cby_1__1__118_left_grid_pin_17_;
  wire [0:0] cby_1__1__118_left_grid_pin_18_;
  wire [0:0] cby_1__1__118_left_grid_pin_19_;
  wire [0:0] cby_1__1__118_left_grid_pin_20_;
  wire [0:0] cby_1__1__118_left_grid_pin_21_;
  wire [0:0] cby_1__1__118_left_grid_pin_22_;
  wire [0:0] cby_1__1__118_left_grid_pin_23_;
  wire [0:0] cby_1__1__118_left_grid_pin_24_;
  wire [0:0] cby_1__1__118_left_grid_pin_25_;
  wire [0:0] cby_1__1__118_left_grid_pin_26_;
  wire [0:0] cby_1__1__118_left_grid_pin_27_;
  wire [0:0] cby_1__1__118_left_grid_pin_28_;
  wire [0:0] cby_1__1__118_left_grid_pin_29_;
  wire [0:0] cby_1__1__118_left_grid_pin_30_;
  wire [0:0] cby_1__1__118_left_grid_pin_31_;
  wire [0:0] cby_1__1__119_ccff_tail;
  wire [0:29] cby_1__1__119_chany_bottom_out;
  wire [0:29] cby_1__1__119_chany_top_out;
  wire [0:0] cby_1__1__119_left_grid_pin_16_;
  wire [0:0] cby_1__1__119_left_grid_pin_17_;
  wire [0:0] cby_1__1__119_left_grid_pin_18_;
  wire [0:0] cby_1__1__119_left_grid_pin_19_;
  wire [0:0] cby_1__1__119_left_grid_pin_20_;
  wire [0:0] cby_1__1__119_left_grid_pin_21_;
  wire [0:0] cby_1__1__119_left_grid_pin_22_;
  wire [0:0] cby_1__1__119_left_grid_pin_23_;
  wire [0:0] cby_1__1__119_left_grid_pin_24_;
  wire [0:0] cby_1__1__119_left_grid_pin_25_;
  wire [0:0] cby_1__1__119_left_grid_pin_26_;
  wire [0:0] cby_1__1__119_left_grid_pin_27_;
  wire [0:0] cby_1__1__119_left_grid_pin_28_;
  wire [0:0] cby_1__1__119_left_grid_pin_29_;
  wire [0:0] cby_1__1__119_left_grid_pin_30_;
  wire [0:0] cby_1__1__119_left_grid_pin_31_;
  wire [0:0] cby_1__1__11_ccff_tail;
  wire [0:29] cby_1__1__11_chany_bottom_out;
  wire [0:29] cby_1__1__11_chany_top_out;
  wire [0:0] cby_1__1__11_left_grid_pin_16_;
  wire [0:0] cby_1__1__11_left_grid_pin_17_;
  wire [0:0] cby_1__1__11_left_grid_pin_18_;
  wire [0:0] cby_1__1__11_left_grid_pin_19_;
  wire [0:0] cby_1__1__11_left_grid_pin_20_;
  wire [0:0] cby_1__1__11_left_grid_pin_21_;
  wire [0:0] cby_1__1__11_left_grid_pin_22_;
  wire [0:0] cby_1__1__11_left_grid_pin_23_;
  wire [0:0] cby_1__1__11_left_grid_pin_24_;
  wire [0:0] cby_1__1__11_left_grid_pin_25_;
  wire [0:0] cby_1__1__11_left_grid_pin_26_;
  wire [0:0] cby_1__1__11_left_grid_pin_27_;
  wire [0:0] cby_1__1__11_left_grid_pin_28_;
  wire [0:0] cby_1__1__11_left_grid_pin_29_;
  wire [0:0] cby_1__1__11_left_grid_pin_30_;
  wire [0:0] cby_1__1__11_left_grid_pin_31_;
  wire [0:0] cby_1__1__120_ccff_tail;
  wire [0:29] cby_1__1__120_chany_bottom_out;
  wire [0:29] cby_1__1__120_chany_top_out;
  wire [0:0] cby_1__1__120_left_grid_pin_16_;
  wire [0:0] cby_1__1__120_left_grid_pin_17_;
  wire [0:0] cby_1__1__120_left_grid_pin_18_;
  wire [0:0] cby_1__1__120_left_grid_pin_19_;
  wire [0:0] cby_1__1__120_left_grid_pin_20_;
  wire [0:0] cby_1__1__120_left_grid_pin_21_;
  wire [0:0] cby_1__1__120_left_grid_pin_22_;
  wire [0:0] cby_1__1__120_left_grid_pin_23_;
  wire [0:0] cby_1__1__120_left_grid_pin_24_;
  wire [0:0] cby_1__1__120_left_grid_pin_25_;
  wire [0:0] cby_1__1__120_left_grid_pin_26_;
  wire [0:0] cby_1__1__120_left_grid_pin_27_;
  wire [0:0] cby_1__1__120_left_grid_pin_28_;
  wire [0:0] cby_1__1__120_left_grid_pin_29_;
  wire [0:0] cby_1__1__120_left_grid_pin_30_;
  wire [0:0] cby_1__1__120_left_grid_pin_31_;
  wire [0:0] cby_1__1__121_ccff_tail;
  wire [0:29] cby_1__1__121_chany_bottom_out;
  wire [0:29] cby_1__1__121_chany_top_out;
  wire [0:0] cby_1__1__121_left_grid_pin_16_;
  wire [0:0] cby_1__1__121_left_grid_pin_17_;
  wire [0:0] cby_1__1__121_left_grid_pin_18_;
  wire [0:0] cby_1__1__121_left_grid_pin_19_;
  wire [0:0] cby_1__1__121_left_grid_pin_20_;
  wire [0:0] cby_1__1__121_left_grid_pin_21_;
  wire [0:0] cby_1__1__121_left_grid_pin_22_;
  wire [0:0] cby_1__1__121_left_grid_pin_23_;
  wire [0:0] cby_1__1__121_left_grid_pin_24_;
  wire [0:0] cby_1__1__121_left_grid_pin_25_;
  wire [0:0] cby_1__1__121_left_grid_pin_26_;
  wire [0:0] cby_1__1__121_left_grid_pin_27_;
  wire [0:0] cby_1__1__121_left_grid_pin_28_;
  wire [0:0] cby_1__1__121_left_grid_pin_29_;
  wire [0:0] cby_1__1__121_left_grid_pin_30_;
  wire [0:0] cby_1__1__121_left_grid_pin_31_;
  wire [0:0] cby_1__1__122_ccff_tail;
  wire [0:29] cby_1__1__122_chany_bottom_out;
  wire [0:29] cby_1__1__122_chany_top_out;
  wire [0:0] cby_1__1__122_left_grid_pin_16_;
  wire [0:0] cby_1__1__122_left_grid_pin_17_;
  wire [0:0] cby_1__1__122_left_grid_pin_18_;
  wire [0:0] cby_1__1__122_left_grid_pin_19_;
  wire [0:0] cby_1__1__122_left_grid_pin_20_;
  wire [0:0] cby_1__1__122_left_grid_pin_21_;
  wire [0:0] cby_1__1__122_left_grid_pin_22_;
  wire [0:0] cby_1__1__122_left_grid_pin_23_;
  wire [0:0] cby_1__1__122_left_grid_pin_24_;
  wire [0:0] cby_1__1__122_left_grid_pin_25_;
  wire [0:0] cby_1__1__122_left_grid_pin_26_;
  wire [0:0] cby_1__1__122_left_grid_pin_27_;
  wire [0:0] cby_1__1__122_left_grid_pin_28_;
  wire [0:0] cby_1__1__122_left_grid_pin_29_;
  wire [0:0] cby_1__1__122_left_grid_pin_30_;
  wire [0:0] cby_1__1__122_left_grid_pin_31_;
  wire [0:0] cby_1__1__123_ccff_tail;
  wire [0:29] cby_1__1__123_chany_bottom_out;
  wire [0:29] cby_1__1__123_chany_top_out;
  wire [0:0] cby_1__1__123_left_grid_pin_16_;
  wire [0:0] cby_1__1__123_left_grid_pin_17_;
  wire [0:0] cby_1__1__123_left_grid_pin_18_;
  wire [0:0] cby_1__1__123_left_grid_pin_19_;
  wire [0:0] cby_1__1__123_left_grid_pin_20_;
  wire [0:0] cby_1__1__123_left_grid_pin_21_;
  wire [0:0] cby_1__1__123_left_grid_pin_22_;
  wire [0:0] cby_1__1__123_left_grid_pin_23_;
  wire [0:0] cby_1__1__123_left_grid_pin_24_;
  wire [0:0] cby_1__1__123_left_grid_pin_25_;
  wire [0:0] cby_1__1__123_left_grid_pin_26_;
  wire [0:0] cby_1__1__123_left_grid_pin_27_;
  wire [0:0] cby_1__1__123_left_grid_pin_28_;
  wire [0:0] cby_1__1__123_left_grid_pin_29_;
  wire [0:0] cby_1__1__123_left_grid_pin_30_;
  wire [0:0] cby_1__1__123_left_grid_pin_31_;
  wire [0:0] cby_1__1__124_ccff_tail;
  wire [0:29] cby_1__1__124_chany_bottom_out;
  wire [0:29] cby_1__1__124_chany_top_out;
  wire [0:0] cby_1__1__124_left_grid_pin_16_;
  wire [0:0] cby_1__1__124_left_grid_pin_17_;
  wire [0:0] cby_1__1__124_left_grid_pin_18_;
  wire [0:0] cby_1__1__124_left_grid_pin_19_;
  wire [0:0] cby_1__1__124_left_grid_pin_20_;
  wire [0:0] cby_1__1__124_left_grid_pin_21_;
  wire [0:0] cby_1__1__124_left_grid_pin_22_;
  wire [0:0] cby_1__1__124_left_grid_pin_23_;
  wire [0:0] cby_1__1__124_left_grid_pin_24_;
  wire [0:0] cby_1__1__124_left_grid_pin_25_;
  wire [0:0] cby_1__1__124_left_grid_pin_26_;
  wire [0:0] cby_1__1__124_left_grid_pin_27_;
  wire [0:0] cby_1__1__124_left_grid_pin_28_;
  wire [0:0] cby_1__1__124_left_grid_pin_29_;
  wire [0:0] cby_1__1__124_left_grid_pin_30_;
  wire [0:0] cby_1__1__124_left_grid_pin_31_;
  wire [0:0] cby_1__1__125_ccff_tail;
  wire [0:29] cby_1__1__125_chany_bottom_out;
  wire [0:29] cby_1__1__125_chany_top_out;
  wire [0:0] cby_1__1__125_left_grid_pin_16_;
  wire [0:0] cby_1__1__125_left_grid_pin_17_;
  wire [0:0] cby_1__1__125_left_grid_pin_18_;
  wire [0:0] cby_1__1__125_left_grid_pin_19_;
  wire [0:0] cby_1__1__125_left_grid_pin_20_;
  wire [0:0] cby_1__1__125_left_grid_pin_21_;
  wire [0:0] cby_1__1__125_left_grid_pin_22_;
  wire [0:0] cby_1__1__125_left_grid_pin_23_;
  wire [0:0] cby_1__1__125_left_grid_pin_24_;
  wire [0:0] cby_1__1__125_left_grid_pin_25_;
  wire [0:0] cby_1__1__125_left_grid_pin_26_;
  wire [0:0] cby_1__1__125_left_grid_pin_27_;
  wire [0:0] cby_1__1__125_left_grid_pin_28_;
  wire [0:0] cby_1__1__125_left_grid_pin_29_;
  wire [0:0] cby_1__1__125_left_grid_pin_30_;
  wire [0:0] cby_1__1__125_left_grid_pin_31_;
  wire [0:0] cby_1__1__126_ccff_tail;
  wire [0:29] cby_1__1__126_chany_bottom_out;
  wire [0:29] cby_1__1__126_chany_top_out;
  wire [0:0] cby_1__1__126_left_grid_pin_16_;
  wire [0:0] cby_1__1__126_left_grid_pin_17_;
  wire [0:0] cby_1__1__126_left_grid_pin_18_;
  wire [0:0] cby_1__1__126_left_grid_pin_19_;
  wire [0:0] cby_1__1__126_left_grid_pin_20_;
  wire [0:0] cby_1__1__126_left_grid_pin_21_;
  wire [0:0] cby_1__1__126_left_grid_pin_22_;
  wire [0:0] cby_1__1__126_left_grid_pin_23_;
  wire [0:0] cby_1__1__126_left_grid_pin_24_;
  wire [0:0] cby_1__1__126_left_grid_pin_25_;
  wire [0:0] cby_1__1__126_left_grid_pin_26_;
  wire [0:0] cby_1__1__126_left_grid_pin_27_;
  wire [0:0] cby_1__1__126_left_grid_pin_28_;
  wire [0:0] cby_1__1__126_left_grid_pin_29_;
  wire [0:0] cby_1__1__126_left_grid_pin_30_;
  wire [0:0] cby_1__1__126_left_grid_pin_31_;
  wire [0:0] cby_1__1__127_ccff_tail;
  wire [0:29] cby_1__1__127_chany_bottom_out;
  wire [0:29] cby_1__1__127_chany_top_out;
  wire [0:0] cby_1__1__127_left_grid_pin_16_;
  wire [0:0] cby_1__1__127_left_grid_pin_17_;
  wire [0:0] cby_1__1__127_left_grid_pin_18_;
  wire [0:0] cby_1__1__127_left_grid_pin_19_;
  wire [0:0] cby_1__1__127_left_grid_pin_20_;
  wire [0:0] cby_1__1__127_left_grid_pin_21_;
  wire [0:0] cby_1__1__127_left_grid_pin_22_;
  wire [0:0] cby_1__1__127_left_grid_pin_23_;
  wire [0:0] cby_1__1__127_left_grid_pin_24_;
  wire [0:0] cby_1__1__127_left_grid_pin_25_;
  wire [0:0] cby_1__1__127_left_grid_pin_26_;
  wire [0:0] cby_1__1__127_left_grid_pin_27_;
  wire [0:0] cby_1__1__127_left_grid_pin_28_;
  wire [0:0] cby_1__1__127_left_grid_pin_29_;
  wire [0:0] cby_1__1__127_left_grid_pin_30_;
  wire [0:0] cby_1__1__127_left_grid_pin_31_;
  wire [0:0] cby_1__1__128_ccff_tail;
  wire [0:29] cby_1__1__128_chany_bottom_out;
  wire [0:29] cby_1__1__128_chany_top_out;
  wire [0:0] cby_1__1__128_left_grid_pin_16_;
  wire [0:0] cby_1__1__128_left_grid_pin_17_;
  wire [0:0] cby_1__1__128_left_grid_pin_18_;
  wire [0:0] cby_1__1__128_left_grid_pin_19_;
  wire [0:0] cby_1__1__128_left_grid_pin_20_;
  wire [0:0] cby_1__1__128_left_grid_pin_21_;
  wire [0:0] cby_1__1__128_left_grid_pin_22_;
  wire [0:0] cby_1__1__128_left_grid_pin_23_;
  wire [0:0] cby_1__1__128_left_grid_pin_24_;
  wire [0:0] cby_1__1__128_left_grid_pin_25_;
  wire [0:0] cby_1__1__128_left_grid_pin_26_;
  wire [0:0] cby_1__1__128_left_grid_pin_27_;
  wire [0:0] cby_1__1__128_left_grid_pin_28_;
  wire [0:0] cby_1__1__128_left_grid_pin_29_;
  wire [0:0] cby_1__1__128_left_grid_pin_30_;
  wire [0:0] cby_1__1__128_left_grid_pin_31_;
  wire [0:0] cby_1__1__129_ccff_tail;
  wire [0:29] cby_1__1__129_chany_bottom_out;
  wire [0:29] cby_1__1__129_chany_top_out;
  wire [0:0] cby_1__1__129_left_grid_pin_16_;
  wire [0:0] cby_1__1__129_left_grid_pin_17_;
  wire [0:0] cby_1__1__129_left_grid_pin_18_;
  wire [0:0] cby_1__1__129_left_grid_pin_19_;
  wire [0:0] cby_1__1__129_left_grid_pin_20_;
  wire [0:0] cby_1__1__129_left_grid_pin_21_;
  wire [0:0] cby_1__1__129_left_grid_pin_22_;
  wire [0:0] cby_1__1__129_left_grid_pin_23_;
  wire [0:0] cby_1__1__129_left_grid_pin_24_;
  wire [0:0] cby_1__1__129_left_grid_pin_25_;
  wire [0:0] cby_1__1__129_left_grid_pin_26_;
  wire [0:0] cby_1__1__129_left_grid_pin_27_;
  wire [0:0] cby_1__1__129_left_grid_pin_28_;
  wire [0:0] cby_1__1__129_left_grid_pin_29_;
  wire [0:0] cby_1__1__129_left_grid_pin_30_;
  wire [0:0] cby_1__1__129_left_grid_pin_31_;
  wire [0:0] cby_1__1__12_ccff_tail;
  wire [0:29] cby_1__1__12_chany_bottom_out;
  wire [0:29] cby_1__1__12_chany_top_out;
  wire [0:0] cby_1__1__12_left_grid_pin_16_;
  wire [0:0] cby_1__1__12_left_grid_pin_17_;
  wire [0:0] cby_1__1__12_left_grid_pin_18_;
  wire [0:0] cby_1__1__12_left_grid_pin_19_;
  wire [0:0] cby_1__1__12_left_grid_pin_20_;
  wire [0:0] cby_1__1__12_left_grid_pin_21_;
  wire [0:0] cby_1__1__12_left_grid_pin_22_;
  wire [0:0] cby_1__1__12_left_grid_pin_23_;
  wire [0:0] cby_1__1__12_left_grid_pin_24_;
  wire [0:0] cby_1__1__12_left_grid_pin_25_;
  wire [0:0] cby_1__1__12_left_grid_pin_26_;
  wire [0:0] cby_1__1__12_left_grid_pin_27_;
  wire [0:0] cby_1__1__12_left_grid_pin_28_;
  wire [0:0] cby_1__1__12_left_grid_pin_29_;
  wire [0:0] cby_1__1__12_left_grid_pin_30_;
  wire [0:0] cby_1__1__12_left_grid_pin_31_;
  wire [0:0] cby_1__1__130_ccff_tail;
  wire [0:29] cby_1__1__130_chany_bottom_out;
  wire [0:29] cby_1__1__130_chany_top_out;
  wire [0:0] cby_1__1__130_left_grid_pin_16_;
  wire [0:0] cby_1__1__130_left_grid_pin_17_;
  wire [0:0] cby_1__1__130_left_grid_pin_18_;
  wire [0:0] cby_1__1__130_left_grid_pin_19_;
  wire [0:0] cby_1__1__130_left_grid_pin_20_;
  wire [0:0] cby_1__1__130_left_grid_pin_21_;
  wire [0:0] cby_1__1__130_left_grid_pin_22_;
  wire [0:0] cby_1__1__130_left_grid_pin_23_;
  wire [0:0] cby_1__1__130_left_grid_pin_24_;
  wire [0:0] cby_1__1__130_left_grid_pin_25_;
  wire [0:0] cby_1__1__130_left_grid_pin_26_;
  wire [0:0] cby_1__1__130_left_grid_pin_27_;
  wire [0:0] cby_1__1__130_left_grid_pin_28_;
  wire [0:0] cby_1__1__130_left_grid_pin_29_;
  wire [0:0] cby_1__1__130_left_grid_pin_30_;
  wire [0:0] cby_1__1__130_left_grid_pin_31_;
  wire [0:0] cby_1__1__131_ccff_tail;
  wire [0:29] cby_1__1__131_chany_bottom_out;
  wire [0:29] cby_1__1__131_chany_top_out;
  wire [0:0] cby_1__1__131_left_grid_pin_16_;
  wire [0:0] cby_1__1__131_left_grid_pin_17_;
  wire [0:0] cby_1__1__131_left_grid_pin_18_;
  wire [0:0] cby_1__1__131_left_grid_pin_19_;
  wire [0:0] cby_1__1__131_left_grid_pin_20_;
  wire [0:0] cby_1__1__131_left_grid_pin_21_;
  wire [0:0] cby_1__1__131_left_grid_pin_22_;
  wire [0:0] cby_1__1__131_left_grid_pin_23_;
  wire [0:0] cby_1__1__131_left_grid_pin_24_;
  wire [0:0] cby_1__1__131_left_grid_pin_25_;
  wire [0:0] cby_1__1__131_left_grid_pin_26_;
  wire [0:0] cby_1__1__131_left_grid_pin_27_;
  wire [0:0] cby_1__1__131_left_grid_pin_28_;
  wire [0:0] cby_1__1__131_left_grid_pin_29_;
  wire [0:0] cby_1__1__131_left_grid_pin_30_;
  wire [0:0] cby_1__1__131_left_grid_pin_31_;
  wire [0:0] cby_1__1__13_ccff_tail;
  wire [0:29] cby_1__1__13_chany_bottom_out;
  wire [0:29] cby_1__1__13_chany_top_out;
  wire [0:0] cby_1__1__13_left_grid_pin_16_;
  wire [0:0] cby_1__1__13_left_grid_pin_17_;
  wire [0:0] cby_1__1__13_left_grid_pin_18_;
  wire [0:0] cby_1__1__13_left_grid_pin_19_;
  wire [0:0] cby_1__1__13_left_grid_pin_20_;
  wire [0:0] cby_1__1__13_left_grid_pin_21_;
  wire [0:0] cby_1__1__13_left_grid_pin_22_;
  wire [0:0] cby_1__1__13_left_grid_pin_23_;
  wire [0:0] cby_1__1__13_left_grid_pin_24_;
  wire [0:0] cby_1__1__13_left_grid_pin_25_;
  wire [0:0] cby_1__1__13_left_grid_pin_26_;
  wire [0:0] cby_1__1__13_left_grid_pin_27_;
  wire [0:0] cby_1__1__13_left_grid_pin_28_;
  wire [0:0] cby_1__1__13_left_grid_pin_29_;
  wire [0:0] cby_1__1__13_left_grid_pin_30_;
  wire [0:0] cby_1__1__13_left_grid_pin_31_;
  wire [0:0] cby_1__1__14_ccff_tail;
  wire [0:29] cby_1__1__14_chany_bottom_out;
  wire [0:29] cby_1__1__14_chany_top_out;
  wire [0:0] cby_1__1__14_left_grid_pin_16_;
  wire [0:0] cby_1__1__14_left_grid_pin_17_;
  wire [0:0] cby_1__1__14_left_grid_pin_18_;
  wire [0:0] cby_1__1__14_left_grid_pin_19_;
  wire [0:0] cby_1__1__14_left_grid_pin_20_;
  wire [0:0] cby_1__1__14_left_grid_pin_21_;
  wire [0:0] cby_1__1__14_left_grid_pin_22_;
  wire [0:0] cby_1__1__14_left_grid_pin_23_;
  wire [0:0] cby_1__1__14_left_grid_pin_24_;
  wire [0:0] cby_1__1__14_left_grid_pin_25_;
  wire [0:0] cby_1__1__14_left_grid_pin_26_;
  wire [0:0] cby_1__1__14_left_grid_pin_27_;
  wire [0:0] cby_1__1__14_left_grid_pin_28_;
  wire [0:0] cby_1__1__14_left_grid_pin_29_;
  wire [0:0] cby_1__1__14_left_grid_pin_30_;
  wire [0:0] cby_1__1__14_left_grid_pin_31_;
  wire [0:0] cby_1__1__15_ccff_tail;
  wire [0:29] cby_1__1__15_chany_bottom_out;
  wire [0:29] cby_1__1__15_chany_top_out;
  wire [0:0] cby_1__1__15_left_grid_pin_16_;
  wire [0:0] cby_1__1__15_left_grid_pin_17_;
  wire [0:0] cby_1__1__15_left_grid_pin_18_;
  wire [0:0] cby_1__1__15_left_grid_pin_19_;
  wire [0:0] cby_1__1__15_left_grid_pin_20_;
  wire [0:0] cby_1__1__15_left_grid_pin_21_;
  wire [0:0] cby_1__1__15_left_grid_pin_22_;
  wire [0:0] cby_1__1__15_left_grid_pin_23_;
  wire [0:0] cby_1__1__15_left_grid_pin_24_;
  wire [0:0] cby_1__1__15_left_grid_pin_25_;
  wire [0:0] cby_1__1__15_left_grid_pin_26_;
  wire [0:0] cby_1__1__15_left_grid_pin_27_;
  wire [0:0] cby_1__1__15_left_grid_pin_28_;
  wire [0:0] cby_1__1__15_left_grid_pin_29_;
  wire [0:0] cby_1__1__15_left_grid_pin_30_;
  wire [0:0] cby_1__1__15_left_grid_pin_31_;
  wire [0:0] cby_1__1__16_ccff_tail;
  wire [0:29] cby_1__1__16_chany_bottom_out;
  wire [0:29] cby_1__1__16_chany_top_out;
  wire [0:0] cby_1__1__16_left_grid_pin_16_;
  wire [0:0] cby_1__1__16_left_grid_pin_17_;
  wire [0:0] cby_1__1__16_left_grid_pin_18_;
  wire [0:0] cby_1__1__16_left_grid_pin_19_;
  wire [0:0] cby_1__1__16_left_grid_pin_20_;
  wire [0:0] cby_1__1__16_left_grid_pin_21_;
  wire [0:0] cby_1__1__16_left_grid_pin_22_;
  wire [0:0] cby_1__1__16_left_grid_pin_23_;
  wire [0:0] cby_1__1__16_left_grid_pin_24_;
  wire [0:0] cby_1__1__16_left_grid_pin_25_;
  wire [0:0] cby_1__1__16_left_grid_pin_26_;
  wire [0:0] cby_1__1__16_left_grid_pin_27_;
  wire [0:0] cby_1__1__16_left_grid_pin_28_;
  wire [0:0] cby_1__1__16_left_grid_pin_29_;
  wire [0:0] cby_1__1__16_left_grid_pin_30_;
  wire [0:0] cby_1__1__16_left_grid_pin_31_;
  wire [0:0] cby_1__1__17_ccff_tail;
  wire [0:29] cby_1__1__17_chany_bottom_out;
  wire [0:29] cby_1__1__17_chany_top_out;
  wire [0:0] cby_1__1__17_left_grid_pin_16_;
  wire [0:0] cby_1__1__17_left_grid_pin_17_;
  wire [0:0] cby_1__1__17_left_grid_pin_18_;
  wire [0:0] cby_1__1__17_left_grid_pin_19_;
  wire [0:0] cby_1__1__17_left_grid_pin_20_;
  wire [0:0] cby_1__1__17_left_grid_pin_21_;
  wire [0:0] cby_1__1__17_left_grid_pin_22_;
  wire [0:0] cby_1__1__17_left_grid_pin_23_;
  wire [0:0] cby_1__1__17_left_grid_pin_24_;
  wire [0:0] cby_1__1__17_left_grid_pin_25_;
  wire [0:0] cby_1__1__17_left_grid_pin_26_;
  wire [0:0] cby_1__1__17_left_grid_pin_27_;
  wire [0:0] cby_1__1__17_left_grid_pin_28_;
  wire [0:0] cby_1__1__17_left_grid_pin_29_;
  wire [0:0] cby_1__1__17_left_grid_pin_30_;
  wire [0:0] cby_1__1__17_left_grid_pin_31_;
  wire [0:0] cby_1__1__18_ccff_tail;
  wire [0:29] cby_1__1__18_chany_bottom_out;
  wire [0:29] cby_1__1__18_chany_top_out;
  wire [0:0] cby_1__1__18_left_grid_pin_16_;
  wire [0:0] cby_1__1__18_left_grid_pin_17_;
  wire [0:0] cby_1__1__18_left_grid_pin_18_;
  wire [0:0] cby_1__1__18_left_grid_pin_19_;
  wire [0:0] cby_1__1__18_left_grid_pin_20_;
  wire [0:0] cby_1__1__18_left_grid_pin_21_;
  wire [0:0] cby_1__1__18_left_grid_pin_22_;
  wire [0:0] cby_1__1__18_left_grid_pin_23_;
  wire [0:0] cby_1__1__18_left_grid_pin_24_;
  wire [0:0] cby_1__1__18_left_grid_pin_25_;
  wire [0:0] cby_1__1__18_left_grid_pin_26_;
  wire [0:0] cby_1__1__18_left_grid_pin_27_;
  wire [0:0] cby_1__1__18_left_grid_pin_28_;
  wire [0:0] cby_1__1__18_left_grid_pin_29_;
  wire [0:0] cby_1__1__18_left_grid_pin_30_;
  wire [0:0] cby_1__1__18_left_grid_pin_31_;
  wire [0:0] cby_1__1__19_ccff_tail;
  wire [0:29] cby_1__1__19_chany_bottom_out;
  wire [0:29] cby_1__1__19_chany_top_out;
  wire [0:0] cby_1__1__19_left_grid_pin_16_;
  wire [0:0] cby_1__1__19_left_grid_pin_17_;
  wire [0:0] cby_1__1__19_left_grid_pin_18_;
  wire [0:0] cby_1__1__19_left_grid_pin_19_;
  wire [0:0] cby_1__1__19_left_grid_pin_20_;
  wire [0:0] cby_1__1__19_left_grid_pin_21_;
  wire [0:0] cby_1__1__19_left_grid_pin_22_;
  wire [0:0] cby_1__1__19_left_grid_pin_23_;
  wire [0:0] cby_1__1__19_left_grid_pin_24_;
  wire [0:0] cby_1__1__19_left_grid_pin_25_;
  wire [0:0] cby_1__1__19_left_grid_pin_26_;
  wire [0:0] cby_1__1__19_left_grid_pin_27_;
  wire [0:0] cby_1__1__19_left_grid_pin_28_;
  wire [0:0] cby_1__1__19_left_grid_pin_29_;
  wire [0:0] cby_1__1__19_left_grid_pin_30_;
  wire [0:0] cby_1__1__19_left_grid_pin_31_;
  wire [0:0] cby_1__1__1_ccff_tail;
  wire [0:29] cby_1__1__1_chany_bottom_out;
  wire [0:29] cby_1__1__1_chany_top_out;
  wire [0:0] cby_1__1__1_left_grid_pin_16_;
  wire [0:0] cby_1__1__1_left_grid_pin_17_;
  wire [0:0] cby_1__1__1_left_grid_pin_18_;
  wire [0:0] cby_1__1__1_left_grid_pin_19_;
  wire [0:0] cby_1__1__1_left_grid_pin_20_;
  wire [0:0] cby_1__1__1_left_grid_pin_21_;
  wire [0:0] cby_1__1__1_left_grid_pin_22_;
  wire [0:0] cby_1__1__1_left_grid_pin_23_;
  wire [0:0] cby_1__1__1_left_grid_pin_24_;
  wire [0:0] cby_1__1__1_left_grid_pin_25_;
  wire [0:0] cby_1__1__1_left_grid_pin_26_;
  wire [0:0] cby_1__1__1_left_grid_pin_27_;
  wire [0:0] cby_1__1__1_left_grid_pin_28_;
  wire [0:0] cby_1__1__1_left_grid_pin_29_;
  wire [0:0] cby_1__1__1_left_grid_pin_30_;
  wire [0:0] cby_1__1__1_left_grid_pin_31_;
  wire [0:0] cby_1__1__20_ccff_tail;
  wire [0:29] cby_1__1__20_chany_bottom_out;
  wire [0:29] cby_1__1__20_chany_top_out;
  wire [0:0] cby_1__1__20_left_grid_pin_16_;
  wire [0:0] cby_1__1__20_left_grid_pin_17_;
  wire [0:0] cby_1__1__20_left_grid_pin_18_;
  wire [0:0] cby_1__1__20_left_grid_pin_19_;
  wire [0:0] cby_1__1__20_left_grid_pin_20_;
  wire [0:0] cby_1__1__20_left_grid_pin_21_;
  wire [0:0] cby_1__1__20_left_grid_pin_22_;
  wire [0:0] cby_1__1__20_left_grid_pin_23_;
  wire [0:0] cby_1__1__20_left_grid_pin_24_;
  wire [0:0] cby_1__1__20_left_grid_pin_25_;
  wire [0:0] cby_1__1__20_left_grid_pin_26_;
  wire [0:0] cby_1__1__20_left_grid_pin_27_;
  wire [0:0] cby_1__1__20_left_grid_pin_28_;
  wire [0:0] cby_1__1__20_left_grid_pin_29_;
  wire [0:0] cby_1__1__20_left_grid_pin_30_;
  wire [0:0] cby_1__1__20_left_grid_pin_31_;
  wire [0:0] cby_1__1__21_ccff_tail;
  wire [0:29] cby_1__1__21_chany_bottom_out;
  wire [0:29] cby_1__1__21_chany_top_out;
  wire [0:0] cby_1__1__21_left_grid_pin_16_;
  wire [0:0] cby_1__1__21_left_grid_pin_17_;
  wire [0:0] cby_1__1__21_left_grid_pin_18_;
  wire [0:0] cby_1__1__21_left_grid_pin_19_;
  wire [0:0] cby_1__1__21_left_grid_pin_20_;
  wire [0:0] cby_1__1__21_left_grid_pin_21_;
  wire [0:0] cby_1__1__21_left_grid_pin_22_;
  wire [0:0] cby_1__1__21_left_grid_pin_23_;
  wire [0:0] cby_1__1__21_left_grid_pin_24_;
  wire [0:0] cby_1__1__21_left_grid_pin_25_;
  wire [0:0] cby_1__1__21_left_grid_pin_26_;
  wire [0:0] cby_1__1__21_left_grid_pin_27_;
  wire [0:0] cby_1__1__21_left_grid_pin_28_;
  wire [0:0] cby_1__1__21_left_grid_pin_29_;
  wire [0:0] cby_1__1__21_left_grid_pin_30_;
  wire [0:0] cby_1__1__21_left_grid_pin_31_;
  wire [0:0] cby_1__1__22_ccff_tail;
  wire [0:29] cby_1__1__22_chany_bottom_out;
  wire [0:29] cby_1__1__22_chany_top_out;
  wire [0:0] cby_1__1__22_left_grid_pin_16_;
  wire [0:0] cby_1__1__22_left_grid_pin_17_;
  wire [0:0] cby_1__1__22_left_grid_pin_18_;
  wire [0:0] cby_1__1__22_left_grid_pin_19_;
  wire [0:0] cby_1__1__22_left_grid_pin_20_;
  wire [0:0] cby_1__1__22_left_grid_pin_21_;
  wire [0:0] cby_1__1__22_left_grid_pin_22_;
  wire [0:0] cby_1__1__22_left_grid_pin_23_;
  wire [0:0] cby_1__1__22_left_grid_pin_24_;
  wire [0:0] cby_1__1__22_left_grid_pin_25_;
  wire [0:0] cby_1__1__22_left_grid_pin_26_;
  wire [0:0] cby_1__1__22_left_grid_pin_27_;
  wire [0:0] cby_1__1__22_left_grid_pin_28_;
  wire [0:0] cby_1__1__22_left_grid_pin_29_;
  wire [0:0] cby_1__1__22_left_grid_pin_30_;
  wire [0:0] cby_1__1__22_left_grid_pin_31_;
  wire [0:0] cby_1__1__23_ccff_tail;
  wire [0:29] cby_1__1__23_chany_bottom_out;
  wire [0:29] cby_1__1__23_chany_top_out;
  wire [0:0] cby_1__1__23_left_grid_pin_16_;
  wire [0:0] cby_1__1__23_left_grid_pin_17_;
  wire [0:0] cby_1__1__23_left_grid_pin_18_;
  wire [0:0] cby_1__1__23_left_grid_pin_19_;
  wire [0:0] cby_1__1__23_left_grid_pin_20_;
  wire [0:0] cby_1__1__23_left_grid_pin_21_;
  wire [0:0] cby_1__1__23_left_grid_pin_22_;
  wire [0:0] cby_1__1__23_left_grid_pin_23_;
  wire [0:0] cby_1__1__23_left_grid_pin_24_;
  wire [0:0] cby_1__1__23_left_grid_pin_25_;
  wire [0:0] cby_1__1__23_left_grid_pin_26_;
  wire [0:0] cby_1__1__23_left_grid_pin_27_;
  wire [0:0] cby_1__1__23_left_grid_pin_28_;
  wire [0:0] cby_1__1__23_left_grid_pin_29_;
  wire [0:0] cby_1__1__23_left_grid_pin_30_;
  wire [0:0] cby_1__1__23_left_grid_pin_31_;
  wire [0:0] cby_1__1__24_ccff_tail;
  wire [0:29] cby_1__1__24_chany_bottom_out;
  wire [0:29] cby_1__1__24_chany_top_out;
  wire [0:0] cby_1__1__24_left_grid_pin_16_;
  wire [0:0] cby_1__1__24_left_grid_pin_17_;
  wire [0:0] cby_1__1__24_left_grid_pin_18_;
  wire [0:0] cby_1__1__24_left_grid_pin_19_;
  wire [0:0] cby_1__1__24_left_grid_pin_20_;
  wire [0:0] cby_1__1__24_left_grid_pin_21_;
  wire [0:0] cby_1__1__24_left_grid_pin_22_;
  wire [0:0] cby_1__1__24_left_grid_pin_23_;
  wire [0:0] cby_1__1__24_left_grid_pin_24_;
  wire [0:0] cby_1__1__24_left_grid_pin_25_;
  wire [0:0] cby_1__1__24_left_grid_pin_26_;
  wire [0:0] cby_1__1__24_left_grid_pin_27_;
  wire [0:0] cby_1__1__24_left_grid_pin_28_;
  wire [0:0] cby_1__1__24_left_grid_pin_29_;
  wire [0:0] cby_1__1__24_left_grid_pin_30_;
  wire [0:0] cby_1__1__24_left_grid_pin_31_;
  wire [0:0] cby_1__1__25_ccff_tail;
  wire [0:29] cby_1__1__25_chany_bottom_out;
  wire [0:29] cby_1__1__25_chany_top_out;
  wire [0:0] cby_1__1__25_left_grid_pin_16_;
  wire [0:0] cby_1__1__25_left_grid_pin_17_;
  wire [0:0] cby_1__1__25_left_grid_pin_18_;
  wire [0:0] cby_1__1__25_left_grid_pin_19_;
  wire [0:0] cby_1__1__25_left_grid_pin_20_;
  wire [0:0] cby_1__1__25_left_grid_pin_21_;
  wire [0:0] cby_1__1__25_left_grid_pin_22_;
  wire [0:0] cby_1__1__25_left_grid_pin_23_;
  wire [0:0] cby_1__1__25_left_grid_pin_24_;
  wire [0:0] cby_1__1__25_left_grid_pin_25_;
  wire [0:0] cby_1__1__25_left_grid_pin_26_;
  wire [0:0] cby_1__1__25_left_grid_pin_27_;
  wire [0:0] cby_1__1__25_left_grid_pin_28_;
  wire [0:0] cby_1__1__25_left_grid_pin_29_;
  wire [0:0] cby_1__1__25_left_grid_pin_30_;
  wire [0:0] cby_1__1__25_left_grid_pin_31_;
  wire [0:0] cby_1__1__26_ccff_tail;
  wire [0:29] cby_1__1__26_chany_bottom_out;
  wire [0:29] cby_1__1__26_chany_top_out;
  wire [0:0] cby_1__1__26_left_grid_pin_16_;
  wire [0:0] cby_1__1__26_left_grid_pin_17_;
  wire [0:0] cby_1__1__26_left_grid_pin_18_;
  wire [0:0] cby_1__1__26_left_grid_pin_19_;
  wire [0:0] cby_1__1__26_left_grid_pin_20_;
  wire [0:0] cby_1__1__26_left_grid_pin_21_;
  wire [0:0] cby_1__1__26_left_grid_pin_22_;
  wire [0:0] cby_1__1__26_left_grid_pin_23_;
  wire [0:0] cby_1__1__26_left_grid_pin_24_;
  wire [0:0] cby_1__1__26_left_grid_pin_25_;
  wire [0:0] cby_1__1__26_left_grid_pin_26_;
  wire [0:0] cby_1__1__26_left_grid_pin_27_;
  wire [0:0] cby_1__1__26_left_grid_pin_28_;
  wire [0:0] cby_1__1__26_left_grid_pin_29_;
  wire [0:0] cby_1__1__26_left_grid_pin_30_;
  wire [0:0] cby_1__1__26_left_grid_pin_31_;
  wire [0:0] cby_1__1__27_ccff_tail;
  wire [0:29] cby_1__1__27_chany_bottom_out;
  wire [0:29] cby_1__1__27_chany_top_out;
  wire [0:0] cby_1__1__27_left_grid_pin_16_;
  wire [0:0] cby_1__1__27_left_grid_pin_17_;
  wire [0:0] cby_1__1__27_left_grid_pin_18_;
  wire [0:0] cby_1__1__27_left_grid_pin_19_;
  wire [0:0] cby_1__1__27_left_grid_pin_20_;
  wire [0:0] cby_1__1__27_left_grid_pin_21_;
  wire [0:0] cby_1__1__27_left_grid_pin_22_;
  wire [0:0] cby_1__1__27_left_grid_pin_23_;
  wire [0:0] cby_1__1__27_left_grid_pin_24_;
  wire [0:0] cby_1__1__27_left_grid_pin_25_;
  wire [0:0] cby_1__1__27_left_grid_pin_26_;
  wire [0:0] cby_1__1__27_left_grid_pin_27_;
  wire [0:0] cby_1__1__27_left_grid_pin_28_;
  wire [0:0] cby_1__1__27_left_grid_pin_29_;
  wire [0:0] cby_1__1__27_left_grid_pin_30_;
  wire [0:0] cby_1__1__27_left_grid_pin_31_;
  wire [0:0] cby_1__1__28_ccff_tail;
  wire [0:29] cby_1__1__28_chany_bottom_out;
  wire [0:29] cby_1__1__28_chany_top_out;
  wire [0:0] cby_1__1__28_left_grid_pin_16_;
  wire [0:0] cby_1__1__28_left_grid_pin_17_;
  wire [0:0] cby_1__1__28_left_grid_pin_18_;
  wire [0:0] cby_1__1__28_left_grid_pin_19_;
  wire [0:0] cby_1__1__28_left_grid_pin_20_;
  wire [0:0] cby_1__1__28_left_grid_pin_21_;
  wire [0:0] cby_1__1__28_left_grid_pin_22_;
  wire [0:0] cby_1__1__28_left_grid_pin_23_;
  wire [0:0] cby_1__1__28_left_grid_pin_24_;
  wire [0:0] cby_1__1__28_left_grid_pin_25_;
  wire [0:0] cby_1__1__28_left_grid_pin_26_;
  wire [0:0] cby_1__1__28_left_grid_pin_27_;
  wire [0:0] cby_1__1__28_left_grid_pin_28_;
  wire [0:0] cby_1__1__28_left_grid_pin_29_;
  wire [0:0] cby_1__1__28_left_grid_pin_30_;
  wire [0:0] cby_1__1__28_left_grid_pin_31_;
  wire [0:0] cby_1__1__29_ccff_tail;
  wire [0:29] cby_1__1__29_chany_bottom_out;
  wire [0:29] cby_1__1__29_chany_top_out;
  wire [0:0] cby_1__1__29_left_grid_pin_16_;
  wire [0:0] cby_1__1__29_left_grid_pin_17_;
  wire [0:0] cby_1__1__29_left_grid_pin_18_;
  wire [0:0] cby_1__1__29_left_grid_pin_19_;
  wire [0:0] cby_1__1__29_left_grid_pin_20_;
  wire [0:0] cby_1__1__29_left_grid_pin_21_;
  wire [0:0] cby_1__1__29_left_grid_pin_22_;
  wire [0:0] cby_1__1__29_left_grid_pin_23_;
  wire [0:0] cby_1__1__29_left_grid_pin_24_;
  wire [0:0] cby_1__1__29_left_grid_pin_25_;
  wire [0:0] cby_1__1__29_left_grid_pin_26_;
  wire [0:0] cby_1__1__29_left_grid_pin_27_;
  wire [0:0] cby_1__1__29_left_grid_pin_28_;
  wire [0:0] cby_1__1__29_left_grid_pin_29_;
  wire [0:0] cby_1__1__29_left_grid_pin_30_;
  wire [0:0] cby_1__1__29_left_grid_pin_31_;
  wire [0:0] cby_1__1__2_ccff_tail;
  wire [0:29] cby_1__1__2_chany_bottom_out;
  wire [0:29] cby_1__1__2_chany_top_out;
  wire [0:0] cby_1__1__2_left_grid_pin_16_;
  wire [0:0] cby_1__1__2_left_grid_pin_17_;
  wire [0:0] cby_1__1__2_left_grid_pin_18_;
  wire [0:0] cby_1__1__2_left_grid_pin_19_;
  wire [0:0] cby_1__1__2_left_grid_pin_20_;
  wire [0:0] cby_1__1__2_left_grid_pin_21_;
  wire [0:0] cby_1__1__2_left_grid_pin_22_;
  wire [0:0] cby_1__1__2_left_grid_pin_23_;
  wire [0:0] cby_1__1__2_left_grid_pin_24_;
  wire [0:0] cby_1__1__2_left_grid_pin_25_;
  wire [0:0] cby_1__1__2_left_grid_pin_26_;
  wire [0:0] cby_1__1__2_left_grid_pin_27_;
  wire [0:0] cby_1__1__2_left_grid_pin_28_;
  wire [0:0] cby_1__1__2_left_grid_pin_29_;
  wire [0:0] cby_1__1__2_left_grid_pin_30_;
  wire [0:0] cby_1__1__2_left_grid_pin_31_;
  wire [0:0] cby_1__1__30_ccff_tail;
  wire [0:29] cby_1__1__30_chany_bottom_out;
  wire [0:29] cby_1__1__30_chany_top_out;
  wire [0:0] cby_1__1__30_left_grid_pin_16_;
  wire [0:0] cby_1__1__30_left_grid_pin_17_;
  wire [0:0] cby_1__1__30_left_grid_pin_18_;
  wire [0:0] cby_1__1__30_left_grid_pin_19_;
  wire [0:0] cby_1__1__30_left_grid_pin_20_;
  wire [0:0] cby_1__1__30_left_grid_pin_21_;
  wire [0:0] cby_1__1__30_left_grid_pin_22_;
  wire [0:0] cby_1__1__30_left_grid_pin_23_;
  wire [0:0] cby_1__1__30_left_grid_pin_24_;
  wire [0:0] cby_1__1__30_left_grid_pin_25_;
  wire [0:0] cby_1__1__30_left_grid_pin_26_;
  wire [0:0] cby_1__1__30_left_grid_pin_27_;
  wire [0:0] cby_1__1__30_left_grid_pin_28_;
  wire [0:0] cby_1__1__30_left_grid_pin_29_;
  wire [0:0] cby_1__1__30_left_grid_pin_30_;
  wire [0:0] cby_1__1__30_left_grid_pin_31_;
  wire [0:0] cby_1__1__31_ccff_tail;
  wire [0:29] cby_1__1__31_chany_bottom_out;
  wire [0:29] cby_1__1__31_chany_top_out;
  wire [0:0] cby_1__1__31_left_grid_pin_16_;
  wire [0:0] cby_1__1__31_left_grid_pin_17_;
  wire [0:0] cby_1__1__31_left_grid_pin_18_;
  wire [0:0] cby_1__1__31_left_grid_pin_19_;
  wire [0:0] cby_1__1__31_left_grid_pin_20_;
  wire [0:0] cby_1__1__31_left_grid_pin_21_;
  wire [0:0] cby_1__1__31_left_grid_pin_22_;
  wire [0:0] cby_1__1__31_left_grid_pin_23_;
  wire [0:0] cby_1__1__31_left_grid_pin_24_;
  wire [0:0] cby_1__1__31_left_grid_pin_25_;
  wire [0:0] cby_1__1__31_left_grid_pin_26_;
  wire [0:0] cby_1__1__31_left_grid_pin_27_;
  wire [0:0] cby_1__1__31_left_grid_pin_28_;
  wire [0:0] cby_1__1__31_left_grid_pin_29_;
  wire [0:0] cby_1__1__31_left_grid_pin_30_;
  wire [0:0] cby_1__1__31_left_grid_pin_31_;
  wire [0:0] cby_1__1__32_ccff_tail;
  wire [0:29] cby_1__1__32_chany_bottom_out;
  wire [0:29] cby_1__1__32_chany_top_out;
  wire [0:0] cby_1__1__32_left_grid_pin_16_;
  wire [0:0] cby_1__1__32_left_grid_pin_17_;
  wire [0:0] cby_1__1__32_left_grid_pin_18_;
  wire [0:0] cby_1__1__32_left_grid_pin_19_;
  wire [0:0] cby_1__1__32_left_grid_pin_20_;
  wire [0:0] cby_1__1__32_left_grid_pin_21_;
  wire [0:0] cby_1__1__32_left_grid_pin_22_;
  wire [0:0] cby_1__1__32_left_grid_pin_23_;
  wire [0:0] cby_1__1__32_left_grid_pin_24_;
  wire [0:0] cby_1__1__32_left_grid_pin_25_;
  wire [0:0] cby_1__1__32_left_grid_pin_26_;
  wire [0:0] cby_1__1__32_left_grid_pin_27_;
  wire [0:0] cby_1__1__32_left_grid_pin_28_;
  wire [0:0] cby_1__1__32_left_grid_pin_29_;
  wire [0:0] cby_1__1__32_left_grid_pin_30_;
  wire [0:0] cby_1__1__32_left_grid_pin_31_;
  wire [0:0] cby_1__1__33_ccff_tail;
  wire [0:29] cby_1__1__33_chany_bottom_out;
  wire [0:29] cby_1__1__33_chany_top_out;
  wire [0:0] cby_1__1__33_left_grid_pin_16_;
  wire [0:0] cby_1__1__33_left_grid_pin_17_;
  wire [0:0] cby_1__1__33_left_grid_pin_18_;
  wire [0:0] cby_1__1__33_left_grid_pin_19_;
  wire [0:0] cby_1__1__33_left_grid_pin_20_;
  wire [0:0] cby_1__1__33_left_grid_pin_21_;
  wire [0:0] cby_1__1__33_left_grid_pin_22_;
  wire [0:0] cby_1__1__33_left_grid_pin_23_;
  wire [0:0] cby_1__1__33_left_grid_pin_24_;
  wire [0:0] cby_1__1__33_left_grid_pin_25_;
  wire [0:0] cby_1__1__33_left_grid_pin_26_;
  wire [0:0] cby_1__1__33_left_grid_pin_27_;
  wire [0:0] cby_1__1__33_left_grid_pin_28_;
  wire [0:0] cby_1__1__33_left_grid_pin_29_;
  wire [0:0] cby_1__1__33_left_grid_pin_30_;
  wire [0:0] cby_1__1__33_left_grid_pin_31_;
  wire [0:0] cby_1__1__34_ccff_tail;
  wire [0:29] cby_1__1__34_chany_bottom_out;
  wire [0:29] cby_1__1__34_chany_top_out;
  wire [0:0] cby_1__1__34_left_grid_pin_16_;
  wire [0:0] cby_1__1__34_left_grid_pin_17_;
  wire [0:0] cby_1__1__34_left_grid_pin_18_;
  wire [0:0] cby_1__1__34_left_grid_pin_19_;
  wire [0:0] cby_1__1__34_left_grid_pin_20_;
  wire [0:0] cby_1__1__34_left_grid_pin_21_;
  wire [0:0] cby_1__1__34_left_grid_pin_22_;
  wire [0:0] cby_1__1__34_left_grid_pin_23_;
  wire [0:0] cby_1__1__34_left_grid_pin_24_;
  wire [0:0] cby_1__1__34_left_grid_pin_25_;
  wire [0:0] cby_1__1__34_left_grid_pin_26_;
  wire [0:0] cby_1__1__34_left_grid_pin_27_;
  wire [0:0] cby_1__1__34_left_grid_pin_28_;
  wire [0:0] cby_1__1__34_left_grid_pin_29_;
  wire [0:0] cby_1__1__34_left_grid_pin_30_;
  wire [0:0] cby_1__1__34_left_grid_pin_31_;
  wire [0:0] cby_1__1__35_ccff_tail;
  wire [0:29] cby_1__1__35_chany_bottom_out;
  wire [0:29] cby_1__1__35_chany_top_out;
  wire [0:0] cby_1__1__35_left_grid_pin_16_;
  wire [0:0] cby_1__1__35_left_grid_pin_17_;
  wire [0:0] cby_1__1__35_left_grid_pin_18_;
  wire [0:0] cby_1__1__35_left_grid_pin_19_;
  wire [0:0] cby_1__1__35_left_grid_pin_20_;
  wire [0:0] cby_1__1__35_left_grid_pin_21_;
  wire [0:0] cby_1__1__35_left_grid_pin_22_;
  wire [0:0] cby_1__1__35_left_grid_pin_23_;
  wire [0:0] cby_1__1__35_left_grid_pin_24_;
  wire [0:0] cby_1__1__35_left_grid_pin_25_;
  wire [0:0] cby_1__1__35_left_grid_pin_26_;
  wire [0:0] cby_1__1__35_left_grid_pin_27_;
  wire [0:0] cby_1__1__35_left_grid_pin_28_;
  wire [0:0] cby_1__1__35_left_grid_pin_29_;
  wire [0:0] cby_1__1__35_left_grid_pin_30_;
  wire [0:0] cby_1__1__35_left_grid_pin_31_;
  wire [0:0] cby_1__1__36_ccff_tail;
  wire [0:29] cby_1__1__36_chany_bottom_out;
  wire [0:29] cby_1__1__36_chany_top_out;
  wire [0:0] cby_1__1__36_left_grid_pin_16_;
  wire [0:0] cby_1__1__36_left_grid_pin_17_;
  wire [0:0] cby_1__1__36_left_grid_pin_18_;
  wire [0:0] cby_1__1__36_left_grid_pin_19_;
  wire [0:0] cby_1__1__36_left_grid_pin_20_;
  wire [0:0] cby_1__1__36_left_grid_pin_21_;
  wire [0:0] cby_1__1__36_left_grid_pin_22_;
  wire [0:0] cby_1__1__36_left_grid_pin_23_;
  wire [0:0] cby_1__1__36_left_grid_pin_24_;
  wire [0:0] cby_1__1__36_left_grid_pin_25_;
  wire [0:0] cby_1__1__36_left_grid_pin_26_;
  wire [0:0] cby_1__1__36_left_grid_pin_27_;
  wire [0:0] cby_1__1__36_left_grid_pin_28_;
  wire [0:0] cby_1__1__36_left_grid_pin_29_;
  wire [0:0] cby_1__1__36_left_grid_pin_30_;
  wire [0:0] cby_1__1__36_left_grid_pin_31_;
  wire [0:0] cby_1__1__37_ccff_tail;
  wire [0:29] cby_1__1__37_chany_bottom_out;
  wire [0:29] cby_1__1__37_chany_top_out;
  wire [0:0] cby_1__1__37_left_grid_pin_16_;
  wire [0:0] cby_1__1__37_left_grid_pin_17_;
  wire [0:0] cby_1__1__37_left_grid_pin_18_;
  wire [0:0] cby_1__1__37_left_grid_pin_19_;
  wire [0:0] cby_1__1__37_left_grid_pin_20_;
  wire [0:0] cby_1__1__37_left_grid_pin_21_;
  wire [0:0] cby_1__1__37_left_grid_pin_22_;
  wire [0:0] cby_1__1__37_left_grid_pin_23_;
  wire [0:0] cby_1__1__37_left_grid_pin_24_;
  wire [0:0] cby_1__1__37_left_grid_pin_25_;
  wire [0:0] cby_1__1__37_left_grid_pin_26_;
  wire [0:0] cby_1__1__37_left_grid_pin_27_;
  wire [0:0] cby_1__1__37_left_grid_pin_28_;
  wire [0:0] cby_1__1__37_left_grid_pin_29_;
  wire [0:0] cby_1__1__37_left_grid_pin_30_;
  wire [0:0] cby_1__1__37_left_grid_pin_31_;
  wire [0:0] cby_1__1__38_ccff_tail;
  wire [0:29] cby_1__1__38_chany_bottom_out;
  wire [0:29] cby_1__1__38_chany_top_out;
  wire [0:0] cby_1__1__38_left_grid_pin_16_;
  wire [0:0] cby_1__1__38_left_grid_pin_17_;
  wire [0:0] cby_1__1__38_left_grid_pin_18_;
  wire [0:0] cby_1__1__38_left_grid_pin_19_;
  wire [0:0] cby_1__1__38_left_grid_pin_20_;
  wire [0:0] cby_1__1__38_left_grid_pin_21_;
  wire [0:0] cby_1__1__38_left_grid_pin_22_;
  wire [0:0] cby_1__1__38_left_grid_pin_23_;
  wire [0:0] cby_1__1__38_left_grid_pin_24_;
  wire [0:0] cby_1__1__38_left_grid_pin_25_;
  wire [0:0] cby_1__1__38_left_grid_pin_26_;
  wire [0:0] cby_1__1__38_left_grid_pin_27_;
  wire [0:0] cby_1__1__38_left_grid_pin_28_;
  wire [0:0] cby_1__1__38_left_grid_pin_29_;
  wire [0:0] cby_1__1__38_left_grid_pin_30_;
  wire [0:0] cby_1__1__38_left_grid_pin_31_;
  wire [0:0] cby_1__1__39_ccff_tail;
  wire [0:29] cby_1__1__39_chany_bottom_out;
  wire [0:29] cby_1__1__39_chany_top_out;
  wire [0:0] cby_1__1__39_left_grid_pin_16_;
  wire [0:0] cby_1__1__39_left_grid_pin_17_;
  wire [0:0] cby_1__1__39_left_grid_pin_18_;
  wire [0:0] cby_1__1__39_left_grid_pin_19_;
  wire [0:0] cby_1__1__39_left_grid_pin_20_;
  wire [0:0] cby_1__1__39_left_grid_pin_21_;
  wire [0:0] cby_1__1__39_left_grid_pin_22_;
  wire [0:0] cby_1__1__39_left_grid_pin_23_;
  wire [0:0] cby_1__1__39_left_grid_pin_24_;
  wire [0:0] cby_1__1__39_left_grid_pin_25_;
  wire [0:0] cby_1__1__39_left_grid_pin_26_;
  wire [0:0] cby_1__1__39_left_grid_pin_27_;
  wire [0:0] cby_1__1__39_left_grid_pin_28_;
  wire [0:0] cby_1__1__39_left_grid_pin_29_;
  wire [0:0] cby_1__1__39_left_grid_pin_30_;
  wire [0:0] cby_1__1__39_left_grid_pin_31_;
  wire [0:0] cby_1__1__3_ccff_tail;
  wire [0:29] cby_1__1__3_chany_bottom_out;
  wire [0:29] cby_1__1__3_chany_top_out;
  wire [0:0] cby_1__1__3_left_grid_pin_16_;
  wire [0:0] cby_1__1__3_left_grid_pin_17_;
  wire [0:0] cby_1__1__3_left_grid_pin_18_;
  wire [0:0] cby_1__1__3_left_grid_pin_19_;
  wire [0:0] cby_1__1__3_left_grid_pin_20_;
  wire [0:0] cby_1__1__3_left_grid_pin_21_;
  wire [0:0] cby_1__1__3_left_grid_pin_22_;
  wire [0:0] cby_1__1__3_left_grid_pin_23_;
  wire [0:0] cby_1__1__3_left_grid_pin_24_;
  wire [0:0] cby_1__1__3_left_grid_pin_25_;
  wire [0:0] cby_1__1__3_left_grid_pin_26_;
  wire [0:0] cby_1__1__3_left_grid_pin_27_;
  wire [0:0] cby_1__1__3_left_grid_pin_28_;
  wire [0:0] cby_1__1__3_left_grid_pin_29_;
  wire [0:0] cby_1__1__3_left_grid_pin_30_;
  wire [0:0] cby_1__1__3_left_grid_pin_31_;
  wire [0:0] cby_1__1__40_ccff_tail;
  wire [0:29] cby_1__1__40_chany_bottom_out;
  wire [0:29] cby_1__1__40_chany_top_out;
  wire [0:0] cby_1__1__40_left_grid_pin_16_;
  wire [0:0] cby_1__1__40_left_grid_pin_17_;
  wire [0:0] cby_1__1__40_left_grid_pin_18_;
  wire [0:0] cby_1__1__40_left_grid_pin_19_;
  wire [0:0] cby_1__1__40_left_grid_pin_20_;
  wire [0:0] cby_1__1__40_left_grid_pin_21_;
  wire [0:0] cby_1__1__40_left_grid_pin_22_;
  wire [0:0] cby_1__1__40_left_grid_pin_23_;
  wire [0:0] cby_1__1__40_left_grid_pin_24_;
  wire [0:0] cby_1__1__40_left_grid_pin_25_;
  wire [0:0] cby_1__1__40_left_grid_pin_26_;
  wire [0:0] cby_1__1__40_left_grid_pin_27_;
  wire [0:0] cby_1__1__40_left_grid_pin_28_;
  wire [0:0] cby_1__1__40_left_grid_pin_29_;
  wire [0:0] cby_1__1__40_left_grid_pin_30_;
  wire [0:0] cby_1__1__40_left_grid_pin_31_;
  wire [0:0] cby_1__1__41_ccff_tail;
  wire [0:29] cby_1__1__41_chany_bottom_out;
  wire [0:29] cby_1__1__41_chany_top_out;
  wire [0:0] cby_1__1__41_left_grid_pin_16_;
  wire [0:0] cby_1__1__41_left_grid_pin_17_;
  wire [0:0] cby_1__1__41_left_grid_pin_18_;
  wire [0:0] cby_1__1__41_left_grid_pin_19_;
  wire [0:0] cby_1__1__41_left_grid_pin_20_;
  wire [0:0] cby_1__1__41_left_grid_pin_21_;
  wire [0:0] cby_1__1__41_left_grid_pin_22_;
  wire [0:0] cby_1__1__41_left_grid_pin_23_;
  wire [0:0] cby_1__1__41_left_grid_pin_24_;
  wire [0:0] cby_1__1__41_left_grid_pin_25_;
  wire [0:0] cby_1__1__41_left_grid_pin_26_;
  wire [0:0] cby_1__1__41_left_grid_pin_27_;
  wire [0:0] cby_1__1__41_left_grid_pin_28_;
  wire [0:0] cby_1__1__41_left_grid_pin_29_;
  wire [0:0] cby_1__1__41_left_grid_pin_30_;
  wire [0:0] cby_1__1__41_left_grid_pin_31_;
  wire [0:0] cby_1__1__42_ccff_tail;
  wire [0:29] cby_1__1__42_chany_bottom_out;
  wire [0:29] cby_1__1__42_chany_top_out;
  wire [0:0] cby_1__1__42_left_grid_pin_16_;
  wire [0:0] cby_1__1__42_left_grid_pin_17_;
  wire [0:0] cby_1__1__42_left_grid_pin_18_;
  wire [0:0] cby_1__1__42_left_grid_pin_19_;
  wire [0:0] cby_1__1__42_left_grid_pin_20_;
  wire [0:0] cby_1__1__42_left_grid_pin_21_;
  wire [0:0] cby_1__1__42_left_grid_pin_22_;
  wire [0:0] cby_1__1__42_left_grid_pin_23_;
  wire [0:0] cby_1__1__42_left_grid_pin_24_;
  wire [0:0] cby_1__1__42_left_grid_pin_25_;
  wire [0:0] cby_1__1__42_left_grid_pin_26_;
  wire [0:0] cby_1__1__42_left_grid_pin_27_;
  wire [0:0] cby_1__1__42_left_grid_pin_28_;
  wire [0:0] cby_1__1__42_left_grid_pin_29_;
  wire [0:0] cby_1__1__42_left_grid_pin_30_;
  wire [0:0] cby_1__1__42_left_grid_pin_31_;
  wire [0:0] cby_1__1__43_ccff_tail;
  wire [0:29] cby_1__1__43_chany_bottom_out;
  wire [0:29] cby_1__1__43_chany_top_out;
  wire [0:0] cby_1__1__43_left_grid_pin_16_;
  wire [0:0] cby_1__1__43_left_grid_pin_17_;
  wire [0:0] cby_1__1__43_left_grid_pin_18_;
  wire [0:0] cby_1__1__43_left_grid_pin_19_;
  wire [0:0] cby_1__1__43_left_grid_pin_20_;
  wire [0:0] cby_1__1__43_left_grid_pin_21_;
  wire [0:0] cby_1__1__43_left_grid_pin_22_;
  wire [0:0] cby_1__1__43_left_grid_pin_23_;
  wire [0:0] cby_1__1__43_left_grid_pin_24_;
  wire [0:0] cby_1__1__43_left_grid_pin_25_;
  wire [0:0] cby_1__1__43_left_grid_pin_26_;
  wire [0:0] cby_1__1__43_left_grid_pin_27_;
  wire [0:0] cby_1__1__43_left_grid_pin_28_;
  wire [0:0] cby_1__1__43_left_grid_pin_29_;
  wire [0:0] cby_1__1__43_left_grid_pin_30_;
  wire [0:0] cby_1__1__43_left_grid_pin_31_;
  wire [0:0] cby_1__1__44_ccff_tail;
  wire [0:29] cby_1__1__44_chany_bottom_out;
  wire [0:29] cby_1__1__44_chany_top_out;
  wire [0:0] cby_1__1__44_left_grid_pin_16_;
  wire [0:0] cby_1__1__44_left_grid_pin_17_;
  wire [0:0] cby_1__1__44_left_grid_pin_18_;
  wire [0:0] cby_1__1__44_left_grid_pin_19_;
  wire [0:0] cby_1__1__44_left_grid_pin_20_;
  wire [0:0] cby_1__1__44_left_grid_pin_21_;
  wire [0:0] cby_1__1__44_left_grid_pin_22_;
  wire [0:0] cby_1__1__44_left_grid_pin_23_;
  wire [0:0] cby_1__1__44_left_grid_pin_24_;
  wire [0:0] cby_1__1__44_left_grid_pin_25_;
  wire [0:0] cby_1__1__44_left_grid_pin_26_;
  wire [0:0] cby_1__1__44_left_grid_pin_27_;
  wire [0:0] cby_1__1__44_left_grid_pin_28_;
  wire [0:0] cby_1__1__44_left_grid_pin_29_;
  wire [0:0] cby_1__1__44_left_grid_pin_30_;
  wire [0:0] cby_1__1__44_left_grid_pin_31_;
  wire [0:0] cby_1__1__45_ccff_tail;
  wire [0:29] cby_1__1__45_chany_bottom_out;
  wire [0:29] cby_1__1__45_chany_top_out;
  wire [0:0] cby_1__1__45_left_grid_pin_16_;
  wire [0:0] cby_1__1__45_left_grid_pin_17_;
  wire [0:0] cby_1__1__45_left_grid_pin_18_;
  wire [0:0] cby_1__1__45_left_grid_pin_19_;
  wire [0:0] cby_1__1__45_left_grid_pin_20_;
  wire [0:0] cby_1__1__45_left_grid_pin_21_;
  wire [0:0] cby_1__1__45_left_grid_pin_22_;
  wire [0:0] cby_1__1__45_left_grid_pin_23_;
  wire [0:0] cby_1__1__45_left_grid_pin_24_;
  wire [0:0] cby_1__1__45_left_grid_pin_25_;
  wire [0:0] cby_1__1__45_left_grid_pin_26_;
  wire [0:0] cby_1__1__45_left_grid_pin_27_;
  wire [0:0] cby_1__1__45_left_grid_pin_28_;
  wire [0:0] cby_1__1__45_left_grid_pin_29_;
  wire [0:0] cby_1__1__45_left_grid_pin_30_;
  wire [0:0] cby_1__1__45_left_grid_pin_31_;
  wire [0:0] cby_1__1__46_ccff_tail;
  wire [0:29] cby_1__1__46_chany_bottom_out;
  wire [0:29] cby_1__1__46_chany_top_out;
  wire [0:0] cby_1__1__46_left_grid_pin_16_;
  wire [0:0] cby_1__1__46_left_grid_pin_17_;
  wire [0:0] cby_1__1__46_left_grid_pin_18_;
  wire [0:0] cby_1__1__46_left_grid_pin_19_;
  wire [0:0] cby_1__1__46_left_grid_pin_20_;
  wire [0:0] cby_1__1__46_left_grid_pin_21_;
  wire [0:0] cby_1__1__46_left_grid_pin_22_;
  wire [0:0] cby_1__1__46_left_grid_pin_23_;
  wire [0:0] cby_1__1__46_left_grid_pin_24_;
  wire [0:0] cby_1__1__46_left_grid_pin_25_;
  wire [0:0] cby_1__1__46_left_grid_pin_26_;
  wire [0:0] cby_1__1__46_left_grid_pin_27_;
  wire [0:0] cby_1__1__46_left_grid_pin_28_;
  wire [0:0] cby_1__1__46_left_grid_pin_29_;
  wire [0:0] cby_1__1__46_left_grid_pin_30_;
  wire [0:0] cby_1__1__46_left_grid_pin_31_;
  wire [0:0] cby_1__1__47_ccff_tail;
  wire [0:29] cby_1__1__47_chany_bottom_out;
  wire [0:29] cby_1__1__47_chany_top_out;
  wire [0:0] cby_1__1__47_left_grid_pin_16_;
  wire [0:0] cby_1__1__47_left_grid_pin_17_;
  wire [0:0] cby_1__1__47_left_grid_pin_18_;
  wire [0:0] cby_1__1__47_left_grid_pin_19_;
  wire [0:0] cby_1__1__47_left_grid_pin_20_;
  wire [0:0] cby_1__1__47_left_grid_pin_21_;
  wire [0:0] cby_1__1__47_left_grid_pin_22_;
  wire [0:0] cby_1__1__47_left_grid_pin_23_;
  wire [0:0] cby_1__1__47_left_grid_pin_24_;
  wire [0:0] cby_1__1__47_left_grid_pin_25_;
  wire [0:0] cby_1__1__47_left_grid_pin_26_;
  wire [0:0] cby_1__1__47_left_grid_pin_27_;
  wire [0:0] cby_1__1__47_left_grid_pin_28_;
  wire [0:0] cby_1__1__47_left_grid_pin_29_;
  wire [0:0] cby_1__1__47_left_grid_pin_30_;
  wire [0:0] cby_1__1__47_left_grid_pin_31_;
  wire [0:0] cby_1__1__48_ccff_tail;
  wire [0:29] cby_1__1__48_chany_bottom_out;
  wire [0:29] cby_1__1__48_chany_top_out;
  wire [0:0] cby_1__1__48_left_grid_pin_16_;
  wire [0:0] cby_1__1__48_left_grid_pin_17_;
  wire [0:0] cby_1__1__48_left_grid_pin_18_;
  wire [0:0] cby_1__1__48_left_grid_pin_19_;
  wire [0:0] cby_1__1__48_left_grid_pin_20_;
  wire [0:0] cby_1__1__48_left_grid_pin_21_;
  wire [0:0] cby_1__1__48_left_grid_pin_22_;
  wire [0:0] cby_1__1__48_left_grid_pin_23_;
  wire [0:0] cby_1__1__48_left_grid_pin_24_;
  wire [0:0] cby_1__1__48_left_grid_pin_25_;
  wire [0:0] cby_1__1__48_left_grid_pin_26_;
  wire [0:0] cby_1__1__48_left_grid_pin_27_;
  wire [0:0] cby_1__1__48_left_grid_pin_28_;
  wire [0:0] cby_1__1__48_left_grid_pin_29_;
  wire [0:0] cby_1__1__48_left_grid_pin_30_;
  wire [0:0] cby_1__1__48_left_grid_pin_31_;
  wire [0:0] cby_1__1__49_ccff_tail;
  wire [0:29] cby_1__1__49_chany_bottom_out;
  wire [0:29] cby_1__1__49_chany_top_out;
  wire [0:0] cby_1__1__49_left_grid_pin_16_;
  wire [0:0] cby_1__1__49_left_grid_pin_17_;
  wire [0:0] cby_1__1__49_left_grid_pin_18_;
  wire [0:0] cby_1__1__49_left_grid_pin_19_;
  wire [0:0] cby_1__1__49_left_grid_pin_20_;
  wire [0:0] cby_1__1__49_left_grid_pin_21_;
  wire [0:0] cby_1__1__49_left_grid_pin_22_;
  wire [0:0] cby_1__1__49_left_grid_pin_23_;
  wire [0:0] cby_1__1__49_left_grid_pin_24_;
  wire [0:0] cby_1__1__49_left_grid_pin_25_;
  wire [0:0] cby_1__1__49_left_grid_pin_26_;
  wire [0:0] cby_1__1__49_left_grid_pin_27_;
  wire [0:0] cby_1__1__49_left_grid_pin_28_;
  wire [0:0] cby_1__1__49_left_grid_pin_29_;
  wire [0:0] cby_1__1__49_left_grid_pin_30_;
  wire [0:0] cby_1__1__49_left_grid_pin_31_;
  wire [0:0] cby_1__1__4_ccff_tail;
  wire [0:29] cby_1__1__4_chany_bottom_out;
  wire [0:29] cby_1__1__4_chany_top_out;
  wire [0:0] cby_1__1__4_left_grid_pin_16_;
  wire [0:0] cby_1__1__4_left_grid_pin_17_;
  wire [0:0] cby_1__1__4_left_grid_pin_18_;
  wire [0:0] cby_1__1__4_left_grid_pin_19_;
  wire [0:0] cby_1__1__4_left_grid_pin_20_;
  wire [0:0] cby_1__1__4_left_grid_pin_21_;
  wire [0:0] cby_1__1__4_left_grid_pin_22_;
  wire [0:0] cby_1__1__4_left_grid_pin_23_;
  wire [0:0] cby_1__1__4_left_grid_pin_24_;
  wire [0:0] cby_1__1__4_left_grid_pin_25_;
  wire [0:0] cby_1__1__4_left_grid_pin_26_;
  wire [0:0] cby_1__1__4_left_grid_pin_27_;
  wire [0:0] cby_1__1__4_left_grid_pin_28_;
  wire [0:0] cby_1__1__4_left_grid_pin_29_;
  wire [0:0] cby_1__1__4_left_grid_pin_30_;
  wire [0:0] cby_1__1__4_left_grid_pin_31_;
  wire [0:0] cby_1__1__50_ccff_tail;
  wire [0:29] cby_1__1__50_chany_bottom_out;
  wire [0:29] cby_1__1__50_chany_top_out;
  wire [0:0] cby_1__1__50_left_grid_pin_16_;
  wire [0:0] cby_1__1__50_left_grid_pin_17_;
  wire [0:0] cby_1__1__50_left_grid_pin_18_;
  wire [0:0] cby_1__1__50_left_grid_pin_19_;
  wire [0:0] cby_1__1__50_left_grid_pin_20_;
  wire [0:0] cby_1__1__50_left_grid_pin_21_;
  wire [0:0] cby_1__1__50_left_grid_pin_22_;
  wire [0:0] cby_1__1__50_left_grid_pin_23_;
  wire [0:0] cby_1__1__50_left_grid_pin_24_;
  wire [0:0] cby_1__1__50_left_grid_pin_25_;
  wire [0:0] cby_1__1__50_left_grid_pin_26_;
  wire [0:0] cby_1__1__50_left_grid_pin_27_;
  wire [0:0] cby_1__1__50_left_grid_pin_28_;
  wire [0:0] cby_1__1__50_left_grid_pin_29_;
  wire [0:0] cby_1__1__50_left_grid_pin_30_;
  wire [0:0] cby_1__1__50_left_grid_pin_31_;
  wire [0:0] cby_1__1__51_ccff_tail;
  wire [0:29] cby_1__1__51_chany_bottom_out;
  wire [0:29] cby_1__1__51_chany_top_out;
  wire [0:0] cby_1__1__51_left_grid_pin_16_;
  wire [0:0] cby_1__1__51_left_grid_pin_17_;
  wire [0:0] cby_1__1__51_left_grid_pin_18_;
  wire [0:0] cby_1__1__51_left_grid_pin_19_;
  wire [0:0] cby_1__1__51_left_grid_pin_20_;
  wire [0:0] cby_1__1__51_left_grid_pin_21_;
  wire [0:0] cby_1__1__51_left_grid_pin_22_;
  wire [0:0] cby_1__1__51_left_grid_pin_23_;
  wire [0:0] cby_1__1__51_left_grid_pin_24_;
  wire [0:0] cby_1__1__51_left_grid_pin_25_;
  wire [0:0] cby_1__1__51_left_grid_pin_26_;
  wire [0:0] cby_1__1__51_left_grid_pin_27_;
  wire [0:0] cby_1__1__51_left_grid_pin_28_;
  wire [0:0] cby_1__1__51_left_grid_pin_29_;
  wire [0:0] cby_1__1__51_left_grid_pin_30_;
  wire [0:0] cby_1__1__51_left_grid_pin_31_;
  wire [0:0] cby_1__1__52_ccff_tail;
  wire [0:29] cby_1__1__52_chany_bottom_out;
  wire [0:29] cby_1__1__52_chany_top_out;
  wire [0:0] cby_1__1__52_left_grid_pin_16_;
  wire [0:0] cby_1__1__52_left_grid_pin_17_;
  wire [0:0] cby_1__1__52_left_grid_pin_18_;
  wire [0:0] cby_1__1__52_left_grid_pin_19_;
  wire [0:0] cby_1__1__52_left_grid_pin_20_;
  wire [0:0] cby_1__1__52_left_grid_pin_21_;
  wire [0:0] cby_1__1__52_left_grid_pin_22_;
  wire [0:0] cby_1__1__52_left_grid_pin_23_;
  wire [0:0] cby_1__1__52_left_grid_pin_24_;
  wire [0:0] cby_1__1__52_left_grid_pin_25_;
  wire [0:0] cby_1__1__52_left_grid_pin_26_;
  wire [0:0] cby_1__1__52_left_grid_pin_27_;
  wire [0:0] cby_1__1__52_left_grid_pin_28_;
  wire [0:0] cby_1__1__52_left_grid_pin_29_;
  wire [0:0] cby_1__1__52_left_grid_pin_30_;
  wire [0:0] cby_1__1__52_left_grid_pin_31_;
  wire [0:0] cby_1__1__53_ccff_tail;
  wire [0:29] cby_1__1__53_chany_bottom_out;
  wire [0:29] cby_1__1__53_chany_top_out;
  wire [0:0] cby_1__1__53_left_grid_pin_16_;
  wire [0:0] cby_1__1__53_left_grid_pin_17_;
  wire [0:0] cby_1__1__53_left_grid_pin_18_;
  wire [0:0] cby_1__1__53_left_grid_pin_19_;
  wire [0:0] cby_1__1__53_left_grid_pin_20_;
  wire [0:0] cby_1__1__53_left_grid_pin_21_;
  wire [0:0] cby_1__1__53_left_grid_pin_22_;
  wire [0:0] cby_1__1__53_left_grid_pin_23_;
  wire [0:0] cby_1__1__53_left_grid_pin_24_;
  wire [0:0] cby_1__1__53_left_grid_pin_25_;
  wire [0:0] cby_1__1__53_left_grid_pin_26_;
  wire [0:0] cby_1__1__53_left_grid_pin_27_;
  wire [0:0] cby_1__1__53_left_grid_pin_28_;
  wire [0:0] cby_1__1__53_left_grid_pin_29_;
  wire [0:0] cby_1__1__53_left_grid_pin_30_;
  wire [0:0] cby_1__1__53_left_grid_pin_31_;
  wire [0:0] cby_1__1__54_ccff_tail;
  wire [0:29] cby_1__1__54_chany_bottom_out;
  wire [0:29] cby_1__1__54_chany_top_out;
  wire [0:0] cby_1__1__54_left_grid_pin_16_;
  wire [0:0] cby_1__1__54_left_grid_pin_17_;
  wire [0:0] cby_1__1__54_left_grid_pin_18_;
  wire [0:0] cby_1__1__54_left_grid_pin_19_;
  wire [0:0] cby_1__1__54_left_grid_pin_20_;
  wire [0:0] cby_1__1__54_left_grid_pin_21_;
  wire [0:0] cby_1__1__54_left_grid_pin_22_;
  wire [0:0] cby_1__1__54_left_grid_pin_23_;
  wire [0:0] cby_1__1__54_left_grid_pin_24_;
  wire [0:0] cby_1__1__54_left_grid_pin_25_;
  wire [0:0] cby_1__1__54_left_grid_pin_26_;
  wire [0:0] cby_1__1__54_left_grid_pin_27_;
  wire [0:0] cby_1__1__54_left_grid_pin_28_;
  wire [0:0] cby_1__1__54_left_grid_pin_29_;
  wire [0:0] cby_1__1__54_left_grid_pin_30_;
  wire [0:0] cby_1__1__54_left_grid_pin_31_;
  wire [0:0] cby_1__1__55_ccff_tail;
  wire [0:29] cby_1__1__55_chany_bottom_out;
  wire [0:29] cby_1__1__55_chany_top_out;
  wire [0:0] cby_1__1__55_left_grid_pin_16_;
  wire [0:0] cby_1__1__55_left_grid_pin_17_;
  wire [0:0] cby_1__1__55_left_grid_pin_18_;
  wire [0:0] cby_1__1__55_left_grid_pin_19_;
  wire [0:0] cby_1__1__55_left_grid_pin_20_;
  wire [0:0] cby_1__1__55_left_grid_pin_21_;
  wire [0:0] cby_1__1__55_left_grid_pin_22_;
  wire [0:0] cby_1__1__55_left_grid_pin_23_;
  wire [0:0] cby_1__1__55_left_grid_pin_24_;
  wire [0:0] cby_1__1__55_left_grid_pin_25_;
  wire [0:0] cby_1__1__55_left_grid_pin_26_;
  wire [0:0] cby_1__1__55_left_grid_pin_27_;
  wire [0:0] cby_1__1__55_left_grid_pin_28_;
  wire [0:0] cby_1__1__55_left_grid_pin_29_;
  wire [0:0] cby_1__1__55_left_grid_pin_30_;
  wire [0:0] cby_1__1__55_left_grid_pin_31_;
  wire [0:0] cby_1__1__56_ccff_tail;
  wire [0:29] cby_1__1__56_chany_bottom_out;
  wire [0:29] cby_1__1__56_chany_top_out;
  wire [0:0] cby_1__1__56_left_grid_pin_16_;
  wire [0:0] cby_1__1__56_left_grid_pin_17_;
  wire [0:0] cby_1__1__56_left_grid_pin_18_;
  wire [0:0] cby_1__1__56_left_grid_pin_19_;
  wire [0:0] cby_1__1__56_left_grid_pin_20_;
  wire [0:0] cby_1__1__56_left_grid_pin_21_;
  wire [0:0] cby_1__1__56_left_grid_pin_22_;
  wire [0:0] cby_1__1__56_left_grid_pin_23_;
  wire [0:0] cby_1__1__56_left_grid_pin_24_;
  wire [0:0] cby_1__1__56_left_grid_pin_25_;
  wire [0:0] cby_1__1__56_left_grid_pin_26_;
  wire [0:0] cby_1__1__56_left_grid_pin_27_;
  wire [0:0] cby_1__1__56_left_grid_pin_28_;
  wire [0:0] cby_1__1__56_left_grid_pin_29_;
  wire [0:0] cby_1__1__56_left_grid_pin_30_;
  wire [0:0] cby_1__1__56_left_grid_pin_31_;
  wire [0:0] cby_1__1__57_ccff_tail;
  wire [0:29] cby_1__1__57_chany_bottom_out;
  wire [0:29] cby_1__1__57_chany_top_out;
  wire [0:0] cby_1__1__57_left_grid_pin_16_;
  wire [0:0] cby_1__1__57_left_grid_pin_17_;
  wire [0:0] cby_1__1__57_left_grid_pin_18_;
  wire [0:0] cby_1__1__57_left_grid_pin_19_;
  wire [0:0] cby_1__1__57_left_grid_pin_20_;
  wire [0:0] cby_1__1__57_left_grid_pin_21_;
  wire [0:0] cby_1__1__57_left_grid_pin_22_;
  wire [0:0] cby_1__1__57_left_grid_pin_23_;
  wire [0:0] cby_1__1__57_left_grid_pin_24_;
  wire [0:0] cby_1__1__57_left_grid_pin_25_;
  wire [0:0] cby_1__1__57_left_grid_pin_26_;
  wire [0:0] cby_1__1__57_left_grid_pin_27_;
  wire [0:0] cby_1__1__57_left_grid_pin_28_;
  wire [0:0] cby_1__1__57_left_grid_pin_29_;
  wire [0:0] cby_1__1__57_left_grid_pin_30_;
  wire [0:0] cby_1__1__57_left_grid_pin_31_;
  wire [0:0] cby_1__1__58_ccff_tail;
  wire [0:29] cby_1__1__58_chany_bottom_out;
  wire [0:29] cby_1__1__58_chany_top_out;
  wire [0:0] cby_1__1__58_left_grid_pin_16_;
  wire [0:0] cby_1__1__58_left_grid_pin_17_;
  wire [0:0] cby_1__1__58_left_grid_pin_18_;
  wire [0:0] cby_1__1__58_left_grid_pin_19_;
  wire [0:0] cby_1__1__58_left_grid_pin_20_;
  wire [0:0] cby_1__1__58_left_grid_pin_21_;
  wire [0:0] cby_1__1__58_left_grid_pin_22_;
  wire [0:0] cby_1__1__58_left_grid_pin_23_;
  wire [0:0] cby_1__1__58_left_grid_pin_24_;
  wire [0:0] cby_1__1__58_left_grid_pin_25_;
  wire [0:0] cby_1__1__58_left_grid_pin_26_;
  wire [0:0] cby_1__1__58_left_grid_pin_27_;
  wire [0:0] cby_1__1__58_left_grid_pin_28_;
  wire [0:0] cby_1__1__58_left_grid_pin_29_;
  wire [0:0] cby_1__1__58_left_grid_pin_30_;
  wire [0:0] cby_1__1__58_left_grid_pin_31_;
  wire [0:0] cby_1__1__59_ccff_tail;
  wire [0:29] cby_1__1__59_chany_bottom_out;
  wire [0:29] cby_1__1__59_chany_top_out;
  wire [0:0] cby_1__1__59_left_grid_pin_16_;
  wire [0:0] cby_1__1__59_left_grid_pin_17_;
  wire [0:0] cby_1__1__59_left_grid_pin_18_;
  wire [0:0] cby_1__1__59_left_grid_pin_19_;
  wire [0:0] cby_1__1__59_left_grid_pin_20_;
  wire [0:0] cby_1__1__59_left_grid_pin_21_;
  wire [0:0] cby_1__1__59_left_grid_pin_22_;
  wire [0:0] cby_1__1__59_left_grid_pin_23_;
  wire [0:0] cby_1__1__59_left_grid_pin_24_;
  wire [0:0] cby_1__1__59_left_grid_pin_25_;
  wire [0:0] cby_1__1__59_left_grid_pin_26_;
  wire [0:0] cby_1__1__59_left_grid_pin_27_;
  wire [0:0] cby_1__1__59_left_grid_pin_28_;
  wire [0:0] cby_1__1__59_left_grid_pin_29_;
  wire [0:0] cby_1__1__59_left_grid_pin_30_;
  wire [0:0] cby_1__1__59_left_grid_pin_31_;
  wire [0:0] cby_1__1__5_ccff_tail;
  wire [0:29] cby_1__1__5_chany_bottom_out;
  wire [0:29] cby_1__1__5_chany_top_out;
  wire [0:0] cby_1__1__5_left_grid_pin_16_;
  wire [0:0] cby_1__1__5_left_grid_pin_17_;
  wire [0:0] cby_1__1__5_left_grid_pin_18_;
  wire [0:0] cby_1__1__5_left_grid_pin_19_;
  wire [0:0] cby_1__1__5_left_grid_pin_20_;
  wire [0:0] cby_1__1__5_left_grid_pin_21_;
  wire [0:0] cby_1__1__5_left_grid_pin_22_;
  wire [0:0] cby_1__1__5_left_grid_pin_23_;
  wire [0:0] cby_1__1__5_left_grid_pin_24_;
  wire [0:0] cby_1__1__5_left_grid_pin_25_;
  wire [0:0] cby_1__1__5_left_grid_pin_26_;
  wire [0:0] cby_1__1__5_left_grid_pin_27_;
  wire [0:0] cby_1__1__5_left_grid_pin_28_;
  wire [0:0] cby_1__1__5_left_grid_pin_29_;
  wire [0:0] cby_1__1__5_left_grid_pin_30_;
  wire [0:0] cby_1__1__5_left_grid_pin_31_;
  wire [0:0] cby_1__1__60_ccff_tail;
  wire [0:29] cby_1__1__60_chany_bottom_out;
  wire [0:29] cby_1__1__60_chany_top_out;
  wire [0:0] cby_1__1__60_left_grid_pin_16_;
  wire [0:0] cby_1__1__60_left_grid_pin_17_;
  wire [0:0] cby_1__1__60_left_grid_pin_18_;
  wire [0:0] cby_1__1__60_left_grid_pin_19_;
  wire [0:0] cby_1__1__60_left_grid_pin_20_;
  wire [0:0] cby_1__1__60_left_grid_pin_21_;
  wire [0:0] cby_1__1__60_left_grid_pin_22_;
  wire [0:0] cby_1__1__60_left_grid_pin_23_;
  wire [0:0] cby_1__1__60_left_grid_pin_24_;
  wire [0:0] cby_1__1__60_left_grid_pin_25_;
  wire [0:0] cby_1__1__60_left_grid_pin_26_;
  wire [0:0] cby_1__1__60_left_grid_pin_27_;
  wire [0:0] cby_1__1__60_left_grid_pin_28_;
  wire [0:0] cby_1__1__60_left_grid_pin_29_;
  wire [0:0] cby_1__1__60_left_grid_pin_30_;
  wire [0:0] cby_1__1__60_left_grid_pin_31_;
  wire [0:0] cby_1__1__61_ccff_tail;
  wire [0:29] cby_1__1__61_chany_bottom_out;
  wire [0:29] cby_1__1__61_chany_top_out;
  wire [0:0] cby_1__1__61_left_grid_pin_16_;
  wire [0:0] cby_1__1__61_left_grid_pin_17_;
  wire [0:0] cby_1__1__61_left_grid_pin_18_;
  wire [0:0] cby_1__1__61_left_grid_pin_19_;
  wire [0:0] cby_1__1__61_left_grid_pin_20_;
  wire [0:0] cby_1__1__61_left_grid_pin_21_;
  wire [0:0] cby_1__1__61_left_grid_pin_22_;
  wire [0:0] cby_1__1__61_left_grid_pin_23_;
  wire [0:0] cby_1__1__61_left_grid_pin_24_;
  wire [0:0] cby_1__1__61_left_grid_pin_25_;
  wire [0:0] cby_1__1__61_left_grid_pin_26_;
  wire [0:0] cby_1__1__61_left_grid_pin_27_;
  wire [0:0] cby_1__1__61_left_grid_pin_28_;
  wire [0:0] cby_1__1__61_left_grid_pin_29_;
  wire [0:0] cby_1__1__61_left_grid_pin_30_;
  wire [0:0] cby_1__1__61_left_grid_pin_31_;
  wire [0:0] cby_1__1__62_ccff_tail;
  wire [0:29] cby_1__1__62_chany_bottom_out;
  wire [0:29] cby_1__1__62_chany_top_out;
  wire [0:0] cby_1__1__62_left_grid_pin_16_;
  wire [0:0] cby_1__1__62_left_grid_pin_17_;
  wire [0:0] cby_1__1__62_left_grid_pin_18_;
  wire [0:0] cby_1__1__62_left_grid_pin_19_;
  wire [0:0] cby_1__1__62_left_grid_pin_20_;
  wire [0:0] cby_1__1__62_left_grid_pin_21_;
  wire [0:0] cby_1__1__62_left_grid_pin_22_;
  wire [0:0] cby_1__1__62_left_grid_pin_23_;
  wire [0:0] cby_1__1__62_left_grid_pin_24_;
  wire [0:0] cby_1__1__62_left_grid_pin_25_;
  wire [0:0] cby_1__1__62_left_grid_pin_26_;
  wire [0:0] cby_1__1__62_left_grid_pin_27_;
  wire [0:0] cby_1__1__62_left_grid_pin_28_;
  wire [0:0] cby_1__1__62_left_grid_pin_29_;
  wire [0:0] cby_1__1__62_left_grid_pin_30_;
  wire [0:0] cby_1__1__62_left_grid_pin_31_;
  wire [0:0] cby_1__1__63_ccff_tail;
  wire [0:29] cby_1__1__63_chany_bottom_out;
  wire [0:29] cby_1__1__63_chany_top_out;
  wire [0:0] cby_1__1__63_left_grid_pin_16_;
  wire [0:0] cby_1__1__63_left_grid_pin_17_;
  wire [0:0] cby_1__1__63_left_grid_pin_18_;
  wire [0:0] cby_1__1__63_left_grid_pin_19_;
  wire [0:0] cby_1__1__63_left_grid_pin_20_;
  wire [0:0] cby_1__1__63_left_grid_pin_21_;
  wire [0:0] cby_1__1__63_left_grid_pin_22_;
  wire [0:0] cby_1__1__63_left_grid_pin_23_;
  wire [0:0] cby_1__1__63_left_grid_pin_24_;
  wire [0:0] cby_1__1__63_left_grid_pin_25_;
  wire [0:0] cby_1__1__63_left_grid_pin_26_;
  wire [0:0] cby_1__1__63_left_grid_pin_27_;
  wire [0:0] cby_1__1__63_left_grid_pin_28_;
  wire [0:0] cby_1__1__63_left_grid_pin_29_;
  wire [0:0] cby_1__1__63_left_grid_pin_30_;
  wire [0:0] cby_1__1__63_left_grid_pin_31_;
  wire [0:0] cby_1__1__64_ccff_tail;
  wire [0:29] cby_1__1__64_chany_bottom_out;
  wire [0:29] cby_1__1__64_chany_top_out;
  wire [0:0] cby_1__1__64_left_grid_pin_16_;
  wire [0:0] cby_1__1__64_left_grid_pin_17_;
  wire [0:0] cby_1__1__64_left_grid_pin_18_;
  wire [0:0] cby_1__1__64_left_grid_pin_19_;
  wire [0:0] cby_1__1__64_left_grid_pin_20_;
  wire [0:0] cby_1__1__64_left_grid_pin_21_;
  wire [0:0] cby_1__1__64_left_grid_pin_22_;
  wire [0:0] cby_1__1__64_left_grid_pin_23_;
  wire [0:0] cby_1__1__64_left_grid_pin_24_;
  wire [0:0] cby_1__1__64_left_grid_pin_25_;
  wire [0:0] cby_1__1__64_left_grid_pin_26_;
  wire [0:0] cby_1__1__64_left_grid_pin_27_;
  wire [0:0] cby_1__1__64_left_grid_pin_28_;
  wire [0:0] cby_1__1__64_left_grid_pin_29_;
  wire [0:0] cby_1__1__64_left_grid_pin_30_;
  wire [0:0] cby_1__1__64_left_grid_pin_31_;
  wire [0:0] cby_1__1__65_ccff_tail;
  wire [0:29] cby_1__1__65_chany_bottom_out;
  wire [0:29] cby_1__1__65_chany_top_out;
  wire [0:0] cby_1__1__65_left_grid_pin_16_;
  wire [0:0] cby_1__1__65_left_grid_pin_17_;
  wire [0:0] cby_1__1__65_left_grid_pin_18_;
  wire [0:0] cby_1__1__65_left_grid_pin_19_;
  wire [0:0] cby_1__1__65_left_grid_pin_20_;
  wire [0:0] cby_1__1__65_left_grid_pin_21_;
  wire [0:0] cby_1__1__65_left_grid_pin_22_;
  wire [0:0] cby_1__1__65_left_grid_pin_23_;
  wire [0:0] cby_1__1__65_left_grid_pin_24_;
  wire [0:0] cby_1__1__65_left_grid_pin_25_;
  wire [0:0] cby_1__1__65_left_grid_pin_26_;
  wire [0:0] cby_1__1__65_left_grid_pin_27_;
  wire [0:0] cby_1__1__65_left_grid_pin_28_;
  wire [0:0] cby_1__1__65_left_grid_pin_29_;
  wire [0:0] cby_1__1__65_left_grid_pin_30_;
  wire [0:0] cby_1__1__65_left_grid_pin_31_;
  wire [0:0] cby_1__1__66_ccff_tail;
  wire [0:29] cby_1__1__66_chany_bottom_out;
  wire [0:29] cby_1__1__66_chany_top_out;
  wire [0:0] cby_1__1__66_left_grid_pin_16_;
  wire [0:0] cby_1__1__66_left_grid_pin_17_;
  wire [0:0] cby_1__1__66_left_grid_pin_18_;
  wire [0:0] cby_1__1__66_left_grid_pin_19_;
  wire [0:0] cby_1__1__66_left_grid_pin_20_;
  wire [0:0] cby_1__1__66_left_grid_pin_21_;
  wire [0:0] cby_1__1__66_left_grid_pin_22_;
  wire [0:0] cby_1__1__66_left_grid_pin_23_;
  wire [0:0] cby_1__1__66_left_grid_pin_24_;
  wire [0:0] cby_1__1__66_left_grid_pin_25_;
  wire [0:0] cby_1__1__66_left_grid_pin_26_;
  wire [0:0] cby_1__1__66_left_grid_pin_27_;
  wire [0:0] cby_1__1__66_left_grid_pin_28_;
  wire [0:0] cby_1__1__66_left_grid_pin_29_;
  wire [0:0] cby_1__1__66_left_grid_pin_30_;
  wire [0:0] cby_1__1__66_left_grid_pin_31_;
  wire [0:0] cby_1__1__67_ccff_tail;
  wire [0:29] cby_1__1__67_chany_bottom_out;
  wire [0:29] cby_1__1__67_chany_top_out;
  wire [0:0] cby_1__1__67_left_grid_pin_16_;
  wire [0:0] cby_1__1__67_left_grid_pin_17_;
  wire [0:0] cby_1__1__67_left_grid_pin_18_;
  wire [0:0] cby_1__1__67_left_grid_pin_19_;
  wire [0:0] cby_1__1__67_left_grid_pin_20_;
  wire [0:0] cby_1__1__67_left_grid_pin_21_;
  wire [0:0] cby_1__1__67_left_grid_pin_22_;
  wire [0:0] cby_1__1__67_left_grid_pin_23_;
  wire [0:0] cby_1__1__67_left_grid_pin_24_;
  wire [0:0] cby_1__1__67_left_grid_pin_25_;
  wire [0:0] cby_1__1__67_left_grid_pin_26_;
  wire [0:0] cby_1__1__67_left_grid_pin_27_;
  wire [0:0] cby_1__1__67_left_grid_pin_28_;
  wire [0:0] cby_1__1__67_left_grid_pin_29_;
  wire [0:0] cby_1__1__67_left_grid_pin_30_;
  wire [0:0] cby_1__1__67_left_grid_pin_31_;
  wire [0:0] cby_1__1__68_ccff_tail;
  wire [0:29] cby_1__1__68_chany_bottom_out;
  wire [0:29] cby_1__1__68_chany_top_out;
  wire [0:0] cby_1__1__68_left_grid_pin_16_;
  wire [0:0] cby_1__1__68_left_grid_pin_17_;
  wire [0:0] cby_1__1__68_left_grid_pin_18_;
  wire [0:0] cby_1__1__68_left_grid_pin_19_;
  wire [0:0] cby_1__1__68_left_grid_pin_20_;
  wire [0:0] cby_1__1__68_left_grid_pin_21_;
  wire [0:0] cby_1__1__68_left_grid_pin_22_;
  wire [0:0] cby_1__1__68_left_grid_pin_23_;
  wire [0:0] cby_1__1__68_left_grid_pin_24_;
  wire [0:0] cby_1__1__68_left_grid_pin_25_;
  wire [0:0] cby_1__1__68_left_grid_pin_26_;
  wire [0:0] cby_1__1__68_left_grid_pin_27_;
  wire [0:0] cby_1__1__68_left_grid_pin_28_;
  wire [0:0] cby_1__1__68_left_grid_pin_29_;
  wire [0:0] cby_1__1__68_left_grid_pin_30_;
  wire [0:0] cby_1__1__68_left_grid_pin_31_;
  wire [0:0] cby_1__1__69_ccff_tail;
  wire [0:29] cby_1__1__69_chany_bottom_out;
  wire [0:29] cby_1__1__69_chany_top_out;
  wire [0:0] cby_1__1__69_left_grid_pin_16_;
  wire [0:0] cby_1__1__69_left_grid_pin_17_;
  wire [0:0] cby_1__1__69_left_grid_pin_18_;
  wire [0:0] cby_1__1__69_left_grid_pin_19_;
  wire [0:0] cby_1__1__69_left_grid_pin_20_;
  wire [0:0] cby_1__1__69_left_grid_pin_21_;
  wire [0:0] cby_1__1__69_left_grid_pin_22_;
  wire [0:0] cby_1__1__69_left_grid_pin_23_;
  wire [0:0] cby_1__1__69_left_grid_pin_24_;
  wire [0:0] cby_1__1__69_left_grid_pin_25_;
  wire [0:0] cby_1__1__69_left_grid_pin_26_;
  wire [0:0] cby_1__1__69_left_grid_pin_27_;
  wire [0:0] cby_1__1__69_left_grid_pin_28_;
  wire [0:0] cby_1__1__69_left_grid_pin_29_;
  wire [0:0] cby_1__1__69_left_grid_pin_30_;
  wire [0:0] cby_1__1__69_left_grid_pin_31_;
  wire [0:0] cby_1__1__6_ccff_tail;
  wire [0:29] cby_1__1__6_chany_bottom_out;
  wire [0:29] cby_1__1__6_chany_top_out;
  wire [0:0] cby_1__1__6_left_grid_pin_16_;
  wire [0:0] cby_1__1__6_left_grid_pin_17_;
  wire [0:0] cby_1__1__6_left_grid_pin_18_;
  wire [0:0] cby_1__1__6_left_grid_pin_19_;
  wire [0:0] cby_1__1__6_left_grid_pin_20_;
  wire [0:0] cby_1__1__6_left_grid_pin_21_;
  wire [0:0] cby_1__1__6_left_grid_pin_22_;
  wire [0:0] cby_1__1__6_left_grid_pin_23_;
  wire [0:0] cby_1__1__6_left_grid_pin_24_;
  wire [0:0] cby_1__1__6_left_grid_pin_25_;
  wire [0:0] cby_1__1__6_left_grid_pin_26_;
  wire [0:0] cby_1__1__6_left_grid_pin_27_;
  wire [0:0] cby_1__1__6_left_grid_pin_28_;
  wire [0:0] cby_1__1__6_left_grid_pin_29_;
  wire [0:0] cby_1__1__6_left_grid_pin_30_;
  wire [0:0] cby_1__1__6_left_grid_pin_31_;
  wire [0:0] cby_1__1__70_ccff_tail;
  wire [0:29] cby_1__1__70_chany_bottom_out;
  wire [0:29] cby_1__1__70_chany_top_out;
  wire [0:0] cby_1__1__70_left_grid_pin_16_;
  wire [0:0] cby_1__1__70_left_grid_pin_17_;
  wire [0:0] cby_1__1__70_left_grid_pin_18_;
  wire [0:0] cby_1__1__70_left_grid_pin_19_;
  wire [0:0] cby_1__1__70_left_grid_pin_20_;
  wire [0:0] cby_1__1__70_left_grid_pin_21_;
  wire [0:0] cby_1__1__70_left_grid_pin_22_;
  wire [0:0] cby_1__1__70_left_grid_pin_23_;
  wire [0:0] cby_1__1__70_left_grid_pin_24_;
  wire [0:0] cby_1__1__70_left_grid_pin_25_;
  wire [0:0] cby_1__1__70_left_grid_pin_26_;
  wire [0:0] cby_1__1__70_left_grid_pin_27_;
  wire [0:0] cby_1__1__70_left_grid_pin_28_;
  wire [0:0] cby_1__1__70_left_grid_pin_29_;
  wire [0:0] cby_1__1__70_left_grid_pin_30_;
  wire [0:0] cby_1__1__70_left_grid_pin_31_;
  wire [0:0] cby_1__1__71_ccff_tail;
  wire [0:29] cby_1__1__71_chany_bottom_out;
  wire [0:29] cby_1__1__71_chany_top_out;
  wire [0:0] cby_1__1__71_left_grid_pin_16_;
  wire [0:0] cby_1__1__71_left_grid_pin_17_;
  wire [0:0] cby_1__1__71_left_grid_pin_18_;
  wire [0:0] cby_1__1__71_left_grid_pin_19_;
  wire [0:0] cby_1__1__71_left_grid_pin_20_;
  wire [0:0] cby_1__1__71_left_grid_pin_21_;
  wire [0:0] cby_1__1__71_left_grid_pin_22_;
  wire [0:0] cby_1__1__71_left_grid_pin_23_;
  wire [0:0] cby_1__1__71_left_grid_pin_24_;
  wire [0:0] cby_1__1__71_left_grid_pin_25_;
  wire [0:0] cby_1__1__71_left_grid_pin_26_;
  wire [0:0] cby_1__1__71_left_grid_pin_27_;
  wire [0:0] cby_1__1__71_left_grid_pin_28_;
  wire [0:0] cby_1__1__71_left_grid_pin_29_;
  wire [0:0] cby_1__1__71_left_grid_pin_30_;
  wire [0:0] cby_1__1__71_left_grid_pin_31_;
  wire [0:0] cby_1__1__72_ccff_tail;
  wire [0:29] cby_1__1__72_chany_bottom_out;
  wire [0:29] cby_1__1__72_chany_top_out;
  wire [0:0] cby_1__1__72_left_grid_pin_16_;
  wire [0:0] cby_1__1__72_left_grid_pin_17_;
  wire [0:0] cby_1__1__72_left_grid_pin_18_;
  wire [0:0] cby_1__1__72_left_grid_pin_19_;
  wire [0:0] cby_1__1__72_left_grid_pin_20_;
  wire [0:0] cby_1__1__72_left_grid_pin_21_;
  wire [0:0] cby_1__1__72_left_grid_pin_22_;
  wire [0:0] cby_1__1__72_left_grid_pin_23_;
  wire [0:0] cby_1__1__72_left_grid_pin_24_;
  wire [0:0] cby_1__1__72_left_grid_pin_25_;
  wire [0:0] cby_1__1__72_left_grid_pin_26_;
  wire [0:0] cby_1__1__72_left_grid_pin_27_;
  wire [0:0] cby_1__1__72_left_grid_pin_28_;
  wire [0:0] cby_1__1__72_left_grid_pin_29_;
  wire [0:0] cby_1__1__72_left_grid_pin_30_;
  wire [0:0] cby_1__1__72_left_grid_pin_31_;
  wire [0:0] cby_1__1__73_ccff_tail;
  wire [0:29] cby_1__1__73_chany_bottom_out;
  wire [0:29] cby_1__1__73_chany_top_out;
  wire [0:0] cby_1__1__73_left_grid_pin_16_;
  wire [0:0] cby_1__1__73_left_grid_pin_17_;
  wire [0:0] cby_1__1__73_left_grid_pin_18_;
  wire [0:0] cby_1__1__73_left_grid_pin_19_;
  wire [0:0] cby_1__1__73_left_grid_pin_20_;
  wire [0:0] cby_1__1__73_left_grid_pin_21_;
  wire [0:0] cby_1__1__73_left_grid_pin_22_;
  wire [0:0] cby_1__1__73_left_grid_pin_23_;
  wire [0:0] cby_1__1__73_left_grid_pin_24_;
  wire [0:0] cby_1__1__73_left_grid_pin_25_;
  wire [0:0] cby_1__1__73_left_grid_pin_26_;
  wire [0:0] cby_1__1__73_left_grid_pin_27_;
  wire [0:0] cby_1__1__73_left_grid_pin_28_;
  wire [0:0] cby_1__1__73_left_grid_pin_29_;
  wire [0:0] cby_1__1__73_left_grid_pin_30_;
  wire [0:0] cby_1__1__73_left_grid_pin_31_;
  wire [0:0] cby_1__1__74_ccff_tail;
  wire [0:29] cby_1__1__74_chany_bottom_out;
  wire [0:29] cby_1__1__74_chany_top_out;
  wire [0:0] cby_1__1__74_left_grid_pin_16_;
  wire [0:0] cby_1__1__74_left_grid_pin_17_;
  wire [0:0] cby_1__1__74_left_grid_pin_18_;
  wire [0:0] cby_1__1__74_left_grid_pin_19_;
  wire [0:0] cby_1__1__74_left_grid_pin_20_;
  wire [0:0] cby_1__1__74_left_grid_pin_21_;
  wire [0:0] cby_1__1__74_left_grid_pin_22_;
  wire [0:0] cby_1__1__74_left_grid_pin_23_;
  wire [0:0] cby_1__1__74_left_grid_pin_24_;
  wire [0:0] cby_1__1__74_left_grid_pin_25_;
  wire [0:0] cby_1__1__74_left_grid_pin_26_;
  wire [0:0] cby_1__1__74_left_grid_pin_27_;
  wire [0:0] cby_1__1__74_left_grid_pin_28_;
  wire [0:0] cby_1__1__74_left_grid_pin_29_;
  wire [0:0] cby_1__1__74_left_grid_pin_30_;
  wire [0:0] cby_1__1__74_left_grid_pin_31_;
  wire [0:0] cby_1__1__75_ccff_tail;
  wire [0:29] cby_1__1__75_chany_bottom_out;
  wire [0:29] cby_1__1__75_chany_top_out;
  wire [0:0] cby_1__1__75_left_grid_pin_16_;
  wire [0:0] cby_1__1__75_left_grid_pin_17_;
  wire [0:0] cby_1__1__75_left_grid_pin_18_;
  wire [0:0] cby_1__1__75_left_grid_pin_19_;
  wire [0:0] cby_1__1__75_left_grid_pin_20_;
  wire [0:0] cby_1__1__75_left_grid_pin_21_;
  wire [0:0] cby_1__1__75_left_grid_pin_22_;
  wire [0:0] cby_1__1__75_left_grid_pin_23_;
  wire [0:0] cby_1__1__75_left_grid_pin_24_;
  wire [0:0] cby_1__1__75_left_grid_pin_25_;
  wire [0:0] cby_1__1__75_left_grid_pin_26_;
  wire [0:0] cby_1__1__75_left_grid_pin_27_;
  wire [0:0] cby_1__1__75_left_grid_pin_28_;
  wire [0:0] cby_1__1__75_left_grid_pin_29_;
  wire [0:0] cby_1__1__75_left_grid_pin_30_;
  wire [0:0] cby_1__1__75_left_grid_pin_31_;
  wire [0:0] cby_1__1__76_ccff_tail;
  wire [0:29] cby_1__1__76_chany_bottom_out;
  wire [0:29] cby_1__1__76_chany_top_out;
  wire [0:0] cby_1__1__76_left_grid_pin_16_;
  wire [0:0] cby_1__1__76_left_grid_pin_17_;
  wire [0:0] cby_1__1__76_left_grid_pin_18_;
  wire [0:0] cby_1__1__76_left_grid_pin_19_;
  wire [0:0] cby_1__1__76_left_grid_pin_20_;
  wire [0:0] cby_1__1__76_left_grid_pin_21_;
  wire [0:0] cby_1__1__76_left_grid_pin_22_;
  wire [0:0] cby_1__1__76_left_grid_pin_23_;
  wire [0:0] cby_1__1__76_left_grid_pin_24_;
  wire [0:0] cby_1__1__76_left_grid_pin_25_;
  wire [0:0] cby_1__1__76_left_grid_pin_26_;
  wire [0:0] cby_1__1__76_left_grid_pin_27_;
  wire [0:0] cby_1__1__76_left_grid_pin_28_;
  wire [0:0] cby_1__1__76_left_grid_pin_29_;
  wire [0:0] cby_1__1__76_left_grid_pin_30_;
  wire [0:0] cby_1__1__76_left_grid_pin_31_;
  wire [0:0] cby_1__1__77_ccff_tail;
  wire [0:29] cby_1__1__77_chany_bottom_out;
  wire [0:29] cby_1__1__77_chany_top_out;
  wire [0:0] cby_1__1__77_left_grid_pin_16_;
  wire [0:0] cby_1__1__77_left_grid_pin_17_;
  wire [0:0] cby_1__1__77_left_grid_pin_18_;
  wire [0:0] cby_1__1__77_left_grid_pin_19_;
  wire [0:0] cby_1__1__77_left_grid_pin_20_;
  wire [0:0] cby_1__1__77_left_grid_pin_21_;
  wire [0:0] cby_1__1__77_left_grid_pin_22_;
  wire [0:0] cby_1__1__77_left_grid_pin_23_;
  wire [0:0] cby_1__1__77_left_grid_pin_24_;
  wire [0:0] cby_1__1__77_left_grid_pin_25_;
  wire [0:0] cby_1__1__77_left_grid_pin_26_;
  wire [0:0] cby_1__1__77_left_grid_pin_27_;
  wire [0:0] cby_1__1__77_left_grid_pin_28_;
  wire [0:0] cby_1__1__77_left_grid_pin_29_;
  wire [0:0] cby_1__1__77_left_grid_pin_30_;
  wire [0:0] cby_1__1__77_left_grid_pin_31_;
  wire [0:0] cby_1__1__78_ccff_tail;
  wire [0:29] cby_1__1__78_chany_bottom_out;
  wire [0:29] cby_1__1__78_chany_top_out;
  wire [0:0] cby_1__1__78_left_grid_pin_16_;
  wire [0:0] cby_1__1__78_left_grid_pin_17_;
  wire [0:0] cby_1__1__78_left_grid_pin_18_;
  wire [0:0] cby_1__1__78_left_grid_pin_19_;
  wire [0:0] cby_1__1__78_left_grid_pin_20_;
  wire [0:0] cby_1__1__78_left_grid_pin_21_;
  wire [0:0] cby_1__1__78_left_grid_pin_22_;
  wire [0:0] cby_1__1__78_left_grid_pin_23_;
  wire [0:0] cby_1__1__78_left_grid_pin_24_;
  wire [0:0] cby_1__1__78_left_grid_pin_25_;
  wire [0:0] cby_1__1__78_left_grid_pin_26_;
  wire [0:0] cby_1__1__78_left_grid_pin_27_;
  wire [0:0] cby_1__1__78_left_grid_pin_28_;
  wire [0:0] cby_1__1__78_left_grid_pin_29_;
  wire [0:0] cby_1__1__78_left_grid_pin_30_;
  wire [0:0] cby_1__1__78_left_grid_pin_31_;
  wire [0:0] cby_1__1__79_ccff_tail;
  wire [0:29] cby_1__1__79_chany_bottom_out;
  wire [0:29] cby_1__1__79_chany_top_out;
  wire [0:0] cby_1__1__79_left_grid_pin_16_;
  wire [0:0] cby_1__1__79_left_grid_pin_17_;
  wire [0:0] cby_1__1__79_left_grid_pin_18_;
  wire [0:0] cby_1__1__79_left_grid_pin_19_;
  wire [0:0] cby_1__1__79_left_grid_pin_20_;
  wire [0:0] cby_1__1__79_left_grid_pin_21_;
  wire [0:0] cby_1__1__79_left_grid_pin_22_;
  wire [0:0] cby_1__1__79_left_grid_pin_23_;
  wire [0:0] cby_1__1__79_left_grid_pin_24_;
  wire [0:0] cby_1__1__79_left_grid_pin_25_;
  wire [0:0] cby_1__1__79_left_grid_pin_26_;
  wire [0:0] cby_1__1__79_left_grid_pin_27_;
  wire [0:0] cby_1__1__79_left_grid_pin_28_;
  wire [0:0] cby_1__1__79_left_grid_pin_29_;
  wire [0:0] cby_1__1__79_left_grid_pin_30_;
  wire [0:0] cby_1__1__79_left_grid_pin_31_;
  wire [0:0] cby_1__1__7_ccff_tail;
  wire [0:29] cby_1__1__7_chany_bottom_out;
  wire [0:29] cby_1__1__7_chany_top_out;
  wire [0:0] cby_1__1__7_left_grid_pin_16_;
  wire [0:0] cby_1__1__7_left_grid_pin_17_;
  wire [0:0] cby_1__1__7_left_grid_pin_18_;
  wire [0:0] cby_1__1__7_left_grid_pin_19_;
  wire [0:0] cby_1__1__7_left_grid_pin_20_;
  wire [0:0] cby_1__1__7_left_grid_pin_21_;
  wire [0:0] cby_1__1__7_left_grid_pin_22_;
  wire [0:0] cby_1__1__7_left_grid_pin_23_;
  wire [0:0] cby_1__1__7_left_grid_pin_24_;
  wire [0:0] cby_1__1__7_left_grid_pin_25_;
  wire [0:0] cby_1__1__7_left_grid_pin_26_;
  wire [0:0] cby_1__1__7_left_grid_pin_27_;
  wire [0:0] cby_1__1__7_left_grid_pin_28_;
  wire [0:0] cby_1__1__7_left_grid_pin_29_;
  wire [0:0] cby_1__1__7_left_grid_pin_30_;
  wire [0:0] cby_1__1__7_left_grid_pin_31_;
  wire [0:0] cby_1__1__80_ccff_tail;
  wire [0:29] cby_1__1__80_chany_bottom_out;
  wire [0:29] cby_1__1__80_chany_top_out;
  wire [0:0] cby_1__1__80_left_grid_pin_16_;
  wire [0:0] cby_1__1__80_left_grid_pin_17_;
  wire [0:0] cby_1__1__80_left_grid_pin_18_;
  wire [0:0] cby_1__1__80_left_grid_pin_19_;
  wire [0:0] cby_1__1__80_left_grid_pin_20_;
  wire [0:0] cby_1__1__80_left_grid_pin_21_;
  wire [0:0] cby_1__1__80_left_grid_pin_22_;
  wire [0:0] cby_1__1__80_left_grid_pin_23_;
  wire [0:0] cby_1__1__80_left_grid_pin_24_;
  wire [0:0] cby_1__1__80_left_grid_pin_25_;
  wire [0:0] cby_1__1__80_left_grid_pin_26_;
  wire [0:0] cby_1__1__80_left_grid_pin_27_;
  wire [0:0] cby_1__1__80_left_grid_pin_28_;
  wire [0:0] cby_1__1__80_left_grid_pin_29_;
  wire [0:0] cby_1__1__80_left_grid_pin_30_;
  wire [0:0] cby_1__1__80_left_grid_pin_31_;
  wire [0:0] cby_1__1__81_ccff_tail;
  wire [0:29] cby_1__1__81_chany_bottom_out;
  wire [0:29] cby_1__1__81_chany_top_out;
  wire [0:0] cby_1__1__81_left_grid_pin_16_;
  wire [0:0] cby_1__1__81_left_grid_pin_17_;
  wire [0:0] cby_1__1__81_left_grid_pin_18_;
  wire [0:0] cby_1__1__81_left_grid_pin_19_;
  wire [0:0] cby_1__1__81_left_grid_pin_20_;
  wire [0:0] cby_1__1__81_left_grid_pin_21_;
  wire [0:0] cby_1__1__81_left_grid_pin_22_;
  wire [0:0] cby_1__1__81_left_grid_pin_23_;
  wire [0:0] cby_1__1__81_left_grid_pin_24_;
  wire [0:0] cby_1__1__81_left_grid_pin_25_;
  wire [0:0] cby_1__1__81_left_grid_pin_26_;
  wire [0:0] cby_1__1__81_left_grid_pin_27_;
  wire [0:0] cby_1__1__81_left_grid_pin_28_;
  wire [0:0] cby_1__1__81_left_grid_pin_29_;
  wire [0:0] cby_1__1__81_left_grid_pin_30_;
  wire [0:0] cby_1__1__81_left_grid_pin_31_;
  wire [0:0] cby_1__1__82_ccff_tail;
  wire [0:29] cby_1__1__82_chany_bottom_out;
  wire [0:29] cby_1__1__82_chany_top_out;
  wire [0:0] cby_1__1__82_left_grid_pin_16_;
  wire [0:0] cby_1__1__82_left_grid_pin_17_;
  wire [0:0] cby_1__1__82_left_grid_pin_18_;
  wire [0:0] cby_1__1__82_left_grid_pin_19_;
  wire [0:0] cby_1__1__82_left_grid_pin_20_;
  wire [0:0] cby_1__1__82_left_grid_pin_21_;
  wire [0:0] cby_1__1__82_left_grid_pin_22_;
  wire [0:0] cby_1__1__82_left_grid_pin_23_;
  wire [0:0] cby_1__1__82_left_grid_pin_24_;
  wire [0:0] cby_1__1__82_left_grid_pin_25_;
  wire [0:0] cby_1__1__82_left_grid_pin_26_;
  wire [0:0] cby_1__1__82_left_grid_pin_27_;
  wire [0:0] cby_1__1__82_left_grid_pin_28_;
  wire [0:0] cby_1__1__82_left_grid_pin_29_;
  wire [0:0] cby_1__1__82_left_grid_pin_30_;
  wire [0:0] cby_1__1__82_left_grid_pin_31_;
  wire [0:0] cby_1__1__83_ccff_tail;
  wire [0:29] cby_1__1__83_chany_bottom_out;
  wire [0:29] cby_1__1__83_chany_top_out;
  wire [0:0] cby_1__1__83_left_grid_pin_16_;
  wire [0:0] cby_1__1__83_left_grid_pin_17_;
  wire [0:0] cby_1__1__83_left_grid_pin_18_;
  wire [0:0] cby_1__1__83_left_grid_pin_19_;
  wire [0:0] cby_1__1__83_left_grid_pin_20_;
  wire [0:0] cby_1__1__83_left_grid_pin_21_;
  wire [0:0] cby_1__1__83_left_grid_pin_22_;
  wire [0:0] cby_1__1__83_left_grid_pin_23_;
  wire [0:0] cby_1__1__83_left_grid_pin_24_;
  wire [0:0] cby_1__1__83_left_grid_pin_25_;
  wire [0:0] cby_1__1__83_left_grid_pin_26_;
  wire [0:0] cby_1__1__83_left_grid_pin_27_;
  wire [0:0] cby_1__1__83_left_grid_pin_28_;
  wire [0:0] cby_1__1__83_left_grid_pin_29_;
  wire [0:0] cby_1__1__83_left_grid_pin_30_;
  wire [0:0] cby_1__1__83_left_grid_pin_31_;
  wire [0:0] cby_1__1__84_ccff_tail;
  wire [0:29] cby_1__1__84_chany_bottom_out;
  wire [0:29] cby_1__1__84_chany_top_out;
  wire [0:0] cby_1__1__84_left_grid_pin_16_;
  wire [0:0] cby_1__1__84_left_grid_pin_17_;
  wire [0:0] cby_1__1__84_left_grid_pin_18_;
  wire [0:0] cby_1__1__84_left_grid_pin_19_;
  wire [0:0] cby_1__1__84_left_grid_pin_20_;
  wire [0:0] cby_1__1__84_left_grid_pin_21_;
  wire [0:0] cby_1__1__84_left_grid_pin_22_;
  wire [0:0] cby_1__1__84_left_grid_pin_23_;
  wire [0:0] cby_1__1__84_left_grid_pin_24_;
  wire [0:0] cby_1__1__84_left_grid_pin_25_;
  wire [0:0] cby_1__1__84_left_grid_pin_26_;
  wire [0:0] cby_1__1__84_left_grid_pin_27_;
  wire [0:0] cby_1__1__84_left_grid_pin_28_;
  wire [0:0] cby_1__1__84_left_grid_pin_29_;
  wire [0:0] cby_1__1__84_left_grid_pin_30_;
  wire [0:0] cby_1__1__84_left_grid_pin_31_;
  wire [0:0] cby_1__1__85_ccff_tail;
  wire [0:29] cby_1__1__85_chany_bottom_out;
  wire [0:29] cby_1__1__85_chany_top_out;
  wire [0:0] cby_1__1__85_left_grid_pin_16_;
  wire [0:0] cby_1__1__85_left_grid_pin_17_;
  wire [0:0] cby_1__1__85_left_grid_pin_18_;
  wire [0:0] cby_1__1__85_left_grid_pin_19_;
  wire [0:0] cby_1__1__85_left_grid_pin_20_;
  wire [0:0] cby_1__1__85_left_grid_pin_21_;
  wire [0:0] cby_1__1__85_left_grid_pin_22_;
  wire [0:0] cby_1__1__85_left_grid_pin_23_;
  wire [0:0] cby_1__1__85_left_grid_pin_24_;
  wire [0:0] cby_1__1__85_left_grid_pin_25_;
  wire [0:0] cby_1__1__85_left_grid_pin_26_;
  wire [0:0] cby_1__1__85_left_grid_pin_27_;
  wire [0:0] cby_1__1__85_left_grid_pin_28_;
  wire [0:0] cby_1__1__85_left_grid_pin_29_;
  wire [0:0] cby_1__1__85_left_grid_pin_30_;
  wire [0:0] cby_1__1__85_left_grid_pin_31_;
  wire [0:0] cby_1__1__86_ccff_tail;
  wire [0:29] cby_1__1__86_chany_bottom_out;
  wire [0:29] cby_1__1__86_chany_top_out;
  wire [0:0] cby_1__1__86_left_grid_pin_16_;
  wire [0:0] cby_1__1__86_left_grid_pin_17_;
  wire [0:0] cby_1__1__86_left_grid_pin_18_;
  wire [0:0] cby_1__1__86_left_grid_pin_19_;
  wire [0:0] cby_1__1__86_left_grid_pin_20_;
  wire [0:0] cby_1__1__86_left_grid_pin_21_;
  wire [0:0] cby_1__1__86_left_grid_pin_22_;
  wire [0:0] cby_1__1__86_left_grid_pin_23_;
  wire [0:0] cby_1__1__86_left_grid_pin_24_;
  wire [0:0] cby_1__1__86_left_grid_pin_25_;
  wire [0:0] cby_1__1__86_left_grid_pin_26_;
  wire [0:0] cby_1__1__86_left_grid_pin_27_;
  wire [0:0] cby_1__1__86_left_grid_pin_28_;
  wire [0:0] cby_1__1__86_left_grid_pin_29_;
  wire [0:0] cby_1__1__86_left_grid_pin_30_;
  wire [0:0] cby_1__1__86_left_grid_pin_31_;
  wire [0:0] cby_1__1__87_ccff_tail;
  wire [0:29] cby_1__1__87_chany_bottom_out;
  wire [0:29] cby_1__1__87_chany_top_out;
  wire [0:0] cby_1__1__87_left_grid_pin_16_;
  wire [0:0] cby_1__1__87_left_grid_pin_17_;
  wire [0:0] cby_1__1__87_left_grid_pin_18_;
  wire [0:0] cby_1__1__87_left_grid_pin_19_;
  wire [0:0] cby_1__1__87_left_grid_pin_20_;
  wire [0:0] cby_1__1__87_left_grid_pin_21_;
  wire [0:0] cby_1__1__87_left_grid_pin_22_;
  wire [0:0] cby_1__1__87_left_grid_pin_23_;
  wire [0:0] cby_1__1__87_left_grid_pin_24_;
  wire [0:0] cby_1__1__87_left_grid_pin_25_;
  wire [0:0] cby_1__1__87_left_grid_pin_26_;
  wire [0:0] cby_1__1__87_left_grid_pin_27_;
  wire [0:0] cby_1__1__87_left_grid_pin_28_;
  wire [0:0] cby_1__1__87_left_grid_pin_29_;
  wire [0:0] cby_1__1__87_left_grid_pin_30_;
  wire [0:0] cby_1__1__87_left_grid_pin_31_;
  wire [0:0] cby_1__1__88_ccff_tail;
  wire [0:29] cby_1__1__88_chany_bottom_out;
  wire [0:29] cby_1__1__88_chany_top_out;
  wire [0:0] cby_1__1__88_left_grid_pin_16_;
  wire [0:0] cby_1__1__88_left_grid_pin_17_;
  wire [0:0] cby_1__1__88_left_grid_pin_18_;
  wire [0:0] cby_1__1__88_left_grid_pin_19_;
  wire [0:0] cby_1__1__88_left_grid_pin_20_;
  wire [0:0] cby_1__1__88_left_grid_pin_21_;
  wire [0:0] cby_1__1__88_left_grid_pin_22_;
  wire [0:0] cby_1__1__88_left_grid_pin_23_;
  wire [0:0] cby_1__1__88_left_grid_pin_24_;
  wire [0:0] cby_1__1__88_left_grid_pin_25_;
  wire [0:0] cby_1__1__88_left_grid_pin_26_;
  wire [0:0] cby_1__1__88_left_grid_pin_27_;
  wire [0:0] cby_1__1__88_left_grid_pin_28_;
  wire [0:0] cby_1__1__88_left_grid_pin_29_;
  wire [0:0] cby_1__1__88_left_grid_pin_30_;
  wire [0:0] cby_1__1__88_left_grid_pin_31_;
  wire [0:0] cby_1__1__89_ccff_tail;
  wire [0:29] cby_1__1__89_chany_bottom_out;
  wire [0:29] cby_1__1__89_chany_top_out;
  wire [0:0] cby_1__1__89_left_grid_pin_16_;
  wire [0:0] cby_1__1__89_left_grid_pin_17_;
  wire [0:0] cby_1__1__89_left_grid_pin_18_;
  wire [0:0] cby_1__1__89_left_grid_pin_19_;
  wire [0:0] cby_1__1__89_left_grid_pin_20_;
  wire [0:0] cby_1__1__89_left_grid_pin_21_;
  wire [0:0] cby_1__1__89_left_grid_pin_22_;
  wire [0:0] cby_1__1__89_left_grid_pin_23_;
  wire [0:0] cby_1__1__89_left_grid_pin_24_;
  wire [0:0] cby_1__1__89_left_grid_pin_25_;
  wire [0:0] cby_1__1__89_left_grid_pin_26_;
  wire [0:0] cby_1__1__89_left_grid_pin_27_;
  wire [0:0] cby_1__1__89_left_grid_pin_28_;
  wire [0:0] cby_1__1__89_left_grid_pin_29_;
  wire [0:0] cby_1__1__89_left_grid_pin_30_;
  wire [0:0] cby_1__1__89_left_grid_pin_31_;
  wire [0:0] cby_1__1__8_ccff_tail;
  wire [0:29] cby_1__1__8_chany_bottom_out;
  wire [0:29] cby_1__1__8_chany_top_out;
  wire [0:0] cby_1__1__8_left_grid_pin_16_;
  wire [0:0] cby_1__1__8_left_grid_pin_17_;
  wire [0:0] cby_1__1__8_left_grid_pin_18_;
  wire [0:0] cby_1__1__8_left_grid_pin_19_;
  wire [0:0] cby_1__1__8_left_grid_pin_20_;
  wire [0:0] cby_1__1__8_left_grid_pin_21_;
  wire [0:0] cby_1__1__8_left_grid_pin_22_;
  wire [0:0] cby_1__1__8_left_grid_pin_23_;
  wire [0:0] cby_1__1__8_left_grid_pin_24_;
  wire [0:0] cby_1__1__8_left_grid_pin_25_;
  wire [0:0] cby_1__1__8_left_grid_pin_26_;
  wire [0:0] cby_1__1__8_left_grid_pin_27_;
  wire [0:0] cby_1__1__8_left_grid_pin_28_;
  wire [0:0] cby_1__1__8_left_grid_pin_29_;
  wire [0:0] cby_1__1__8_left_grid_pin_30_;
  wire [0:0] cby_1__1__8_left_grid_pin_31_;
  wire [0:0] cby_1__1__90_ccff_tail;
  wire [0:29] cby_1__1__90_chany_bottom_out;
  wire [0:29] cby_1__1__90_chany_top_out;
  wire [0:0] cby_1__1__90_left_grid_pin_16_;
  wire [0:0] cby_1__1__90_left_grid_pin_17_;
  wire [0:0] cby_1__1__90_left_grid_pin_18_;
  wire [0:0] cby_1__1__90_left_grid_pin_19_;
  wire [0:0] cby_1__1__90_left_grid_pin_20_;
  wire [0:0] cby_1__1__90_left_grid_pin_21_;
  wire [0:0] cby_1__1__90_left_grid_pin_22_;
  wire [0:0] cby_1__1__90_left_grid_pin_23_;
  wire [0:0] cby_1__1__90_left_grid_pin_24_;
  wire [0:0] cby_1__1__90_left_grid_pin_25_;
  wire [0:0] cby_1__1__90_left_grid_pin_26_;
  wire [0:0] cby_1__1__90_left_grid_pin_27_;
  wire [0:0] cby_1__1__90_left_grid_pin_28_;
  wire [0:0] cby_1__1__90_left_grid_pin_29_;
  wire [0:0] cby_1__1__90_left_grid_pin_30_;
  wire [0:0] cby_1__1__90_left_grid_pin_31_;
  wire [0:0] cby_1__1__91_ccff_tail;
  wire [0:29] cby_1__1__91_chany_bottom_out;
  wire [0:29] cby_1__1__91_chany_top_out;
  wire [0:0] cby_1__1__91_left_grid_pin_16_;
  wire [0:0] cby_1__1__91_left_grid_pin_17_;
  wire [0:0] cby_1__1__91_left_grid_pin_18_;
  wire [0:0] cby_1__1__91_left_grid_pin_19_;
  wire [0:0] cby_1__1__91_left_grid_pin_20_;
  wire [0:0] cby_1__1__91_left_grid_pin_21_;
  wire [0:0] cby_1__1__91_left_grid_pin_22_;
  wire [0:0] cby_1__1__91_left_grid_pin_23_;
  wire [0:0] cby_1__1__91_left_grid_pin_24_;
  wire [0:0] cby_1__1__91_left_grid_pin_25_;
  wire [0:0] cby_1__1__91_left_grid_pin_26_;
  wire [0:0] cby_1__1__91_left_grid_pin_27_;
  wire [0:0] cby_1__1__91_left_grid_pin_28_;
  wire [0:0] cby_1__1__91_left_grid_pin_29_;
  wire [0:0] cby_1__1__91_left_grid_pin_30_;
  wire [0:0] cby_1__1__91_left_grid_pin_31_;
  wire [0:0] cby_1__1__92_ccff_tail;
  wire [0:29] cby_1__1__92_chany_bottom_out;
  wire [0:29] cby_1__1__92_chany_top_out;
  wire [0:0] cby_1__1__92_left_grid_pin_16_;
  wire [0:0] cby_1__1__92_left_grid_pin_17_;
  wire [0:0] cby_1__1__92_left_grid_pin_18_;
  wire [0:0] cby_1__1__92_left_grid_pin_19_;
  wire [0:0] cby_1__1__92_left_grid_pin_20_;
  wire [0:0] cby_1__1__92_left_grid_pin_21_;
  wire [0:0] cby_1__1__92_left_grid_pin_22_;
  wire [0:0] cby_1__1__92_left_grid_pin_23_;
  wire [0:0] cby_1__1__92_left_grid_pin_24_;
  wire [0:0] cby_1__1__92_left_grid_pin_25_;
  wire [0:0] cby_1__1__92_left_grid_pin_26_;
  wire [0:0] cby_1__1__92_left_grid_pin_27_;
  wire [0:0] cby_1__1__92_left_grid_pin_28_;
  wire [0:0] cby_1__1__92_left_grid_pin_29_;
  wire [0:0] cby_1__1__92_left_grid_pin_30_;
  wire [0:0] cby_1__1__92_left_grid_pin_31_;
  wire [0:0] cby_1__1__93_ccff_tail;
  wire [0:29] cby_1__1__93_chany_bottom_out;
  wire [0:29] cby_1__1__93_chany_top_out;
  wire [0:0] cby_1__1__93_left_grid_pin_16_;
  wire [0:0] cby_1__1__93_left_grid_pin_17_;
  wire [0:0] cby_1__1__93_left_grid_pin_18_;
  wire [0:0] cby_1__1__93_left_grid_pin_19_;
  wire [0:0] cby_1__1__93_left_grid_pin_20_;
  wire [0:0] cby_1__1__93_left_grid_pin_21_;
  wire [0:0] cby_1__1__93_left_grid_pin_22_;
  wire [0:0] cby_1__1__93_left_grid_pin_23_;
  wire [0:0] cby_1__1__93_left_grid_pin_24_;
  wire [0:0] cby_1__1__93_left_grid_pin_25_;
  wire [0:0] cby_1__1__93_left_grid_pin_26_;
  wire [0:0] cby_1__1__93_left_grid_pin_27_;
  wire [0:0] cby_1__1__93_left_grid_pin_28_;
  wire [0:0] cby_1__1__93_left_grid_pin_29_;
  wire [0:0] cby_1__1__93_left_grid_pin_30_;
  wire [0:0] cby_1__1__93_left_grid_pin_31_;
  wire [0:0] cby_1__1__94_ccff_tail;
  wire [0:29] cby_1__1__94_chany_bottom_out;
  wire [0:29] cby_1__1__94_chany_top_out;
  wire [0:0] cby_1__1__94_left_grid_pin_16_;
  wire [0:0] cby_1__1__94_left_grid_pin_17_;
  wire [0:0] cby_1__1__94_left_grid_pin_18_;
  wire [0:0] cby_1__1__94_left_grid_pin_19_;
  wire [0:0] cby_1__1__94_left_grid_pin_20_;
  wire [0:0] cby_1__1__94_left_grid_pin_21_;
  wire [0:0] cby_1__1__94_left_grid_pin_22_;
  wire [0:0] cby_1__1__94_left_grid_pin_23_;
  wire [0:0] cby_1__1__94_left_grid_pin_24_;
  wire [0:0] cby_1__1__94_left_grid_pin_25_;
  wire [0:0] cby_1__1__94_left_grid_pin_26_;
  wire [0:0] cby_1__1__94_left_grid_pin_27_;
  wire [0:0] cby_1__1__94_left_grid_pin_28_;
  wire [0:0] cby_1__1__94_left_grid_pin_29_;
  wire [0:0] cby_1__1__94_left_grid_pin_30_;
  wire [0:0] cby_1__1__94_left_grid_pin_31_;
  wire [0:0] cby_1__1__95_ccff_tail;
  wire [0:29] cby_1__1__95_chany_bottom_out;
  wire [0:29] cby_1__1__95_chany_top_out;
  wire [0:0] cby_1__1__95_left_grid_pin_16_;
  wire [0:0] cby_1__1__95_left_grid_pin_17_;
  wire [0:0] cby_1__1__95_left_grid_pin_18_;
  wire [0:0] cby_1__1__95_left_grid_pin_19_;
  wire [0:0] cby_1__1__95_left_grid_pin_20_;
  wire [0:0] cby_1__1__95_left_grid_pin_21_;
  wire [0:0] cby_1__1__95_left_grid_pin_22_;
  wire [0:0] cby_1__1__95_left_grid_pin_23_;
  wire [0:0] cby_1__1__95_left_grid_pin_24_;
  wire [0:0] cby_1__1__95_left_grid_pin_25_;
  wire [0:0] cby_1__1__95_left_grid_pin_26_;
  wire [0:0] cby_1__1__95_left_grid_pin_27_;
  wire [0:0] cby_1__1__95_left_grid_pin_28_;
  wire [0:0] cby_1__1__95_left_grid_pin_29_;
  wire [0:0] cby_1__1__95_left_grid_pin_30_;
  wire [0:0] cby_1__1__95_left_grid_pin_31_;
  wire [0:0] cby_1__1__96_ccff_tail;
  wire [0:29] cby_1__1__96_chany_bottom_out;
  wire [0:29] cby_1__1__96_chany_top_out;
  wire [0:0] cby_1__1__96_left_grid_pin_16_;
  wire [0:0] cby_1__1__96_left_grid_pin_17_;
  wire [0:0] cby_1__1__96_left_grid_pin_18_;
  wire [0:0] cby_1__1__96_left_grid_pin_19_;
  wire [0:0] cby_1__1__96_left_grid_pin_20_;
  wire [0:0] cby_1__1__96_left_grid_pin_21_;
  wire [0:0] cby_1__1__96_left_grid_pin_22_;
  wire [0:0] cby_1__1__96_left_grid_pin_23_;
  wire [0:0] cby_1__1__96_left_grid_pin_24_;
  wire [0:0] cby_1__1__96_left_grid_pin_25_;
  wire [0:0] cby_1__1__96_left_grid_pin_26_;
  wire [0:0] cby_1__1__96_left_grid_pin_27_;
  wire [0:0] cby_1__1__96_left_grid_pin_28_;
  wire [0:0] cby_1__1__96_left_grid_pin_29_;
  wire [0:0] cby_1__1__96_left_grid_pin_30_;
  wire [0:0] cby_1__1__96_left_grid_pin_31_;
  wire [0:0] cby_1__1__97_ccff_tail;
  wire [0:29] cby_1__1__97_chany_bottom_out;
  wire [0:29] cby_1__1__97_chany_top_out;
  wire [0:0] cby_1__1__97_left_grid_pin_16_;
  wire [0:0] cby_1__1__97_left_grid_pin_17_;
  wire [0:0] cby_1__1__97_left_grid_pin_18_;
  wire [0:0] cby_1__1__97_left_grid_pin_19_;
  wire [0:0] cby_1__1__97_left_grid_pin_20_;
  wire [0:0] cby_1__1__97_left_grid_pin_21_;
  wire [0:0] cby_1__1__97_left_grid_pin_22_;
  wire [0:0] cby_1__1__97_left_grid_pin_23_;
  wire [0:0] cby_1__1__97_left_grid_pin_24_;
  wire [0:0] cby_1__1__97_left_grid_pin_25_;
  wire [0:0] cby_1__1__97_left_grid_pin_26_;
  wire [0:0] cby_1__1__97_left_grid_pin_27_;
  wire [0:0] cby_1__1__97_left_grid_pin_28_;
  wire [0:0] cby_1__1__97_left_grid_pin_29_;
  wire [0:0] cby_1__1__97_left_grid_pin_30_;
  wire [0:0] cby_1__1__97_left_grid_pin_31_;
  wire [0:0] cby_1__1__98_ccff_tail;
  wire [0:29] cby_1__1__98_chany_bottom_out;
  wire [0:29] cby_1__1__98_chany_top_out;
  wire [0:0] cby_1__1__98_left_grid_pin_16_;
  wire [0:0] cby_1__1__98_left_grid_pin_17_;
  wire [0:0] cby_1__1__98_left_grid_pin_18_;
  wire [0:0] cby_1__1__98_left_grid_pin_19_;
  wire [0:0] cby_1__1__98_left_grid_pin_20_;
  wire [0:0] cby_1__1__98_left_grid_pin_21_;
  wire [0:0] cby_1__1__98_left_grid_pin_22_;
  wire [0:0] cby_1__1__98_left_grid_pin_23_;
  wire [0:0] cby_1__1__98_left_grid_pin_24_;
  wire [0:0] cby_1__1__98_left_grid_pin_25_;
  wire [0:0] cby_1__1__98_left_grid_pin_26_;
  wire [0:0] cby_1__1__98_left_grid_pin_27_;
  wire [0:0] cby_1__1__98_left_grid_pin_28_;
  wire [0:0] cby_1__1__98_left_grid_pin_29_;
  wire [0:0] cby_1__1__98_left_grid_pin_30_;
  wire [0:0] cby_1__1__98_left_grid_pin_31_;
  wire [0:0] cby_1__1__99_ccff_tail;
  wire [0:29] cby_1__1__99_chany_bottom_out;
  wire [0:29] cby_1__1__99_chany_top_out;
  wire [0:0] cby_1__1__99_left_grid_pin_16_;
  wire [0:0] cby_1__1__99_left_grid_pin_17_;
  wire [0:0] cby_1__1__99_left_grid_pin_18_;
  wire [0:0] cby_1__1__99_left_grid_pin_19_;
  wire [0:0] cby_1__1__99_left_grid_pin_20_;
  wire [0:0] cby_1__1__99_left_grid_pin_21_;
  wire [0:0] cby_1__1__99_left_grid_pin_22_;
  wire [0:0] cby_1__1__99_left_grid_pin_23_;
  wire [0:0] cby_1__1__99_left_grid_pin_24_;
  wire [0:0] cby_1__1__99_left_grid_pin_25_;
  wire [0:0] cby_1__1__99_left_grid_pin_26_;
  wire [0:0] cby_1__1__99_left_grid_pin_27_;
  wire [0:0] cby_1__1__99_left_grid_pin_28_;
  wire [0:0] cby_1__1__99_left_grid_pin_29_;
  wire [0:0] cby_1__1__99_left_grid_pin_30_;
  wire [0:0] cby_1__1__99_left_grid_pin_31_;
  wire [0:0] cby_1__1__9_ccff_tail;
  wire [0:29] cby_1__1__9_chany_bottom_out;
  wire [0:29] cby_1__1__9_chany_top_out;
  wire [0:0] cby_1__1__9_left_grid_pin_16_;
  wire [0:0] cby_1__1__9_left_grid_pin_17_;
  wire [0:0] cby_1__1__9_left_grid_pin_18_;
  wire [0:0] cby_1__1__9_left_grid_pin_19_;
  wire [0:0] cby_1__1__9_left_grid_pin_20_;
  wire [0:0] cby_1__1__9_left_grid_pin_21_;
  wire [0:0] cby_1__1__9_left_grid_pin_22_;
  wire [0:0] cby_1__1__9_left_grid_pin_23_;
  wire [0:0] cby_1__1__9_left_grid_pin_24_;
  wire [0:0] cby_1__1__9_left_grid_pin_25_;
  wire [0:0] cby_1__1__9_left_grid_pin_26_;
  wire [0:0] cby_1__1__9_left_grid_pin_27_;
  wire [0:0] cby_1__1__9_left_grid_pin_28_;
  wire [0:0] cby_1__1__9_left_grid_pin_29_;
  wire [0:0] cby_1__1__9_left_grid_pin_30_;
  wire [0:0] cby_1__1__9_left_grid_pin_31_;
  wire [0:0] direct_interc_0_out;
  wire [0:0] direct_interc_100_out;
  wire [0:0] direct_interc_101_out;
  wire [0:0] direct_interc_102_out;
  wire [0:0] direct_interc_103_out;
  wire [0:0] direct_interc_104_out;
  wire [0:0] direct_interc_105_out;
  wire [0:0] direct_interc_106_out;
  wire [0:0] direct_interc_107_out;
  wire [0:0] direct_interc_108_out;
  wire [0:0] direct_interc_109_out;
  wire [0:0] direct_interc_10_out;
  wire [0:0] direct_interc_110_out;
  wire [0:0] direct_interc_111_out;
  wire [0:0] direct_interc_112_out;
  wire [0:0] direct_interc_113_out;
  wire [0:0] direct_interc_114_out;
  wire [0:0] direct_interc_115_out;
  wire [0:0] direct_interc_116_out;
  wire [0:0] direct_interc_117_out;
  wire [0:0] direct_interc_118_out;
  wire [0:0] direct_interc_119_out;
  wire [0:0] direct_interc_11_out;
  wire [0:0] direct_interc_120_out;
  wire [0:0] direct_interc_121_out;
  wire [0:0] direct_interc_122_out;
  wire [0:0] direct_interc_123_out;
  wire [0:0] direct_interc_124_out;
  wire [0:0] direct_interc_125_out;
  wire [0:0] direct_interc_126_out;
  wire [0:0] direct_interc_127_out;
  wire [0:0] direct_interc_128_out;
  wire [0:0] direct_interc_129_out;
  wire [0:0] direct_interc_12_out;
  wire [0:0] direct_interc_130_out;
  wire [0:0] direct_interc_131_out;
  wire [0:0] direct_interc_132_out;
  wire [0:0] direct_interc_133_out;
  wire [0:0] direct_interc_134_out;
  wire [0:0] direct_interc_135_out;
  wire [0:0] direct_interc_136_out;
  wire [0:0] direct_interc_137_out;
  wire [0:0] direct_interc_138_out;
  wire [0:0] direct_interc_139_out;
  wire [0:0] direct_interc_13_out;
  wire [0:0] direct_interc_140_out;
  wire [0:0] direct_interc_141_out;
  wire [0:0] direct_interc_142_out;
  wire [0:0] direct_interc_143_out;
  wire [0:0] direct_interc_144_out;
  wire [0:0] direct_interc_145_out;
  wire [0:0] direct_interc_146_out;
  wire [0:0] direct_interc_147_out;
  wire [0:0] direct_interc_148_out;
  wire [0:0] direct_interc_149_out;
  wire [0:0] direct_interc_14_out;
  wire [0:0] direct_interc_150_out;
  wire [0:0] direct_interc_151_out;
  wire [0:0] direct_interc_152_out;
  wire [0:0] direct_interc_153_out;
  wire [0:0] direct_interc_154_out;
  wire [0:0] direct_interc_155_out;
  wire [0:0] direct_interc_156_out;
  wire [0:0] direct_interc_157_out;
  wire [0:0] direct_interc_158_out;
  wire [0:0] direct_interc_159_out;
  wire [0:0] direct_interc_15_out;
  wire [0:0] direct_interc_160_out;
  wire [0:0] direct_interc_161_out;
  wire [0:0] direct_interc_162_out;
  wire [0:0] direct_interc_163_out;
  wire [0:0] direct_interc_164_out;
  wire [0:0] direct_interc_165_out;
  wire [0:0] direct_interc_166_out;
  wire [0:0] direct_interc_167_out;
  wire [0:0] direct_interc_168_out;
  wire [0:0] direct_interc_169_out;
  wire [0:0] direct_interc_16_out;
  wire [0:0] direct_interc_170_out;
  wire [0:0] direct_interc_171_out;
  wire [0:0] direct_interc_172_out;
  wire [0:0] direct_interc_173_out;
  wire [0:0] direct_interc_174_out;
  wire [0:0] direct_interc_175_out;
  wire [0:0] direct_interc_176_out;
  wire [0:0] direct_interc_177_out;
  wire [0:0] direct_interc_178_out;
  wire [0:0] direct_interc_179_out;
  wire [0:0] direct_interc_17_out;
  wire [0:0] direct_interc_180_out;
  wire [0:0] direct_interc_181_out;
  wire [0:0] direct_interc_182_out;
  wire [0:0] direct_interc_183_out;
  wire [0:0] direct_interc_184_out;
  wire [0:0] direct_interc_185_out;
  wire [0:0] direct_interc_186_out;
  wire [0:0] direct_interc_187_out;
  wire [0:0] direct_interc_188_out;
  wire [0:0] direct_interc_189_out;
  wire [0:0] direct_interc_18_out;
  wire [0:0] direct_interc_190_out;
  wire [0:0] direct_interc_191_out;
  wire [0:0] direct_interc_192_out;
  wire [0:0] direct_interc_193_out;
  wire [0:0] direct_interc_194_out;
  wire [0:0] direct_interc_195_out;
  wire [0:0] direct_interc_196_out;
  wire [0:0] direct_interc_197_out;
  wire [0:0] direct_interc_198_out;
  wire [0:0] direct_interc_199_out;
  wire [0:0] direct_interc_19_out;
  wire [0:0] direct_interc_1_out;
  wire [0:0] direct_interc_200_out;
  wire [0:0] direct_interc_201_out;
  wire [0:0] direct_interc_202_out;
  wire [0:0] direct_interc_203_out;
  wire [0:0] direct_interc_204_out;
  wire [0:0] direct_interc_205_out;
  wire [0:0] direct_interc_206_out;
  wire [0:0] direct_interc_207_out;
  wire [0:0] direct_interc_208_out;
  wire [0:0] direct_interc_209_out;
  wire [0:0] direct_interc_20_out;
  wire [0:0] direct_interc_210_out;
  wire [0:0] direct_interc_211_out;
  wire [0:0] direct_interc_212_out;
  wire [0:0] direct_interc_213_out;
  wire [0:0] direct_interc_214_out;
  wire [0:0] direct_interc_215_out;
  wire [0:0] direct_interc_216_out;
  wire [0:0] direct_interc_217_out;
  wire [0:0] direct_interc_218_out;
  wire [0:0] direct_interc_219_out;
  wire [0:0] direct_interc_21_out;
  wire [0:0] direct_interc_220_out;
  wire [0:0] direct_interc_221_out;
  wire [0:0] direct_interc_222_out;
  wire [0:0] direct_interc_223_out;
  wire [0:0] direct_interc_224_out;
  wire [0:0] direct_interc_225_out;
  wire [0:0] direct_interc_226_out;
  wire [0:0] direct_interc_227_out;
  wire [0:0] direct_interc_228_out;
  wire [0:0] direct_interc_229_out;
  wire [0:0] direct_interc_22_out;
  wire [0:0] direct_interc_230_out;
  wire [0:0] direct_interc_231_out;
  wire [0:0] direct_interc_232_out;
  wire [0:0] direct_interc_233_out;
  wire [0:0] direct_interc_234_out;
  wire [0:0] direct_interc_235_out;
  wire [0:0] direct_interc_236_out;
  wire [0:0] direct_interc_237_out;
  wire [0:0] direct_interc_238_out;
  wire [0:0] direct_interc_239_out;
  wire [0:0] direct_interc_23_out;
  wire [0:0] direct_interc_240_out;
  wire [0:0] direct_interc_241_out;
  wire [0:0] direct_interc_242_out;
  wire [0:0] direct_interc_243_out;
  wire [0:0] direct_interc_244_out;
  wire [0:0] direct_interc_245_out;
  wire [0:0] direct_interc_246_out;
  wire [0:0] direct_interc_247_out;
  wire [0:0] direct_interc_248_out;
  wire [0:0] direct_interc_249_out;
  wire [0:0] direct_interc_24_out;
  wire [0:0] direct_interc_250_out;
  wire [0:0] direct_interc_251_out;
  wire [0:0] direct_interc_252_out;
  wire [0:0] direct_interc_253_out;
  wire [0:0] direct_interc_254_out;
  wire [0:0] direct_interc_255_out;
  wire [0:0] direct_interc_256_out;
  wire [0:0] direct_interc_257_out;
  wire [0:0] direct_interc_258_out;
  wire [0:0] direct_interc_259_out;
  wire [0:0] direct_interc_25_out;
  wire [0:0] direct_interc_260_out;
  wire [0:0] direct_interc_261_out;
  wire [0:0] direct_interc_262_out;
  wire [0:0] direct_interc_263_out;
  wire [0:0] direct_interc_264_out;
  wire [0:0] direct_interc_265_out;
  wire [0:0] direct_interc_266_out;
  wire [0:0] direct_interc_267_out;
  wire [0:0] direct_interc_268_out;
  wire [0:0] direct_interc_269_out;
  wire [0:0] direct_interc_26_out;
  wire [0:0] direct_interc_270_out;
  wire [0:0] direct_interc_271_out;
  wire [0:0] direct_interc_272_out;
  wire [0:0] direct_interc_273_out;
  wire [0:0] direct_interc_274_out;
  wire [0:0] direct_interc_275_out;
  wire [0:0] direct_interc_276_out;
  wire [0:0] direct_interc_277_out;
  wire [0:0] direct_interc_278_out;
  wire [0:0] direct_interc_279_out;
  wire [0:0] direct_interc_27_out;
  wire [0:0] direct_interc_280_out;
  wire [0:0] direct_interc_281_out;
  wire [0:0] direct_interc_282_out;
  wire [0:0] direct_interc_283_out;
  wire [0:0] direct_interc_284_out;
  wire [0:0] direct_interc_285_out;
  wire [0:0] direct_interc_286_out;
  wire [0:0] direct_interc_287_out;
  wire [0:0] direct_interc_288_out;
  wire [0:0] direct_interc_289_out;
  wire [0:0] direct_interc_28_out;
  wire [0:0] direct_interc_290_out;
  wire [0:0] direct_interc_291_out;
  wire [0:0] direct_interc_292_out;
  wire [0:0] direct_interc_293_out;
  wire [0:0] direct_interc_294_out;
  wire [0:0] direct_interc_295_out;
  wire [0:0] direct_interc_296_out;
  wire [0:0] direct_interc_297_out;
  wire [0:0] direct_interc_298_out;
  wire [0:0] direct_interc_299_out;
  wire [0:0] direct_interc_29_out;
  wire [0:0] direct_interc_2_out;
  wire [0:0] direct_interc_300_out;
  wire [0:0] direct_interc_301_out;
  wire [0:0] direct_interc_302_out;
  wire [0:0] direct_interc_303_out;
  wire [0:0] direct_interc_304_out;
  wire [0:0] direct_interc_305_out;
  wire [0:0] direct_interc_306_out;
  wire [0:0] direct_interc_307_out;
  wire [0:0] direct_interc_308_out;
  wire [0:0] direct_interc_309_out;
  wire [0:0] direct_interc_30_out;
  wire [0:0] direct_interc_310_out;
  wire [0:0] direct_interc_311_out;
  wire [0:0] direct_interc_312_out;
  wire [0:0] direct_interc_313_out;
  wire [0:0] direct_interc_314_out;
  wire [0:0] direct_interc_315_out;
  wire [0:0] direct_interc_316_out;
  wire [0:0] direct_interc_317_out;
  wire [0:0] direct_interc_318_out;
  wire [0:0] direct_interc_319_out;
  wire [0:0] direct_interc_31_out;
  wire [0:0] direct_interc_320_out;
  wire [0:0] direct_interc_321_out;
  wire [0:0] direct_interc_322_out;
  wire [0:0] direct_interc_323_out;
  wire [0:0] direct_interc_324_out;
  wire [0:0] direct_interc_325_out;
  wire [0:0] direct_interc_326_out;
  wire [0:0] direct_interc_327_out;
  wire [0:0] direct_interc_328_out;
  wire [0:0] direct_interc_329_out;
  wire [0:0] direct_interc_32_out;
  wire [0:0] direct_interc_330_out;
  wire [0:0] direct_interc_331_out;
  wire [0:0] direct_interc_332_out;
  wire [0:0] direct_interc_333_out;
  wire [0:0] direct_interc_334_out;
  wire [0:0] direct_interc_335_out;
  wire [0:0] direct_interc_336_out;
  wire [0:0] direct_interc_337_out;
  wire [0:0] direct_interc_338_out;
  wire [0:0] direct_interc_339_out;
  wire [0:0] direct_interc_33_out;
  wire [0:0] direct_interc_340_out;
  wire [0:0] direct_interc_341_out;
  wire [0:0] direct_interc_342_out;
  wire [0:0] direct_interc_343_out;
  wire [0:0] direct_interc_344_out;
  wire [0:0] direct_interc_345_out;
  wire [0:0] direct_interc_346_out;
  wire [0:0] direct_interc_347_out;
  wire [0:0] direct_interc_348_out;
  wire [0:0] direct_interc_349_out;
  wire [0:0] direct_interc_34_out;
  wire [0:0] direct_interc_350_out;
  wire [0:0] direct_interc_351_out;
  wire [0:0] direct_interc_352_out;
  wire [0:0] direct_interc_353_out;
  wire [0:0] direct_interc_354_out;
  wire [0:0] direct_interc_355_out;
  wire [0:0] direct_interc_356_out;
  wire [0:0] direct_interc_357_out;
  wire [0:0] direct_interc_358_out;
  wire [0:0] direct_interc_359_out;
  wire [0:0] direct_interc_35_out;
  wire [0:0] direct_interc_360_out;
  wire [0:0] direct_interc_361_out;
  wire [0:0] direct_interc_362_out;
  wire [0:0] direct_interc_363_out;
  wire [0:0] direct_interc_364_out;
  wire [0:0] direct_interc_365_out;
  wire [0:0] direct_interc_366_out;
  wire [0:0] direct_interc_367_out;
  wire [0:0] direct_interc_368_out;
  wire [0:0] direct_interc_369_out;
  wire [0:0] direct_interc_36_out;
  wire [0:0] direct_interc_370_out;
  wire [0:0] direct_interc_371_out;
  wire [0:0] direct_interc_372_out;
  wire [0:0] direct_interc_373_out;
  wire [0:0] direct_interc_374_out;
  wire [0:0] direct_interc_375_out;
  wire [0:0] direct_interc_376_out;
  wire [0:0] direct_interc_377_out;
  wire [0:0] direct_interc_378_out;
  wire [0:0] direct_interc_379_out;
  wire [0:0] direct_interc_37_out;
  wire [0:0] direct_interc_380_out;
  wire [0:0] direct_interc_381_out;
  wire [0:0] direct_interc_382_out;
  wire [0:0] direct_interc_383_out;
  wire [0:0] direct_interc_384_out;
  wire [0:0] direct_interc_385_out;
  wire [0:0] direct_interc_386_out;
  wire [0:0] direct_interc_387_out;
  wire [0:0] direct_interc_388_out;
  wire [0:0] direct_interc_389_out;
  wire [0:0] direct_interc_38_out;
  wire [0:0] direct_interc_390_out;
  wire [0:0] direct_interc_391_out;
  wire [0:0] direct_interc_392_out;
  wire [0:0] direct_interc_393_out;
  wire [0:0] direct_interc_394_out;
  wire [0:0] direct_interc_395_out;
  wire [0:0] direct_interc_396_out;
  wire [0:0] direct_interc_397_out;
  wire [0:0] direct_interc_398_out;
  wire [0:0] direct_interc_399_out;
  wire [0:0] direct_interc_39_out;
  wire [0:0] direct_interc_3_out;
  wire [0:0] direct_interc_400_out;
  wire [0:0] direct_interc_401_out;
  wire [0:0] direct_interc_402_out;
  wire [0:0] direct_interc_403_out;
  wire [0:0] direct_interc_404_out;
  wire [0:0] direct_interc_405_out;
  wire [0:0] direct_interc_406_out;
  wire [0:0] direct_interc_40_out;
  wire [0:0] direct_interc_41_out;
  wire [0:0] direct_interc_42_out;
  wire [0:0] direct_interc_43_out;
  wire [0:0] direct_interc_44_out;
  wire [0:0] direct_interc_45_out;
  wire [0:0] direct_interc_46_out;
  wire [0:0] direct_interc_47_out;
  wire [0:0] direct_interc_48_out;
  wire [0:0] direct_interc_49_out;
  wire [0:0] direct_interc_4_out;
  wire [0:0] direct_interc_50_out;
  wire [0:0] direct_interc_51_out;
  wire [0:0] direct_interc_52_out;
  wire [0:0] direct_interc_53_out;
  wire [0:0] direct_interc_54_out;
  wire [0:0] direct_interc_55_out;
  wire [0:0] direct_interc_56_out;
  wire [0:0] direct_interc_57_out;
  wire [0:0] direct_interc_58_out;
  wire [0:0] direct_interc_59_out;
  wire [0:0] direct_interc_5_out;
  wire [0:0] direct_interc_60_out;
  wire [0:0] direct_interc_61_out;
  wire [0:0] direct_interc_62_out;
  wire [0:0] direct_interc_63_out;
  wire [0:0] direct_interc_64_out;
  wire [0:0] direct_interc_65_out;
  wire [0:0] direct_interc_66_out;
  wire [0:0] direct_interc_67_out;
  wire [0:0] direct_interc_68_out;
  wire [0:0] direct_interc_69_out;
  wire [0:0] direct_interc_6_out;
  wire [0:0] direct_interc_70_out;
  wire [0:0] direct_interc_71_out;
  wire [0:0] direct_interc_72_out;
  wire [0:0] direct_interc_73_out;
  wire [0:0] direct_interc_74_out;
  wire [0:0] direct_interc_75_out;
  wire [0:0] direct_interc_76_out;
  wire [0:0] direct_interc_77_out;
  wire [0:0] direct_interc_78_out;
  wire [0:0] direct_interc_79_out;
  wire [0:0] direct_interc_7_out;
  wire [0:0] direct_interc_80_out;
  wire [0:0] direct_interc_81_out;
  wire [0:0] direct_interc_82_out;
  wire [0:0] direct_interc_83_out;
  wire [0:0] direct_interc_84_out;
  wire [0:0] direct_interc_85_out;
  wire [0:0] direct_interc_86_out;
  wire [0:0] direct_interc_87_out;
  wire [0:0] direct_interc_88_out;
  wire [0:0] direct_interc_89_out;
  wire [0:0] direct_interc_8_out;
  wire [0:0] direct_interc_90_out;
  wire [0:0] direct_interc_91_out;
  wire [0:0] direct_interc_92_out;
  wire [0:0] direct_interc_93_out;
  wire [0:0] direct_interc_94_out;
  wire [0:0] direct_interc_95_out;
  wire [0:0] direct_interc_96_out;
  wire [0:0] direct_interc_97_out;
  wire [0:0] direct_interc_98_out;
  wire [0:0] direct_interc_99_out;
  wire [0:0] direct_interc_9_out;
  wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_0_ccff_tail;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_100_ccff_tail;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_100_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_100_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_101_ccff_tail;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_101_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_101_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_102_ccff_tail;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_102_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_102_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_103_ccff_tail;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_103_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_103_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_104_ccff_tail;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_104_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_104_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_105_ccff_tail;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_105_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_105_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_106_ccff_tail;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_106_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_106_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_107_ccff_tail;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_107_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_107_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_108_ccff_tail;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_108_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_108_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_109_ccff_tail;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_109_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_109_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_10__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_10__12__undriven_top_width_0_height_0__pin_34_;
  wire [0:0] grid_clb_10__1__undriven_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_10__1__undriven_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_10_ccff_tail;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_110_ccff_tail;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_110_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_110_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_111_ccff_tail;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_111_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_111_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_112_ccff_tail;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_112_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_112_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_113_ccff_tail;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_113_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_113_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_114_ccff_tail;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_114_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_114_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_115_ccff_tail;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_115_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_115_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_116_ccff_tail;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_116_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_116_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_117_ccff_tail;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_117_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_117_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_118_ccff_tail;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_118_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_118_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_119_ccff_tail;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_119_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_119_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_11__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_11__12__undriven_top_width_0_height_0__pin_34_;
  wire [0:0] grid_clb_11__1__undriven_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_11__1__undriven_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_11_ccff_tail;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_120_ccff_tail;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_120_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_120_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_121_ccff_tail;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_121_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_121_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_122_ccff_tail;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_122_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_122_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_123_ccff_tail;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_123_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_123_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_124_ccff_tail;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_124_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_124_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_125_ccff_tail;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_125_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_125_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_126_ccff_tail;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_126_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_126_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_127_ccff_tail;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_127_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_127_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_128_ccff_tail;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_128_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_128_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_129_ccff_tail;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_129_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_129_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_12__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_12__12__undriven_top_width_0_height_0__pin_34_;
  wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_12_ccff_tail;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_130_ccff_tail;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_130_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_130_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_131_ccff_tail;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_131_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_131_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_132_ccff_tail;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_132_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_132_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_133_ccff_tail;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_133_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_133_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_134_ccff_tail;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_134_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_134_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_135_ccff_tail;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_135_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_135_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_136_ccff_tail;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_136_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_136_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_137_ccff_tail;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_137_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_137_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_138_ccff_tail;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_138_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_138_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_139_ccff_tail;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_139_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_139_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_13_ccff_tail;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_140_ccff_tail;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_140_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_140_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_141_ccff_tail;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_141_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_141_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_142_ccff_tail;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_142_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_142_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_143_ccff_tail;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_143_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_143_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_14_ccff_tail;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_15_ccff_tail;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_16_ccff_tail;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_17_ccff_tail;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_18_ccff_tail;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_19_ccff_tail;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_1__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_1__12__undriven_top_width_0_height_0__pin_33_;
  wire [0:0] grid_clb_1__12__undriven_top_width_0_height_0__pin_34_;
  wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_1_ccff_tail;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_20_ccff_tail;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_21_ccff_tail;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_22_ccff_tail;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_23_ccff_tail;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_24_ccff_tail;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_25_ccff_tail;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_26_ccff_tail;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_27_ccff_tail;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_28_ccff_tail;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_29_ccff_tail;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_2__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_2__12__undriven_top_width_0_height_0__pin_34_;
  wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_2_ccff_tail;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_30_ccff_tail;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_31_ccff_tail;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_32_ccff_tail;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_33_ccff_tail;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_34_ccff_tail;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_35_ccff_tail;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_36_ccff_tail;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_37_ccff_tail;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_38_ccff_tail;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_39_ccff_tail;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_3__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_3__12__undriven_top_width_0_height_0__pin_34_;
  wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_3_ccff_tail;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_40_ccff_tail;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_41_ccff_tail;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_42_ccff_tail;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_43_ccff_tail;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_44_ccff_tail;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_45_ccff_tail;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_46_ccff_tail;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_47_ccff_tail;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_48_ccff_tail;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_49_ccff_tail;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_4__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_4__12__undriven_top_width_0_height_0__pin_34_;
  wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_4_ccff_tail;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_50_ccff_tail;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_51_ccff_tail;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_52_ccff_tail;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_53_ccff_tail;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_54_ccff_tail;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_55_ccff_tail;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_56_ccff_tail;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_57_ccff_tail;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_58_ccff_tail;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_59_ccff_tail;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_5__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_5__12__undriven_top_width_0_height_0__pin_34_;
  wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_5_ccff_tail;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_60_ccff_tail;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_61_ccff_tail;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_62_ccff_tail;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_63_ccff_tail;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_64_ccff_tail;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_64_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_64_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_65_ccff_tail;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_65_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_65_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_66_ccff_tail;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_66_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_66_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_67_ccff_tail;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_67_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_67_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_68_ccff_tail;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_68_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_68_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_69_ccff_tail;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_69_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_69_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_6__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_6__12__undriven_top_width_0_height_0__pin_34_;
  wire [0:0] grid_clb_6__1__undriven_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_6__1__undriven_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_6_ccff_tail;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_70_ccff_tail;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_70_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_70_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_71_ccff_tail;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_71_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_71_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_72_ccff_tail;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_72_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_72_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_73_ccff_tail;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_73_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_73_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_74_ccff_tail;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_74_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_74_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_75_ccff_tail;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_75_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_75_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_76_ccff_tail;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_76_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_76_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_77_ccff_tail;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_77_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_77_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_78_ccff_tail;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_78_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_78_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_79_ccff_tail;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_79_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_79_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_7__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_7__12__undriven_top_width_0_height_0__pin_34_;
  wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_7_ccff_tail;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_80_ccff_tail;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_80_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_80_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_81_ccff_tail;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_81_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_81_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_82_ccff_tail;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_82_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_82_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_83_ccff_tail;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_83_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_83_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_84_ccff_tail;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_84_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_84_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_85_ccff_tail;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_85_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_85_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_86_ccff_tail;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_86_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_86_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_87_ccff_tail;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_87_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_87_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_88_ccff_tail;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_88_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_88_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_89_ccff_tail;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_89_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_89_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_8__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_8__12__undriven_top_width_0_height_0__pin_34_;
  wire [0:0] grid_clb_8__1__undriven_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_8__1__undriven_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_8_ccff_tail;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_90_ccff_tail;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_90_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_90_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_91_ccff_tail;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_91_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_91_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_92_ccff_tail;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_92_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_92_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_93_ccff_tail;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_93_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_93_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_94_ccff_tail;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_94_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_94_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_95_ccff_tail;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_95_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_95_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_96_ccff_tail;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_96_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_96_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_97_ccff_tail;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_97_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_97_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_98_ccff_tail;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_98_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_98_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_99_ccff_tail;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_99_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_99_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_9__12__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_9__12__undriven_top_width_0_height_0__pin_34_;
  wire [0:0] grid_clb_9__1__undriven_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_9__1__undriven_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_52_;
  wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_53_;
  wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_54_;
  wire [0:0] grid_clb_9_ccff_tail;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_50_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_50_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_51_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_51_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_43_upper;
  wire [0:0] grid_io_bottom_0_ccff_tail;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_10_ccff_tail;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_11_ccff_tail;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_1_ccff_tail;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_2_ccff_tail;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_3_ccff_tail;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_4_ccff_tail;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_5_ccff_tail;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_6_ccff_tail;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_7_ccff_tail;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_8_ccff_tail;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_9_ccff_tail;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_left_0_ccff_tail;
  wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_10_ccff_tail;
  wire [0:0] grid_io_left_10_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_10_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_11_ccff_tail;
  wire [0:0] grid_io_left_11_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_11_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_1_ccff_tail;
  wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_2_ccff_tail;
  wire [0:0] grid_io_left_2_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_2_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_3_ccff_tail;
  wire [0:0] grid_io_left_3_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_3_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_4_ccff_tail;
  wire [0:0] grid_io_left_4_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_4_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_5_ccff_tail;
  wire [0:0] grid_io_left_5_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_5_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_6_ccff_tail;
  wire [0:0] grid_io_left_6_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_6_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_7_ccff_tail;
  wire [0:0] grid_io_left_7_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_7_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_8_ccff_tail;
  wire [0:0] grid_io_left_8_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_8_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_9_ccff_tail;
  wire [0:0] grid_io_left_9_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_9_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_0_ccff_tail;
  wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_10_ccff_tail;
  wire [0:0] grid_io_right_10_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_10_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_11_ccff_tail;
  wire [0:0] grid_io_right_11_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_11_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_1_ccff_tail;
  wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_2_ccff_tail;
  wire [0:0] grid_io_right_2_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_2_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_3_ccff_tail;
  wire [0:0] grid_io_right_3_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_3_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_4_ccff_tail;
  wire [0:0] grid_io_right_4_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_4_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_5_ccff_tail;
  wire [0:0] grid_io_right_5_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_5_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_6_ccff_tail;
  wire [0:0] grid_io_right_6_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_6_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_7_ccff_tail;
  wire [0:0] grid_io_right_7_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_7_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_8_ccff_tail;
  wire [0:0] grid_io_right_8_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_8_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_9_ccff_tail;
  wire [0:0] grid_io_right_9_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_9_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_0_ccff_tail;
  wire [0:0] grid_io_top_10_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_10_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_10_ccff_tail;
  wire [0:0] grid_io_top_11_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_11_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_11_ccff_tail;
  wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_1_ccff_tail;
  wire [0:0] grid_io_top_2_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_2_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_2_ccff_tail;
  wire [0:0] grid_io_top_3_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_3_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_3_ccff_tail;
  wire [0:0] grid_io_top_4_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_4_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_4_ccff_tail;
  wire [0:0] grid_io_top_5_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_5_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_5_ccff_tail;
  wire [0:0] grid_io_top_6_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_6_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_6_ccff_tail;
  wire [0:0] grid_io_top_7_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_7_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_7_ccff_tail;
  wire [0:0] grid_io_top_8_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_8_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_8_ccff_tail;
  wire [0:0] grid_io_top_9_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_9_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_9_ccff_tail;
  wire [0:29] sb_0__0__0_chanx_right_out;
  wire [0:29] sb_0__0__0_chany_top_out;
  wire [0:0] sb_0__12__0_ccff_tail;
  wire [0:29] sb_0__12__0_chanx_right_out;
  wire [0:29] sb_0__12__0_chany_bottom_out;
  wire [0:0] sb_0__1__0_ccff_tail;
  wire [0:29] sb_0__1__0_chanx_right_out;
  wire [0:29] sb_0__1__0_chany_bottom_out;
  wire [0:29] sb_0__1__0_chany_top_out;
  wire [0:0] sb_0__1__10_ccff_tail;
  wire [0:29] sb_0__1__10_chanx_right_out;
  wire [0:29] sb_0__1__10_chany_bottom_out;
  wire [0:29] sb_0__1__10_chany_top_out;
  wire [0:0] sb_0__1__1_ccff_tail;
  wire [0:29] sb_0__1__1_chanx_right_out;
  wire [0:29] sb_0__1__1_chany_bottom_out;
  wire [0:29] sb_0__1__1_chany_top_out;
  wire [0:0] sb_0__1__2_ccff_tail;
  wire [0:29] sb_0__1__2_chanx_right_out;
  wire [0:29] sb_0__1__2_chany_bottom_out;
  wire [0:29] sb_0__1__2_chany_top_out;
  wire [0:0] sb_0__1__3_ccff_tail;
  wire [0:29] sb_0__1__3_chanx_right_out;
  wire [0:29] sb_0__1__3_chany_bottom_out;
  wire [0:29] sb_0__1__3_chany_top_out;
  wire [0:0] sb_0__1__4_ccff_tail;
  wire [0:29] sb_0__1__4_chanx_right_out;
  wire [0:29] sb_0__1__4_chany_bottom_out;
  wire [0:29] sb_0__1__4_chany_top_out;
  wire [0:0] sb_0__1__5_ccff_tail;
  wire [0:29] sb_0__1__5_chanx_right_out;
  wire [0:29] sb_0__1__5_chany_bottom_out;
  wire [0:29] sb_0__1__5_chany_top_out;
  wire [0:0] sb_0__1__6_ccff_tail;
  wire [0:29] sb_0__1__6_chanx_right_out;
  wire [0:29] sb_0__1__6_chany_bottom_out;
  wire [0:29] sb_0__1__6_chany_top_out;
  wire [0:0] sb_0__1__7_ccff_tail;
  wire [0:29] sb_0__1__7_chanx_right_out;
  wire [0:29] sb_0__1__7_chany_bottom_out;
  wire [0:29] sb_0__1__7_chany_top_out;
  wire [0:0] sb_0__1__8_ccff_tail;
  wire [0:29] sb_0__1__8_chanx_right_out;
  wire [0:29] sb_0__1__8_chany_bottom_out;
  wire [0:29] sb_0__1__8_chany_top_out;
  wire [0:0] sb_0__1__9_ccff_tail;
  wire [0:29] sb_0__1__9_chanx_right_out;
  wire [0:29] sb_0__1__9_chany_bottom_out;
  wire [0:29] sb_0__1__9_chany_top_out;
  wire [0:0] sb_12__0__0_ccff_tail;
  wire [0:29] sb_12__0__0_chanx_left_out;
  wire [0:29] sb_12__0__0_chany_top_out;
  wire [0:0] sb_12__12__0_ccff_tail;
  wire [0:29] sb_12__12__0_chanx_left_out;
  wire [0:29] sb_12__12__0_chany_bottom_out;
  wire [0:0] sb_12__1__0_ccff_tail;
  wire [0:29] sb_12__1__0_chanx_left_out;
  wire [0:29] sb_12__1__0_chany_bottom_out;
  wire [0:29] sb_12__1__0_chany_top_out;
  wire [0:0] sb_12__1__10_ccff_tail;
  wire [0:29] sb_12__1__10_chanx_left_out;
  wire [0:29] sb_12__1__10_chany_bottom_out;
  wire [0:29] sb_12__1__10_chany_top_out;
  wire [0:0] sb_12__1__1_ccff_tail;
  wire [0:29] sb_12__1__1_chanx_left_out;
  wire [0:29] sb_12__1__1_chany_bottom_out;
  wire [0:29] sb_12__1__1_chany_top_out;
  wire [0:0] sb_12__1__2_ccff_tail;
  wire [0:29] sb_12__1__2_chanx_left_out;
  wire [0:29] sb_12__1__2_chany_bottom_out;
  wire [0:29] sb_12__1__2_chany_top_out;
  wire [0:0] sb_12__1__3_ccff_tail;
  wire [0:29] sb_12__1__3_chanx_left_out;
  wire [0:29] sb_12__1__3_chany_bottom_out;
  wire [0:29] sb_12__1__3_chany_top_out;
  wire [0:0] sb_12__1__4_ccff_tail;
  wire [0:29] sb_12__1__4_chanx_left_out;
  wire [0:29] sb_12__1__4_chany_bottom_out;
  wire [0:29] sb_12__1__4_chany_top_out;
  wire [0:0] sb_12__1__5_ccff_tail;
  wire [0:29] sb_12__1__5_chanx_left_out;
  wire [0:29] sb_12__1__5_chany_bottom_out;
  wire [0:29] sb_12__1__5_chany_top_out;
  wire [0:0] sb_12__1__6_ccff_tail;
  wire [0:29] sb_12__1__6_chanx_left_out;
  wire [0:29] sb_12__1__6_chany_bottom_out;
  wire [0:29] sb_12__1__6_chany_top_out;
  wire [0:0] sb_12__1__7_ccff_tail;
  wire [0:29] sb_12__1__7_chanx_left_out;
  wire [0:29] sb_12__1__7_chany_bottom_out;
  wire [0:29] sb_12__1__7_chany_top_out;
  wire [0:0] sb_12__1__8_ccff_tail;
  wire [0:29] sb_12__1__8_chanx_left_out;
  wire [0:29] sb_12__1__8_chany_bottom_out;
  wire [0:29] sb_12__1__8_chany_top_out;
  wire [0:0] sb_12__1__9_ccff_tail;
  wire [0:29] sb_12__1__9_chanx_left_out;
  wire [0:29] sb_12__1__9_chany_bottom_out;
  wire [0:29] sb_12__1__9_chany_top_out;
  wire [0:0] sb_1__0__0_ccff_tail;
  wire [0:29] sb_1__0__0_chanx_left_out;
  wire [0:29] sb_1__0__0_chanx_right_out;
  wire [0:29] sb_1__0__0_chany_top_out;
  wire [0:0] sb_1__0__10_ccff_tail;
  wire [0:29] sb_1__0__10_chanx_left_out;
  wire [0:29] sb_1__0__10_chanx_right_out;
  wire [0:29] sb_1__0__10_chany_top_out;
  wire [0:0] sb_1__0__1_ccff_tail;
  wire [0:29] sb_1__0__1_chanx_left_out;
  wire [0:29] sb_1__0__1_chanx_right_out;
  wire [0:29] sb_1__0__1_chany_top_out;
  wire [0:0] sb_1__0__2_ccff_tail;
  wire [0:29] sb_1__0__2_chanx_left_out;
  wire [0:29] sb_1__0__2_chanx_right_out;
  wire [0:29] sb_1__0__2_chany_top_out;
  wire [0:0] sb_1__0__3_ccff_tail;
  wire [0:29] sb_1__0__3_chanx_left_out;
  wire [0:29] sb_1__0__3_chanx_right_out;
  wire [0:29] sb_1__0__3_chany_top_out;
  wire [0:0] sb_1__0__4_ccff_tail;
  wire [0:29] sb_1__0__4_chanx_left_out;
  wire [0:29] sb_1__0__4_chanx_right_out;
  wire [0:29] sb_1__0__4_chany_top_out;
  wire [0:0] sb_1__0__5_ccff_tail;
  wire [0:29] sb_1__0__5_chanx_left_out;
  wire [0:29] sb_1__0__5_chanx_right_out;
  wire [0:29] sb_1__0__5_chany_top_out;
  wire [0:0] sb_1__0__6_ccff_tail;
  wire [0:29] sb_1__0__6_chanx_left_out;
  wire [0:29] sb_1__0__6_chanx_right_out;
  wire [0:29] sb_1__0__6_chany_top_out;
  wire [0:0] sb_1__0__7_ccff_tail;
  wire [0:29] sb_1__0__7_chanx_left_out;
  wire [0:29] sb_1__0__7_chanx_right_out;
  wire [0:29] sb_1__0__7_chany_top_out;
  wire [0:0] sb_1__0__8_ccff_tail;
  wire [0:29] sb_1__0__8_chanx_left_out;
  wire [0:29] sb_1__0__8_chanx_right_out;
  wire [0:29] sb_1__0__8_chany_top_out;
  wire [0:0] sb_1__0__9_ccff_tail;
  wire [0:29] sb_1__0__9_chanx_left_out;
  wire [0:29] sb_1__0__9_chanx_right_out;
  wire [0:29] sb_1__0__9_chany_top_out;
  wire [0:0] sb_1__12__0_ccff_tail;
  wire [0:29] sb_1__12__0_chanx_left_out;
  wire [0:29] sb_1__12__0_chanx_right_out;
  wire [0:29] sb_1__12__0_chany_bottom_out;
  wire [0:0] sb_1__12__10_ccff_tail;
  wire [0:29] sb_1__12__10_chanx_left_out;
  wire [0:29] sb_1__12__10_chanx_right_out;
  wire [0:29] sb_1__12__10_chany_bottom_out;
  wire [0:0] sb_1__12__1_ccff_tail;
  wire [0:29] sb_1__12__1_chanx_left_out;
  wire [0:29] sb_1__12__1_chanx_right_out;
  wire [0:29] sb_1__12__1_chany_bottom_out;
  wire [0:0] sb_1__12__2_ccff_tail;
  wire [0:29] sb_1__12__2_chanx_left_out;
  wire [0:29] sb_1__12__2_chanx_right_out;
  wire [0:29] sb_1__12__2_chany_bottom_out;
  wire [0:0] sb_1__12__3_ccff_tail;
  wire [0:29] sb_1__12__3_chanx_left_out;
  wire [0:29] sb_1__12__3_chanx_right_out;
  wire [0:29] sb_1__12__3_chany_bottom_out;
  wire [0:0] sb_1__12__4_ccff_tail;
  wire [0:29] sb_1__12__4_chanx_left_out;
  wire [0:29] sb_1__12__4_chanx_right_out;
  wire [0:29] sb_1__12__4_chany_bottom_out;
  wire [0:0] sb_1__12__5_ccff_tail;
  wire [0:29] sb_1__12__5_chanx_left_out;
  wire [0:29] sb_1__12__5_chanx_right_out;
  wire [0:29] sb_1__12__5_chany_bottom_out;
  wire [0:0] sb_1__12__6_ccff_tail;
  wire [0:29] sb_1__12__6_chanx_left_out;
  wire [0:29] sb_1__12__6_chanx_right_out;
  wire [0:29] sb_1__12__6_chany_bottom_out;
  wire [0:0] sb_1__12__7_ccff_tail;
  wire [0:29] sb_1__12__7_chanx_left_out;
  wire [0:29] sb_1__12__7_chanx_right_out;
  wire [0:29] sb_1__12__7_chany_bottom_out;
  wire [0:0] sb_1__12__8_ccff_tail;
  wire [0:29] sb_1__12__8_chanx_left_out;
  wire [0:29] sb_1__12__8_chanx_right_out;
  wire [0:29] sb_1__12__8_chany_bottom_out;
  wire [0:0] sb_1__12__9_ccff_tail;
  wire [0:29] sb_1__12__9_chanx_left_out;
  wire [0:29] sb_1__12__9_chanx_right_out;
  wire [0:29] sb_1__12__9_chany_bottom_out;
  wire [0:0] sb_1__1__0_ccff_tail;
  wire [0:29] sb_1__1__0_chanx_left_out;
  wire [0:29] sb_1__1__0_chanx_right_out;
  wire [0:29] sb_1__1__0_chany_bottom_out;
  wire [0:29] sb_1__1__0_chany_top_out;
  wire [0:0] sb_1__1__100_ccff_tail;
  wire [0:29] sb_1__1__100_chanx_left_out;
  wire [0:29] sb_1__1__100_chanx_right_out;
  wire [0:29] sb_1__1__100_chany_bottom_out;
  wire [0:29] sb_1__1__100_chany_top_out;
  wire [0:0] sb_1__1__101_ccff_tail;
  wire [0:29] sb_1__1__101_chanx_left_out;
  wire [0:29] sb_1__1__101_chanx_right_out;
  wire [0:29] sb_1__1__101_chany_bottom_out;
  wire [0:29] sb_1__1__101_chany_top_out;
  wire [0:0] sb_1__1__102_ccff_tail;
  wire [0:29] sb_1__1__102_chanx_left_out;
  wire [0:29] sb_1__1__102_chanx_right_out;
  wire [0:29] sb_1__1__102_chany_bottom_out;
  wire [0:29] sb_1__1__102_chany_top_out;
  wire [0:0] sb_1__1__103_ccff_tail;
  wire [0:29] sb_1__1__103_chanx_left_out;
  wire [0:29] sb_1__1__103_chanx_right_out;
  wire [0:29] sb_1__1__103_chany_bottom_out;
  wire [0:29] sb_1__1__103_chany_top_out;
  wire [0:0] sb_1__1__104_ccff_tail;
  wire [0:29] sb_1__1__104_chanx_left_out;
  wire [0:29] sb_1__1__104_chanx_right_out;
  wire [0:29] sb_1__1__104_chany_bottom_out;
  wire [0:29] sb_1__1__104_chany_top_out;
  wire [0:0] sb_1__1__105_ccff_tail;
  wire [0:29] sb_1__1__105_chanx_left_out;
  wire [0:29] sb_1__1__105_chanx_right_out;
  wire [0:29] sb_1__1__105_chany_bottom_out;
  wire [0:29] sb_1__1__105_chany_top_out;
  wire [0:0] sb_1__1__106_ccff_tail;
  wire [0:29] sb_1__1__106_chanx_left_out;
  wire [0:29] sb_1__1__106_chanx_right_out;
  wire [0:29] sb_1__1__106_chany_bottom_out;
  wire [0:29] sb_1__1__106_chany_top_out;
  wire [0:0] sb_1__1__107_ccff_tail;
  wire [0:29] sb_1__1__107_chanx_left_out;
  wire [0:29] sb_1__1__107_chanx_right_out;
  wire [0:29] sb_1__1__107_chany_bottom_out;
  wire [0:29] sb_1__1__107_chany_top_out;
  wire [0:0] sb_1__1__108_ccff_tail;
  wire [0:29] sb_1__1__108_chanx_left_out;
  wire [0:29] sb_1__1__108_chanx_right_out;
  wire [0:29] sb_1__1__108_chany_bottom_out;
  wire [0:29] sb_1__1__108_chany_top_out;
  wire [0:0] sb_1__1__109_ccff_tail;
  wire [0:29] sb_1__1__109_chanx_left_out;
  wire [0:29] sb_1__1__109_chanx_right_out;
  wire [0:29] sb_1__1__109_chany_bottom_out;
  wire [0:29] sb_1__1__109_chany_top_out;
  wire [0:0] sb_1__1__10_ccff_tail;
  wire [0:29] sb_1__1__10_chanx_left_out;
  wire [0:29] sb_1__1__10_chanx_right_out;
  wire [0:29] sb_1__1__10_chany_bottom_out;
  wire [0:29] sb_1__1__10_chany_top_out;
  wire [0:0] sb_1__1__110_ccff_tail;
  wire [0:29] sb_1__1__110_chanx_left_out;
  wire [0:29] sb_1__1__110_chanx_right_out;
  wire [0:29] sb_1__1__110_chany_bottom_out;
  wire [0:29] sb_1__1__110_chany_top_out;
  wire [0:0] sb_1__1__111_ccff_tail;
  wire [0:29] sb_1__1__111_chanx_left_out;
  wire [0:29] sb_1__1__111_chanx_right_out;
  wire [0:29] sb_1__1__111_chany_bottom_out;
  wire [0:29] sb_1__1__111_chany_top_out;
  wire [0:0] sb_1__1__112_ccff_tail;
  wire [0:29] sb_1__1__112_chanx_left_out;
  wire [0:29] sb_1__1__112_chanx_right_out;
  wire [0:29] sb_1__1__112_chany_bottom_out;
  wire [0:29] sb_1__1__112_chany_top_out;
  wire [0:0] sb_1__1__113_ccff_tail;
  wire [0:29] sb_1__1__113_chanx_left_out;
  wire [0:29] sb_1__1__113_chanx_right_out;
  wire [0:29] sb_1__1__113_chany_bottom_out;
  wire [0:29] sb_1__1__113_chany_top_out;
  wire [0:0] sb_1__1__114_ccff_tail;
  wire [0:29] sb_1__1__114_chanx_left_out;
  wire [0:29] sb_1__1__114_chanx_right_out;
  wire [0:29] sb_1__1__114_chany_bottom_out;
  wire [0:29] sb_1__1__114_chany_top_out;
  wire [0:0] sb_1__1__115_ccff_tail;
  wire [0:29] sb_1__1__115_chanx_left_out;
  wire [0:29] sb_1__1__115_chanx_right_out;
  wire [0:29] sb_1__1__115_chany_bottom_out;
  wire [0:29] sb_1__1__115_chany_top_out;
  wire [0:0] sb_1__1__116_ccff_tail;
  wire [0:29] sb_1__1__116_chanx_left_out;
  wire [0:29] sb_1__1__116_chanx_right_out;
  wire [0:29] sb_1__1__116_chany_bottom_out;
  wire [0:29] sb_1__1__116_chany_top_out;
  wire [0:0] sb_1__1__117_ccff_tail;
  wire [0:29] sb_1__1__117_chanx_left_out;
  wire [0:29] sb_1__1__117_chanx_right_out;
  wire [0:29] sb_1__1__117_chany_bottom_out;
  wire [0:29] sb_1__1__117_chany_top_out;
  wire [0:0] sb_1__1__118_ccff_tail;
  wire [0:29] sb_1__1__118_chanx_left_out;
  wire [0:29] sb_1__1__118_chanx_right_out;
  wire [0:29] sb_1__1__118_chany_bottom_out;
  wire [0:29] sb_1__1__118_chany_top_out;
  wire [0:0] sb_1__1__119_ccff_tail;
  wire [0:29] sb_1__1__119_chanx_left_out;
  wire [0:29] sb_1__1__119_chanx_right_out;
  wire [0:29] sb_1__1__119_chany_bottom_out;
  wire [0:29] sb_1__1__119_chany_top_out;
  wire [0:0] sb_1__1__11_ccff_tail;
  wire [0:29] sb_1__1__11_chanx_left_out;
  wire [0:29] sb_1__1__11_chanx_right_out;
  wire [0:29] sb_1__1__11_chany_bottom_out;
  wire [0:29] sb_1__1__11_chany_top_out;
  wire [0:0] sb_1__1__120_ccff_tail;
  wire [0:29] sb_1__1__120_chanx_left_out;
  wire [0:29] sb_1__1__120_chanx_right_out;
  wire [0:29] sb_1__1__120_chany_bottom_out;
  wire [0:29] sb_1__1__120_chany_top_out;
  wire [0:0] sb_1__1__12_ccff_tail;
  wire [0:29] sb_1__1__12_chanx_left_out;
  wire [0:29] sb_1__1__12_chanx_right_out;
  wire [0:29] sb_1__1__12_chany_bottom_out;
  wire [0:29] sb_1__1__12_chany_top_out;
  wire [0:0] sb_1__1__13_ccff_tail;
  wire [0:29] sb_1__1__13_chanx_left_out;
  wire [0:29] sb_1__1__13_chanx_right_out;
  wire [0:29] sb_1__1__13_chany_bottom_out;
  wire [0:29] sb_1__1__13_chany_top_out;
  wire [0:0] sb_1__1__14_ccff_tail;
  wire [0:29] sb_1__1__14_chanx_left_out;
  wire [0:29] sb_1__1__14_chanx_right_out;
  wire [0:29] sb_1__1__14_chany_bottom_out;
  wire [0:29] sb_1__1__14_chany_top_out;
  wire [0:0] sb_1__1__15_ccff_tail;
  wire [0:29] sb_1__1__15_chanx_left_out;
  wire [0:29] sb_1__1__15_chanx_right_out;
  wire [0:29] sb_1__1__15_chany_bottom_out;
  wire [0:29] sb_1__1__15_chany_top_out;
  wire [0:0] sb_1__1__16_ccff_tail;
  wire [0:29] sb_1__1__16_chanx_left_out;
  wire [0:29] sb_1__1__16_chanx_right_out;
  wire [0:29] sb_1__1__16_chany_bottom_out;
  wire [0:29] sb_1__1__16_chany_top_out;
  wire [0:0] sb_1__1__17_ccff_tail;
  wire [0:29] sb_1__1__17_chanx_left_out;
  wire [0:29] sb_1__1__17_chanx_right_out;
  wire [0:29] sb_1__1__17_chany_bottom_out;
  wire [0:29] sb_1__1__17_chany_top_out;
  wire [0:0] sb_1__1__18_ccff_tail;
  wire [0:29] sb_1__1__18_chanx_left_out;
  wire [0:29] sb_1__1__18_chanx_right_out;
  wire [0:29] sb_1__1__18_chany_bottom_out;
  wire [0:29] sb_1__1__18_chany_top_out;
  wire [0:0] sb_1__1__19_ccff_tail;
  wire [0:29] sb_1__1__19_chanx_left_out;
  wire [0:29] sb_1__1__19_chanx_right_out;
  wire [0:29] sb_1__1__19_chany_bottom_out;
  wire [0:29] sb_1__1__19_chany_top_out;
  wire [0:0] sb_1__1__1_ccff_tail;
  wire [0:29] sb_1__1__1_chanx_left_out;
  wire [0:29] sb_1__1__1_chanx_right_out;
  wire [0:29] sb_1__1__1_chany_bottom_out;
  wire [0:29] sb_1__1__1_chany_top_out;
  wire [0:0] sb_1__1__20_ccff_tail;
  wire [0:29] sb_1__1__20_chanx_left_out;
  wire [0:29] sb_1__1__20_chanx_right_out;
  wire [0:29] sb_1__1__20_chany_bottom_out;
  wire [0:29] sb_1__1__20_chany_top_out;
  wire [0:0] sb_1__1__21_ccff_tail;
  wire [0:29] sb_1__1__21_chanx_left_out;
  wire [0:29] sb_1__1__21_chanx_right_out;
  wire [0:29] sb_1__1__21_chany_bottom_out;
  wire [0:29] sb_1__1__21_chany_top_out;
  wire [0:0] sb_1__1__22_ccff_tail;
  wire [0:29] sb_1__1__22_chanx_left_out;
  wire [0:29] sb_1__1__22_chanx_right_out;
  wire [0:29] sb_1__1__22_chany_bottom_out;
  wire [0:29] sb_1__1__22_chany_top_out;
  wire [0:0] sb_1__1__23_ccff_tail;
  wire [0:29] sb_1__1__23_chanx_left_out;
  wire [0:29] sb_1__1__23_chanx_right_out;
  wire [0:29] sb_1__1__23_chany_bottom_out;
  wire [0:29] sb_1__1__23_chany_top_out;
  wire [0:0] sb_1__1__24_ccff_tail;
  wire [0:29] sb_1__1__24_chanx_left_out;
  wire [0:29] sb_1__1__24_chanx_right_out;
  wire [0:29] sb_1__1__24_chany_bottom_out;
  wire [0:29] sb_1__1__24_chany_top_out;
  wire [0:0] sb_1__1__25_ccff_tail;
  wire [0:29] sb_1__1__25_chanx_left_out;
  wire [0:29] sb_1__1__25_chanx_right_out;
  wire [0:29] sb_1__1__25_chany_bottom_out;
  wire [0:29] sb_1__1__25_chany_top_out;
  wire [0:0] sb_1__1__26_ccff_tail;
  wire [0:29] sb_1__1__26_chanx_left_out;
  wire [0:29] sb_1__1__26_chanx_right_out;
  wire [0:29] sb_1__1__26_chany_bottom_out;
  wire [0:29] sb_1__1__26_chany_top_out;
  wire [0:0] sb_1__1__27_ccff_tail;
  wire [0:29] sb_1__1__27_chanx_left_out;
  wire [0:29] sb_1__1__27_chanx_right_out;
  wire [0:29] sb_1__1__27_chany_bottom_out;
  wire [0:29] sb_1__1__27_chany_top_out;
  wire [0:0] sb_1__1__28_ccff_tail;
  wire [0:29] sb_1__1__28_chanx_left_out;
  wire [0:29] sb_1__1__28_chanx_right_out;
  wire [0:29] sb_1__1__28_chany_bottom_out;
  wire [0:29] sb_1__1__28_chany_top_out;
  wire [0:0] sb_1__1__29_ccff_tail;
  wire [0:29] sb_1__1__29_chanx_left_out;
  wire [0:29] sb_1__1__29_chanx_right_out;
  wire [0:29] sb_1__1__29_chany_bottom_out;
  wire [0:29] sb_1__1__29_chany_top_out;
  wire [0:0] sb_1__1__2_ccff_tail;
  wire [0:29] sb_1__1__2_chanx_left_out;
  wire [0:29] sb_1__1__2_chanx_right_out;
  wire [0:29] sb_1__1__2_chany_bottom_out;
  wire [0:29] sb_1__1__2_chany_top_out;
  wire [0:0] sb_1__1__30_ccff_tail;
  wire [0:29] sb_1__1__30_chanx_left_out;
  wire [0:29] sb_1__1__30_chanx_right_out;
  wire [0:29] sb_1__1__30_chany_bottom_out;
  wire [0:29] sb_1__1__30_chany_top_out;
  wire [0:0] sb_1__1__31_ccff_tail;
  wire [0:29] sb_1__1__31_chanx_left_out;
  wire [0:29] sb_1__1__31_chanx_right_out;
  wire [0:29] sb_1__1__31_chany_bottom_out;
  wire [0:29] sb_1__1__31_chany_top_out;
  wire [0:0] sb_1__1__32_ccff_tail;
  wire [0:29] sb_1__1__32_chanx_left_out;
  wire [0:29] sb_1__1__32_chanx_right_out;
  wire [0:29] sb_1__1__32_chany_bottom_out;
  wire [0:29] sb_1__1__32_chany_top_out;
  wire [0:0] sb_1__1__33_ccff_tail;
  wire [0:29] sb_1__1__33_chanx_left_out;
  wire [0:29] sb_1__1__33_chanx_right_out;
  wire [0:29] sb_1__1__33_chany_bottom_out;
  wire [0:29] sb_1__1__33_chany_top_out;
  wire [0:0] sb_1__1__34_ccff_tail;
  wire [0:29] sb_1__1__34_chanx_left_out;
  wire [0:29] sb_1__1__34_chanx_right_out;
  wire [0:29] sb_1__1__34_chany_bottom_out;
  wire [0:29] sb_1__1__34_chany_top_out;
  wire [0:0] sb_1__1__35_ccff_tail;
  wire [0:29] sb_1__1__35_chanx_left_out;
  wire [0:29] sb_1__1__35_chanx_right_out;
  wire [0:29] sb_1__1__35_chany_bottom_out;
  wire [0:29] sb_1__1__35_chany_top_out;
  wire [0:0] sb_1__1__36_ccff_tail;
  wire [0:29] sb_1__1__36_chanx_left_out;
  wire [0:29] sb_1__1__36_chanx_right_out;
  wire [0:29] sb_1__1__36_chany_bottom_out;
  wire [0:29] sb_1__1__36_chany_top_out;
  wire [0:0] sb_1__1__37_ccff_tail;
  wire [0:29] sb_1__1__37_chanx_left_out;
  wire [0:29] sb_1__1__37_chanx_right_out;
  wire [0:29] sb_1__1__37_chany_bottom_out;
  wire [0:29] sb_1__1__37_chany_top_out;
  wire [0:0] sb_1__1__38_ccff_tail;
  wire [0:29] sb_1__1__38_chanx_left_out;
  wire [0:29] sb_1__1__38_chanx_right_out;
  wire [0:29] sb_1__1__38_chany_bottom_out;
  wire [0:29] sb_1__1__38_chany_top_out;
  wire [0:0] sb_1__1__39_ccff_tail;
  wire [0:29] sb_1__1__39_chanx_left_out;
  wire [0:29] sb_1__1__39_chanx_right_out;
  wire [0:29] sb_1__1__39_chany_bottom_out;
  wire [0:29] sb_1__1__39_chany_top_out;
  wire [0:0] sb_1__1__3_ccff_tail;
  wire [0:29] sb_1__1__3_chanx_left_out;
  wire [0:29] sb_1__1__3_chanx_right_out;
  wire [0:29] sb_1__1__3_chany_bottom_out;
  wire [0:29] sb_1__1__3_chany_top_out;
  wire [0:0] sb_1__1__40_ccff_tail;
  wire [0:29] sb_1__1__40_chanx_left_out;
  wire [0:29] sb_1__1__40_chanx_right_out;
  wire [0:29] sb_1__1__40_chany_bottom_out;
  wire [0:29] sb_1__1__40_chany_top_out;
  wire [0:0] sb_1__1__41_ccff_tail;
  wire [0:29] sb_1__1__41_chanx_left_out;
  wire [0:29] sb_1__1__41_chanx_right_out;
  wire [0:29] sb_1__1__41_chany_bottom_out;
  wire [0:29] sb_1__1__41_chany_top_out;
  wire [0:0] sb_1__1__42_ccff_tail;
  wire [0:29] sb_1__1__42_chanx_left_out;
  wire [0:29] sb_1__1__42_chanx_right_out;
  wire [0:29] sb_1__1__42_chany_bottom_out;
  wire [0:29] sb_1__1__42_chany_top_out;
  wire [0:0] sb_1__1__43_ccff_tail;
  wire [0:29] sb_1__1__43_chanx_left_out;
  wire [0:29] sb_1__1__43_chanx_right_out;
  wire [0:29] sb_1__1__43_chany_bottom_out;
  wire [0:29] sb_1__1__43_chany_top_out;
  wire [0:0] sb_1__1__44_ccff_tail;
  wire [0:29] sb_1__1__44_chanx_left_out;
  wire [0:29] sb_1__1__44_chanx_right_out;
  wire [0:29] sb_1__1__44_chany_bottom_out;
  wire [0:29] sb_1__1__44_chany_top_out;
  wire [0:0] sb_1__1__45_ccff_tail;
  wire [0:29] sb_1__1__45_chanx_left_out;
  wire [0:29] sb_1__1__45_chanx_right_out;
  wire [0:29] sb_1__1__45_chany_bottom_out;
  wire [0:29] sb_1__1__45_chany_top_out;
  wire [0:0] sb_1__1__46_ccff_tail;
  wire [0:29] sb_1__1__46_chanx_left_out;
  wire [0:29] sb_1__1__46_chanx_right_out;
  wire [0:29] sb_1__1__46_chany_bottom_out;
  wire [0:29] sb_1__1__46_chany_top_out;
  wire [0:0] sb_1__1__47_ccff_tail;
  wire [0:29] sb_1__1__47_chanx_left_out;
  wire [0:29] sb_1__1__47_chanx_right_out;
  wire [0:29] sb_1__1__47_chany_bottom_out;
  wire [0:29] sb_1__1__47_chany_top_out;
  wire [0:0] sb_1__1__48_ccff_tail;
  wire [0:29] sb_1__1__48_chanx_left_out;
  wire [0:29] sb_1__1__48_chanx_right_out;
  wire [0:29] sb_1__1__48_chany_bottom_out;
  wire [0:29] sb_1__1__48_chany_top_out;
  wire [0:0] sb_1__1__49_ccff_tail;
  wire [0:29] sb_1__1__49_chanx_left_out;
  wire [0:29] sb_1__1__49_chanx_right_out;
  wire [0:29] sb_1__1__49_chany_bottom_out;
  wire [0:29] sb_1__1__49_chany_top_out;
  wire [0:0] sb_1__1__4_ccff_tail;
  wire [0:29] sb_1__1__4_chanx_left_out;
  wire [0:29] sb_1__1__4_chanx_right_out;
  wire [0:29] sb_1__1__4_chany_bottom_out;
  wire [0:29] sb_1__1__4_chany_top_out;
  wire [0:0] sb_1__1__50_ccff_tail;
  wire [0:29] sb_1__1__50_chanx_left_out;
  wire [0:29] sb_1__1__50_chanx_right_out;
  wire [0:29] sb_1__1__50_chany_bottom_out;
  wire [0:29] sb_1__1__50_chany_top_out;
  wire [0:0] sb_1__1__51_ccff_tail;
  wire [0:29] sb_1__1__51_chanx_left_out;
  wire [0:29] sb_1__1__51_chanx_right_out;
  wire [0:29] sb_1__1__51_chany_bottom_out;
  wire [0:29] sb_1__1__51_chany_top_out;
  wire [0:0] sb_1__1__52_ccff_tail;
  wire [0:29] sb_1__1__52_chanx_left_out;
  wire [0:29] sb_1__1__52_chanx_right_out;
  wire [0:29] sb_1__1__52_chany_bottom_out;
  wire [0:29] sb_1__1__52_chany_top_out;
  wire [0:0] sb_1__1__53_ccff_tail;
  wire [0:29] sb_1__1__53_chanx_left_out;
  wire [0:29] sb_1__1__53_chanx_right_out;
  wire [0:29] sb_1__1__53_chany_bottom_out;
  wire [0:29] sb_1__1__53_chany_top_out;
  wire [0:0] sb_1__1__54_ccff_tail;
  wire [0:29] sb_1__1__54_chanx_left_out;
  wire [0:29] sb_1__1__54_chanx_right_out;
  wire [0:29] sb_1__1__54_chany_bottom_out;
  wire [0:29] sb_1__1__54_chany_top_out;
  wire [0:0] sb_1__1__55_ccff_tail;
  wire [0:29] sb_1__1__55_chanx_left_out;
  wire [0:29] sb_1__1__55_chanx_right_out;
  wire [0:29] sb_1__1__55_chany_bottom_out;
  wire [0:29] sb_1__1__55_chany_top_out;
  wire [0:0] sb_1__1__56_ccff_tail;
  wire [0:29] sb_1__1__56_chanx_left_out;
  wire [0:29] sb_1__1__56_chanx_right_out;
  wire [0:29] sb_1__1__56_chany_bottom_out;
  wire [0:29] sb_1__1__56_chany_top_out;
  wire [0:0] sb_1__1__57_ccff_tail;
  wire [0:29] sb_1__1__57_chanx_left_out;
  wire [0:29] sb_1__1__57_chanx_right_out;
  wire [0:29] sb_1__1__57_chany_bottom_out;
  wire [0:29] sb_1__1__57_chany_top_out;
  wire [0:0] sb_1__1__58_ccff_tail;
  wire [0:29] sb_1__1__58_chanx_left_out;
  wire [0:29] sb_1__1__58_chanx_right_out;
  wire [0:29] sb_1__1__58_chany_bottom_out;
  wire [0:29] sb_1__1__58_chany_top_out;
  wire [0:0] sb_1__1__59_ccff_tail;
  wire [0:29] sb_1__1__59_chanx_left_out;
  wire [0:29] sb_1__1__59_chanx_right_out;
  wire [0:29] sb_1__1__59_chany_bottom_out;
  wire [0:29] sb_1__1__59_chany_top_out;
  wire [0:0] sb_1__1__5_ccff_tail;
  wire [0:29] sb_1__1__5_chanx_left_out;
  wire [0:29] sb_1__1__5_chanx_right_out;
  wire [0:29] sb_1__1__5_chany_bottom_out;
  wire [0:29] sb_1__1__5_chany_top_out;
  wire [0:0] sb_1__1__60_ccff_tail;
  wire [0:29] sb_1__1__60_chanx_left_out;
  wire [0:29] sb_1__1__60_chanx_right_out;
  wire [0:29] sb_1__1__60_chany_bottom_out;
  wire [0:29] sb_1__1__60_chany_top_out;
  wire [0:0] sb_1__1__61_ccff_tail;
  wire [0:29] sb_1__1__61_chanx_left_out;
  wire [0:29] sb_1__1__61_chanx_right_out;
  wire [0:29] sb_1__1__61_chany_bottom_out;
  wire [0:29] sb_1__1__61_chany_top_out;
  wire [0:0] sb_1__1__62_ccff_tail;
  wire [0:29] sb_1__1__62_chanx_left_out;
  wire [0:29] sb_1__1__62_chanx_right_out;
  wire [0:29] sb_1__1__62_chany_bottom_out;
  wire [0:29] sb_1__1__62_chany_top_out;
  wire [0:0] sb_1__1__63_ccff_tail;
  wire [0:29] sb_1__1__63_chanx_left_out;
  wire [0:29] sb_1__1__63_chanx_right_out;
  wire [0:29] sb_1__1__63_chany_bottom_out;
  wire [0:29] sb_1__1__63_chany_top_out;
  wire [0:0] sb_1__1__64_ccff_tail;
  wire [0:29] sb_1__1__64_chanx_left_out;
  wire [0:29] sb_1__1__64_chanx_right_out;
  wire [0:29] sb_1__1__64_chany_bottom_out;
  wire [0:29] sb_1__1__64_chany_top_out;
  wire [0:0] sb_1__1__65_ccff_tail;
  wire [0:29] sb_1__1__65_chanx_left_out;
  wire [0:29] sb_1__1__65_chanx_right_out;
  wire [0:29] sb_1__1__65_chany_bottom_out;
  wire [0:29] sb_1__1__65_chany_top_out;
  wire [0:0] sb_1__1__66_ccff_tail;
  wire [0:29] sb_1__1__66_chanx_left_out;
  wire [0:29] sb_1__1__66_chanx_right_out;
  wire [0:29] sb_1__1__66_chany_bottom_out;
  wire [0:29] sb_1__1__66_chany_top_out;
  wire [0:0] sb_1__1__67_ccff_tail;
  wire [0:29] sb_1__1__67_chanx_left_out;
  wire [0:29] sb_1__1__67_chanx_right_out;
  wire [0:29] sb_1__1__67_chany_bottom_out;
  wire [0:29] sb_1__1__67_chany_top_out;
  wire [0:0] sb_1__1__68_ccff_tail;
  wire [0:29] sb_1__1__68_chanx_left_out;
  wire [0:29] sb_1__1__68_chanx_right_out;
  wire [0:29] sb_1__1__68_chany_bottom_out;
  wire [0:29] sb_1__1__68_chany_top_out;
  wire [0:0] sb_1__1__69_ccff_tail;
  wire [0:29] sb_1__1__69_chanx_left_out;
  wire [0:29] sb_1__1__69_chanx_right_out;
  wire [0:29] sb_1__1__69_chany_bottom_out;
  wire [0:29] sb_1__1__69_chany_top_out;
  wire [0:0] sb_1__1__6_ccff_tail;
  wire [0:29] sb_1__1__6_chanx_left_out;
  wire [0:29] sb_1__1__6_chanx_right_out;
  wire [0:29] sb_1__1__6_chany_bottom_out;
  wire [0:29] sb_1__1__6_chany_top_out;
  wire [0:0] sb_1__1__70_ccff_tail;
  wire [0:29] sb_1__1__70_chanx_left_out;
  wire [0:29] sb_1__1__70_chanx_right_out;
  wire [0:29] sb_1__1__70_chany_bottom_out;
  wire [0:29] sb_1__1__70_chany_top_out;
  wire [0:0] sb_1__1__71_ccff_tail;
  wire [0:29] sb_1__1__71_chanx_left_out;
  wire [0:29] sb_1__1__71_chanx_right_out;
  wire [0:29] sb_1__1__71_chany_bottom_out;
  wire [0:29] sb_1__1__71_chany_top_out;
  wire [0:0] sb_1__1__72_ccff_tail;
  wire [0:29] sb_1__1__72_chanx_left_out;
  wire [0:29] sb_1__1__72_chanx_right_out;
  wire [0:29] sb_1__1__72_chany_bottom_out;
  wire [0:29] sb_1__1__72_chany_top_out;
  wire [0:0] sb_1__1__73_ccff_tail;
  wire [0:29] sb_1__1__73_chanx_left_out;
  wire [0:29] sb_1__1__73_chanx_right_out;
  wire [0:29] sb_1__1__73_chany_bottom_out;
  wire [0:29] sb_1__1__73_chany_top_out;
  wire [0:0] sb_1__1__74_ccff_tail;
  wire [0:29] sb_1__1__74_chanx_left_out;
  wire [0:29] sb_1__1__74_chanx_right_out;
  wire [0:29] sb_1__1__74_chany_bottom_out;
  wire [0:29] sb_1__1__74_chany_top_out;
  wire [0:0] sb_1__1__75_ccff_tail;
  wire [0:29] sb_1__1__75_chanx_left_out;
  wire [0:29] sb_1__1__75_chanx_right_out;
  wire [0:29] sb_1__1__75_chany_bottom_out;
  wire [0:29] sb_1__1__75_chany_top_out;
  wire [0:0] sb_1__1__76_ccff_tail;
  wire [0:29] sb_1__1__76_chanx_left_out;
  wire [0:29] sb_1__1__76_chanx_right_out;
  wire [0:29] sb_1__1__76_chany_bottom_out;
  wire [0:29] sb_1__1__76_chany_top_out;
  wire [0:0] sb_1__1__77_ccff_tail;
  wire [0:29] sb_1__1__77_chanx_left_out;
  wire [0:29] sb_1__1__77_chanx_right_out;
  wire [0:29] sb_1__1__77_chany_bottom_out;
  wire [0:29] sb_1__1__77_chany_top_out;
  wire [0:0] sb_1__1__78_ccff_tail;
  wire [0:29] sb_1__1__78_chanx_left_out;
  wire [0:29] sb_1__1__78_chanx_right_out;
  wire [0:29] sb_1__1__78_chany_bottom_out;
  wire [0:29] sb_1__1__78_chany_top_out;
  wire [0:0] sb_1__1__79_ccff_tail;
  wire [0:29] sb_1__1__79_chanx_left_out;
  wire [0:29] sb_1__1__79_chanx_right_out;
  wire [0:29] sb_1__1__79_chany_bottom_out;
  wire [0:29] sb_1__1__79_chany_top_out;
  wire [0:0] sb_1__1__7_ccff_tail;
  wire [0:29] sb_1__1__7_chanx_left_out;
  wire [0:29] sb_1__1__7_chanx_right_out;
  wire [0:29] sb_1__1__7_chany_bottom_out;
  wire [0:29] sb_1__1__7_chany_top_out;
  wire [0:0] sb_1__1__80_ccff_tail;
  wire [0:29] sb_1__1__80_chanx_left_out;
  wire [0:29] sb_1__1__80_chanx_right_out;
  wire [0:29] sb_1__1__80_chany_bottom_out;
  wire [0:29] sb_1__1__80_chany_top_out;
  wire [0:0] sb_1__1__81_ccff_tail;
  wire [0:29] sb_1__1__81_chanx_left_out;
  wire [0:29] sb_1__1__81_chanx_right_out;
  wire [0:29] sb_1__1__81_chany_bottom_out;
  wire [0:29] sb_1__1__81_chany_top_out;
  wire [0:0] sb_1__1__82_ccff_tail;
  wire [0:29] sb_1__1__82_chanx_left_out;
  wire [0:29] sb_1__1__82_chanx_right_out;
  wire [0:29] sb_1__1__82_chany_bottom_out;
  wire [0:29] sb_1__1__82_chany_top_out;
  wire [0:0] sb_1__1__83_ccff_tail;
  wire [0:29] sb_1__1__83_chanx_left_out;
  wire [0:29] sb_1__1__83_chanx_right_out;
  wire [0:29] sb_1__1__83_chany_bottom_out;
  wire [0:29] sb_1__1__83_chany_top_out;
  wire [0:0] sb_1__1__84_ccff_tail;
  wire [0:29] sb_1__1__84_chanx_left_out;
  wire [0:29] sb_1__1__84_chanx_right_out;
  wire [0:29] sb_1__1__84_chany_bottom_out;
  wire [0:29] sb_1__1__84_chany_top_out;
  wire [0:0] sb_1__1__85_ccff_tail;
  wire [0:29] sb_1__1__85_chanx_left_out;
  wire [0:29] sb_1__1__85_chanx_right_out;
  wire [0:29] sb_1__1__85_chany_bottom_out;
  wire [0:29] sb_1__1__85_chany_top_out;
  wire [0:0] sb_1__1__86_ccff_tail;
  wire [0:29] sb_1__1__86_chanx_left_out;
  wire [0:29] sb_1__1__86_chanx_right_out;
  wire [0:29] sb_1__1__86_chany_bottom_out;
  wire [0:29] sb_1__1__86_chany_top_out;
  wire [0:0] sb_1__1__87_ccff_tail;
  wire [0:29] sb_1__1__87_chanx_left_out;
  wire [0:29] sb_1__1__87_chanx_right_out;
  wire [0:29] sb_1__1__87_chany_bottom_out;
  wire [0:29] sb_1__1__87_chany_top_out;
  wire [0:0] sb_1__1__88_ccff_tail;
  wire [0:29] sb_1__1__88_chanx_left_out;
  wire [0:29] sb_1__1__88_chanx_right_out;
  wire [0:29] sb_1__1__88_chany_bottom_out;
  wire [0:29] sb_1__1__88_chany_top_out;
  wire [0:0] sb_1__1__89_ccff_tail;
  wire [0:29] sb_1__1__89_chanx_left_out;
  wire [0:29] sb_1__1__89_chanx_right_out;
  wire [0:29] sb_1__1__89_chany_bottom_out;
  wire [0:29] sb_1__1__89_chany_top_out;
  wire [0:0] sb_1__1__8_ccff_tail;
  wire [0:29] sb_1__1__8_chanx_left_out;
  wire [0:29] sb_1__1__8_chanx_right_out;
  wire [0:29] sb_1__1__8_chany_bottom_out;
  wire [0:29] sb_1__1__8_chany_top_out;
  wire [0:0] sb_1__1__90_ccff_tail;
  wire [0:29] sb_1__1__90_chanx_left_out;
  wire [0:29] sb_1__1__90_chanx_right_out;
  wire [0:29] sb_1__1__90_chany_bottom_out;
  wire [0:29] sb_1__1__90_chany_top_out;
  wire [0:0] sb_1__1__91_ccff_tail;
  wire [0:29] sb_1__1__91_chanx_left_out;
  wire [0:29] sb_1__1__91_chanx_right_out;
  wire [0:29] sb_1__1__91_chany_bottom_out;
  wire [0:29] sb_1__1__91_chany_top_out;
  wire [0:0] sb_1__1__92_ccff_tail;
  wire [0:29] sb_1__1__92_chanx_left_out;
  wire [0:29] sb_1__1__92_chanx_right_out;
  wire [0:29] sb_1__1__92_chany_bottom_out;
  wire [0:29] sb_1__1__92_chany_top_out;
  wire [0:0] sb_1__1__93_ccff_tail;
  wire [0:29] sb_1__1__93_chanx_left_out;
  wire [0:29] sb_1__1__93_chanx_right_out;
  wire [0:29] sb_1__1__93_chany_bottom_out;
  wire [0:29] sb_1__1__93_chany_top_out;
  wire [0:0] sb_1__1__94_ccff_tail;
  wire [0:29] sb_1__1__94_chanx_left_out;
  wire [0:29] sb_1__1__94_chanx_right_out;
  wire [0:29] sb_1__1__94_chany_bottom_out;
  wire [0:29] sb_1__1__94_chany_top_out;
  wire [0:0] sb_1__1__95_ccff_tail;
  wire [0:29] sb_1__1__95_chanx_left_out;
  wire [0:29] sb_1__1__95_chanx_right_out;
  wire [0:29] sb_1__1__95_chany_bottom_out;
  wire [0:29] sb_1__1__95_chany_top_out;
  wire [0:0] sb_1__1__96_ccff_tail;
  wire [0:29] sb_1__1__96_chanx_left_out;
  wire [0:29] sb_1__1__96_chanx_right_out;
  wire [0:29] sb_1__1__96_chany_bottom_out;
  wire [0:29] sb_1__1__96_chany_top_out;
  wire [0:0] sb_1__1__97_ccff_tail;
  wire [0:29] sb_1__1__97_chanx_left_out;
  wire [0:29] sb_1__1__97_chanx_right_out;
  wire [0:29] sb_1__1__97_chany_bottom_out;
  wire [0:29] sb_1__1__97_chany_top_out;
  wire [0:0] sb_1__1__98_ccff_tail;
  wire [0:29] sb_1__1__98_chanx_left_out;
  wire [0:29] sb_1__1__98_chanx_right_out;
  wire [0:29] sb_1__1__98_chany_bottom_out;
  wire [0:29] sb_1__1__98_chany_top_out;
  wire [0:0] sb_1__1__99_ccff_tail;
  wire [0:29] sb_1__1__99_chanx_left_out;
  wire [0:29] sb_1__1__99_chanx_right_out;
  wire [0:29] sb_1__1__99_chany_bottom_out;
  wire [0:29] sb_1__1__99_chany_top_out;
  wire [0:0] sb_1__1__9_ccff_tail;
  wire [0:29] sb_1__1__9_chanx_left_out;
  wire [0:29] sb_1__1__9_chanx_right_out;
  wire [0:29] sb_1__1__9_chany_bottom_out;
  wire [0:29] sb_1__1__9_chany_top_out;
  wire [1:0] UNCONN;
  wire [317:0] scff_Wires;
  wire [132:0] regin_feedthrough_wires;
  wire [132:0] regout_feedthrough_wires;
  wire [132:0] cin_feedthrough_wires;
  wire [132:0] cout_feedthrough_wires;
  wire [287:0] Test_enWires;
  wire [636:0] pResetWires;
  wire [287:0] ResetWires;
  wire [624:0] prog_clk_0_wires;
  wire [251:0] prog_clk_1_wires;
  wire [135:0] prog_clk_2_wires;
  wire [100:0] prog_clk_3_wires;
  wire [251:0] clk_1_wires;
  wire [135:0] clk_2_wires;
  wire [100:0] clk_3_wires;

  grid_clb
  grid_clb_1__1_
  (
    .clk_0_N_in(clk_1_wires[4]),
    .prog_clk_0_N_in(prog_clk_1_wires[4]),
    .prog_clk_0_W_out(prog_clk_0_wires[3]),
    .prog_clk_0_E_out(prog_clk_0_wires[1]),
    .prog_clk_0_S_out(prog_clk_0_wires[0]),
    .Reset_E_in(ResetWires[24]),
    .pReset_N_in(pResetWires[63]),
    .Test_en_E_in(Test_enWires[24]),
    .SC_OUT_BOT(scff_Wires[25]),
    .SC_IN_TOP(scff_Wires[23]),
    .top_width_0_height_0__pin_0_(cbx_1__1__0_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__0_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__0_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__0_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__0_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__0_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__0_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__0_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__0_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__0_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__0_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__0_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__0_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__0_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__0_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__0_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[0]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__0_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__0_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__0_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__0_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__0_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__0_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__0_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__0_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__0_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__0_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__0_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__0_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__0_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__0_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__0_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__0_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_0_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_0_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_0_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_0_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_0_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_0_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_0_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_0_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_0_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_0_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_0_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_0_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_0_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_0_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_0_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_0_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_0_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_0_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_0_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_0_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_0_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_0_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_0_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_0_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_0_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_0_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_0_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_0_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_0_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_0_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_0_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_0_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_0_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(grid_clb_1__1__undriven_bottom_width_0_height_0__pin_52_[0]),
    .bottom_width_0_height_0__pin_54_(grid_clb_1__1__undriven_bottom_width_0_height_0__pin_54_[0]),
    .ccff_tail(grid_clb_0_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__2_
  (
    .clk_0_S_in(clk_1_wires[3]),
    .prog_clk_0_S_in(prog_clk_1_wires[3]),
    .prog_clk_0_W_out(prog_clk_0_wires[9]),
    .prog_clk_0_E_out(prog_clk_0_wires[7]),
    .prog_clk_0_S_out(prog_clk_0_wires[6]),
    .Reset_E_in(ResetWires[46]),
    .pReset_N_in(pResetWires[112]),
    .Test_en_E_in(Test_enWires[46]),
    .SC_OUT_BOT(scff_Wires[22]),
    .SC_IN_TOP(scff_Wires[21]),
    .top_width_0_height_0__pin_0_(cbx_1__1__1_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__1_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__1_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__1_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__1_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__1_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__1_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__1_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__1_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__1_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__1_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__1_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__1_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__1_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__1_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__1_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[1]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[1]),
    .right_width_0_height_0__pin_16_(cby_1__1__1_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__1_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__1_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__1_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__1_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__1_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__1_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__1_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__1_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__1_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__1_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__1_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__1_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__1_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__1_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__1_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_1_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_1_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_1_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_1_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_1_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_1_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_1_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_1_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_1_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_1_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_1_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_1_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_1_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_1_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_1_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_1_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_1_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_1_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_1_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_1_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_1_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_1_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_1_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_1_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_1_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_1_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_1_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_1_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_1_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_1_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_1_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_1_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_1_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[0]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[0]),
    .ccff_tail(grid_clb_1_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__3_
  (
    .clk_0_N_in(clk_1_wires[11]),
    .prog_clk_0_N_in(prog_clk_1_wires[11]),
    .prog_clk_0_W_out(prog_clk_0_wires[14]),
    .prog_clk_0_E_out(prog_clk_0_wires[12]),
    .prog_clk_0_S_out(prog_clk_0_wires[11]),
    .Reset_E_in(ResetWires[68]),
    .pReset_N_in(pResetWires[161]),
    .Test_en_E_in(Test_enWires[68]),
    .SC_OUT_BOT(scff_Wires[20]),
    .SC_IN_TOP(scff_Wires[19]),
    .top_width_0_height_0__pin_0_(cbx_1__1__2_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__2_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__2_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__2_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__2_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__2_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__2_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__2_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__2_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__2_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__2_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__2_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__2_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__2_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__2_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__2_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[2]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[2]),
    .right_width_0_height_0__pin_16_(cby_1__1__2_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__2_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__2_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__2_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__2_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__2_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__2_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__2_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__2_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__2_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__2_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__2_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__2_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__2_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__2_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__2_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_2_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_2_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_2_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_2_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_2_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_2_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_2_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_2_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_2_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_2_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_2_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_2_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_2_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_2_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_2_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_2_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_2_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_2_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_2_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_2_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_2_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_2_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_2_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_2_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_2_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_2_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_2_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_2_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_2_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_2_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_2_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_2_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_2_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[1]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[1]),
    .ccff_tail(grid_clb_2_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__4_
  (
    .clk_0_S_in(clk_1_wires[10]),
    .prog_clk_0_S_in(prog_clk_1_wires[10]),
    .prog_clk_0_W_out(prog_clk_0_wires[19]),
    .prog_clk_0_E_out(prog_clk_0_wires[17]),
    .prog_clk_0_S_out(prog_clk_0_wires[16]),
    .Reset_E_in(ResetWires[90]),
    .pReset_N_in(pResetWires[210]),
    .Test_en_E_in(Test_enWires[90]),
    .SC_OUT_BOT(scff_Wires[18]),
    .SC_IN_TOP(scff_Wires[17]),
    .top_width_0_height_0__pin_0_(cbx_1__1__3_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__3_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__3_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__3_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__3_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__3_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__3_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__3_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__3_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__3_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__3_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__3_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__3_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__3_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__3_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__3_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[3]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[3]),
    .right_width_0_height_0__pin_16_(cby_1__1__3_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__3_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__3_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__3_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__3_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__3_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__3_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__3_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__3_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__3_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__3_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__3_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__3_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__3_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__3_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__3_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_3_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_3_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_3_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_3_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_3_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_3_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_3_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_3_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_3_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_3_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_3_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_3_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_3_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_3_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_3_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_3_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_3_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_3_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_3_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_3_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_3_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_3_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_3_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_3_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_3_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_3_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_3_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_3_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_3_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_3_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_3_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_3_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_3_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[2]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[2]),
    .ccff_tail(grid_clb_3_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__5_
  (
    .clk_0_N_in(clk_1_wires[18]),
    .prog_clk_0_N_in(prog_clk_1_wires[18]),
    .prog_clk_0_W_out(prog_clk_0_wires[24]),
    .prog_clk_0_E_out(prog_clk_0_wires[22]),
    .prog_clk_0_S_out(prog_clk_0_wires[21]),
    .Reset_E_in(ResetWires[112]),
    .pReset_N_in(pResetWires[259]),
    .Test_en_E_in(Test_enWires[112]),
    .SC_OUT_BOT(scff_Wires[16]),
    .SC_IN_TOP(scff_Wires[15]),
    .top_width_0_height_0__pin_0_(cbx_1__1__4_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__4_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__4_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__4_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__4_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__4_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__4_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__4_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__4_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__4_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__4_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__4_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__4_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__4_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__4_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__4_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[4]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[4]),
    .right_width_0_height_0__pin_16_(cby_1__1__4_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__4_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__4_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__4_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__4_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__4_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__4_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__4_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__4_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__4_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__4_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__4_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__4_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__4_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__4_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__4_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_4_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_4_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_4_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_4_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_4_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_4_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_4_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_4_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_4_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_4_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_4_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_4_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_4_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_4_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_4_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_4_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_4_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_4_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_4_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_4_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_4_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_4_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_4_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_4_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_4_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_4_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_4_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_4_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_4_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_4_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_4_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_4_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_4_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[3]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[3]),
    .ccff_tail(grid_clb_4_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__6_
  (
    .clk_0_S_in(clk_1_wires[17]),
    .prog_clk_0_S_in(prog_clk_1_wires[17]),
    .prog_clk_0_W_out(prog_clk_0_wires[29]),
    .prog_clk_0_E_out(prog_clk_0_wires[27]),
    .prog_clk_0_S_out(prog_clk_0_wires[26]),
    .Reset_E_in(ResetWires[134]),
    .pReset_N_in(pResetWires[308]),
    .Test_en_E_in(Test_enWires[134]),
    .SC_OUT_BOT(scff_Wires[14]),
    .SC_IN_TOP(scff_Wires[13]),
    .top_width_0_height_0__pin_0_(cbx_1__1__5_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__5_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__5_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__5_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__5_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__5_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__5_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__5_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__5_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__5_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__5_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__5_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__5_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__5_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__5_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__5_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[5]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[5]),
    .right_width_0_height_0__pin_16_(cby_1__1__5_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__5_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__5_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__5_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__5_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__5_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__5_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__5_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__5_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__5_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__5_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__5_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__5_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__5_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__5_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__5_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_5_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_5_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_5_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_5_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_5_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_5_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_5_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_5_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_5_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_5_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_5_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_5_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_5_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_5_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_5_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_5_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_5_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_5_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_5_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_5_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_5_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_5_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_5_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_5_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_5_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_5_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_5_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_5_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_5_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_5_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_5_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_5_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_5_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[4]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[4]),
    .ccff_tail(grid_clb_5_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__7_
  (
    .clk_0_N_in(clk_1_wires[25]),
    .prog_clk_0_N_in(prog_clk_1_wires[25]),
    .prog_clk_0_W_out(prog_clk_0_wires[34]),
    .prog_clk_0_E_out(prog_clk_0_wires[32]),
    .prog_clk_0_S_out(prog_clk_0_wires[31]),
    .Reset_E_in(ResetWires[156]),
    .pReset_N_in(pResetWires[357]),
    .Test_en_E_in(Test_enWires[156]),
    .SC_OUT_BOT(scff_Wires[12]),
    .SC_IN_TOP(scff_Wires[11]),
    .top_width_0_height_0__pin_0_(cbx_1__1__6_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__6_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__6_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__6_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__6_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__6_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__6_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__6_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__6_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__6_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__6_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__6_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__6_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__6_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__6_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__6_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[6]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[6]),
    .right_width_0_height_0__pin_16_(cby_1__1__6_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__6_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__6_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__6_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__6_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__6_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__6_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__6_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__6_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__6_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__6_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__6_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__6_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__6_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__6_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__6_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_6_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_6_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_6_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_6_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_6_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_6_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_6_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_6_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_6_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_6_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_6_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_6_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_6_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_6_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_6_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_6_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_6_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_6_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_6_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_6_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_6_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_6_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_6_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_6_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_6_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_6_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_6_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_6_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_6_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_6_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_6_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_6_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_6_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[5]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[5]),
    .ccff_tail(grid_clb_6_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__8_
  (
    .clk_0_S_in(clk_1_wires[24]),
    .prog_clk_0_S_in(prog_clk_1_wires[24]),
    .prog_clk_0_W_out(prog_clk_0_wires[39]),
    .prog_clk_0_E_out(prog_clk_0_wires[37]),
    .prog_clk_0_S_out(prog_clk_0_wires[36]),
    .Reset_E_in(ResetWires[178]),
    .pReset_N_in(pResetWires[406]),
    .Test_en_E_in(Test_enWires[178]),
    .SC_OUT_BOT(scff_Wires[10]),
    .SC_IN_TOP(scff_Wires[9]),
    .top_width_0_height_0__pin_0_(cbx_1__1__7_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__7_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__7_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__7_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__7_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__7_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__7_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__7_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__7_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__7_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__7_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__7_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__7_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__7_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__7_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__7_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[7]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[7]),
    .right_width_0_height_0__pin_16_(cby_1__1__7_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__7_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__7_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__7_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__7_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__7_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__7_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__7_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__7_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__7_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__7_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__7_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__7_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__7_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__7_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__7_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_7_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_7_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_7_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_7_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_7_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_7_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_7_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_7_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_7_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_7_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_7_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_7_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_7_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_7_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_7_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_7_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_7_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_7_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_7_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_7_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_7_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_7_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_7_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_7_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_7_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_7_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_7_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_7_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_7_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_7_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_7_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_7_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_7_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[6]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[6]),
    .ccff_tail(grid_clb_7_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__9_
  (
    .clk_0_N_in(clk_1_wires[32]),
    .prog_clk_0_N_in(prog_clk_1_wires[32]),
    .prog_clk_0_W_out(prog_clk_0_wires[44]),
    .prog_clk_0_E_out(prog_clk_0_wires[42]),
    .prog_clk_0_S_out(prog_clk_0_wires[41]),
    .Reset_E_in(ResetWires[200]),
    .pReset_N_in(pResetWires[455]),
    .Test_en_E_in(Test_enWires[200]),
    .SC_OUT_BOT(scff_Wires[8]),
    .SC_IN_TOP(scff_Wires[7]),
    .top_width_0_height_0__pin_0_(cbx_1__1__8_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__8_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__8_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__8_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__8_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__8_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__8_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__8_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__8_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__8_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__8_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__8_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__8_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__8_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__8_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__8_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[8]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[8]),
    .right_width_0_height_0__pin_16_(cby_1__1__8_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__8_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__8_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__8_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__8_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__8_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__8_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__8_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__8_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__8_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__8_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__8_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__8_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__8_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__8_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__8_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_8_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_8_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_8_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_8_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_8_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_8_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_8_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_8_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_8_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_8_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_8_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_8_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_8_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_8_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_8_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_8_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_8_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_8_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_8_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_8_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_8_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_8_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_8_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_8_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_8_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_8_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_8_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_8_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_8_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_8_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_8_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_8_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_8_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[7]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[7]),
    .ccff_tail(grid_clb_8_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__10_
  (
    .clk_0_S_in(clk_1_wires[31]),
    .prog_clk_0_S_in(prog_clk_1_wires[31]),
    .prog_clk_0_W_out(prog_clk_0_wires[49]),
    .prog_clk_0_E_out(prog_clk_0_wires[47]),
    .prog_clk_0_S_out(prog_clk_0_wires[46]),
    .Reset_E_in(ResetWires[222]),
    .pReset_N_in(pResetWires[504]),
    .Test_en_E_in(Test_enWires[222]),
    .SC_OUT_BOT(scff_Wires[6]),
    .SC_IN_TOP(scff_Wires[5]),
    .top_width_0_height_0__pin_0_(cbx_1__1__9_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__9_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__9_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__9_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__9_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__9_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__9_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__9_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__9_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__9_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__9_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__9_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__9_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__9_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__9_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__9_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[9]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[9]),
    .right_width_0_height_0__pin_16_(cby_1__1__9_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__9_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__9_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__9_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__9_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__9_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__9_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__9_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__9_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__9_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__9_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__9_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__9_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__9_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__9_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__9_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_9_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_9_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_9_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_9_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_9_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_9_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_9_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_9_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_9_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_9_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_9_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_9_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_9_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_9_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_9_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_9_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_9_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_9_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_9_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_9_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_9_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_9_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_9_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_9_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_9_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_9_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_9_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_9_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_9_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_9_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_9_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_9_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_9_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[8]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[8]),
    .ccff_tail(grid_clb_9_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__11_
  (
    .clk_0_N_in(clk_1_wires[39]),
    .prog_clk_0_N_in(prog_clk_1_wires[39]),
    .prog_clk_0_W_out(prog_clk_0_wires[54]),
    .prog_clk_0_E_out(prog_clk_0_wires[52]),
    .prog_clk_0_S_out(prog_clk_0_wires[51]),
    .Reset_E_in(ResetWires[244]),
    .pReset_N_in(pResetWires[553]),
    .Test_en_E_in(Test_enWires[244]),
    .SC_OUT_BOT(scff_Wires[4]),
    .SC_IN_TOP(scff_Wires[3]),
    .top_width_0_height_0__pin_0_(cbx_1__1__10_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__10_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__10_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__10_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__10_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__10_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__10_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__10_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__10_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__10_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__10_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__10_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__10_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__10_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__10_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__10_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[10]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[10]),
    .right_width_0_height_0__pin_16_(cby_1__1__10_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__10_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__10_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__10_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__10_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__10_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__10_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__10_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__10_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__10_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__10_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__10_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__10_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__10_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__10_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__10_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_10_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_10_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_10_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_10_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_10_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_10_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_10_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_10_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_10_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_10_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_10_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_10_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_10_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_10_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_10_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_10_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_10_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_10_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_10_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_10_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_10_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_10_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_10_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_10_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_10_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_10_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_10_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_10_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_10_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_10_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_10_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_10_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_10_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[9]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[9]),
    .ccff_tail(grid_clb_10_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__12_
  (
    .clk_0_S_in(clk_1_wires[38]),
    .prog_clk_0_S_in(prog_clk_1_wires[38]),
    .prog_clk_0_W_out(prog_clk_0_wires[61]),
    .prog_clk_0_N_out(prog_clk_0_wires[59]),
    .prog_clk_0_E_out(prog_clk_0_wires[57]),
    .prog_clk_0_S_out(prog_clk_0_wires[56]),
    .Reset_E_in(ResetWires[266]),
    .pReset_N_in(pResetWires[602]),
    .Test_en_E_in(Test_enWires[266]),
    .SC_OUT_BOT(scff_Wires[2]),
    .SC_IN_TOP(scff_Wires[1]),
    .top_width_0_height_0__pin_0_(cbx_1__12__0_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__0_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__0_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__0_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__0_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__0_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__0_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__0_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__0_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__0_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__0_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__0_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__0_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__0_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__0_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__0_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_1__12__undriven_top_width_0_height_0__pin_32_[0]),
    .top_width_0_height_0__pin_34_(grid_clb_1__12__undriven_top_width_0_height_0__pin_34_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__11_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__11_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__11_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__11_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__11_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__11_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__11_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__11_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__11_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__11_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__11_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__11_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__11_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__11_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__11_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__11_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_11_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_11_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_11_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_11_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_11_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_11_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_11_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_11_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_11_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_11_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_11_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_11_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_11_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_11_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_11_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_11_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_11_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_11_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_11_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_11_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_11_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_11_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_11_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_11_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_11_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_11_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_11_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_11_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_11_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_11_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_11_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_11_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_11_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[10]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[10]),
    .ccff_tail(grid_clb_11_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__1_
  (
    .clk_0_N_in(clk_1_wires[6]),
    .prog_clk_0_N_in(prog_clk_1_wires[6]),
    .prog_clk_0_E_out(prog_clk_0_wires[64]),
    .prog_clk_0_S_out(prog_clk_0_wires[63]),
    .Reset_W_out(ResetWires[26]),
    .Reset_E_in(ResetWires[25]),
    .pReset_N_in(pResetWires[68]),
    .Test_en_W_out(Test_enWires[26]),
    .Test_en_E_in(Test_enWires[25]),
    .SC_OUT_TOP(scff_Wires[29]),
    .SC_IN_BOT(scff_Wires[28]),
    .top_width_0_height_0__pin_0_(cbx_1__1__11_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__11_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__11_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__11_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__11_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__11_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__11_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__11_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__11_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__11_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__11_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__11_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__11_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__11_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__11_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__11_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[11]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[11]),
    .right_width_0_height_0__pin_16_(cby_1__1__12_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__12_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__12_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__12_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__12_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__12_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__12_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__12_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__12_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__12_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__12_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__12_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__12_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__12_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__12_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__12_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__0_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_12_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_12_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_12_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_12_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_12_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_12_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_12_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_12_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_12_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_12_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_12_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_12_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_12_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_12_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_12_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_12_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_12_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_12_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_12_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_12_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_12_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_12_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_12_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_12_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_12_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_12_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_12_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_12_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_12_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_12_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_12_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_12_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(grid_clb_2__1__undriven_bottom_width_0_height_0__pin_52_[0]),
    .bottom_width_0_height_0__pin_54_(grid_clb_2__1__undriven_bottom_width_0_height_0__pin_54_[0]),
    .ccff_tail(grid_clb_12_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__2_
  (
    .clk_0_S_in(clk_1_wires[5]),
    .prog_clk_0_S_in(prog_clk_1_wires[5]),
    .prog_clk_0_E_out(prog_clk_0_wires[67]),
    .prog_clk_0_S_out(prog_clk_0_wires[66]),
    .Reset_W_out(ResetWires[48]),
    .Reset_E_in(ResetWires[47]),
    .pReset_N_in(pResetWires[117]),
    .Test_en_W_out(Test_enWires[48]),
    .Test_en_E_in(Test_enWires[47]),
    .SC_OUT_TOP(scff_Wires[31]),
    .SC_IN_BOT(scff_Wires[30]),
    .top_width_0_height_0__pin_0_(cbx_1__1__12_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__12_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__12_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__12_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__12_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__12_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__12_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__12_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__12_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__12_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__12_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__12_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__12_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__12_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__12_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__12_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[12]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[12]),
    .right_width_0_height_0__pin_16_(cby_1__1__13_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__13_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__13_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__13_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__13_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__13_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__13_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__13_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__13_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__13_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__13_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__13_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__13_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__13_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__13_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__13_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__1_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_13_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_13_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_13_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_13_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_13_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_13_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_13_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_13_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_13_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_13_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_13_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_13_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_13_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_13_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_13_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_13_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_13_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_13_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_13_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_13_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_13_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_13_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_13_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_13_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_13_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_13_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_13_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_13_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_13_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_13_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_13_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_13_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[11]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[11]),
    .ccff_tail(grid_clb_13_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__3_
  (
    .clk_0_N_in(clk_1_wires[13]),
    .prog_clk_0_N_in(prog_clk_1_wires[13]),
    .prog_clk_0_E_out(prog_clk_0_wires[70]),
    .prog_clk_0_S_out(prog_clk_0_wires[69]),
    .Reset_W_out(ResetWires[70]),
    .Reset_E_in(ResetWires[69]),
    .pReset_N_in(pResetWires[166]),
    .Test_en_W_out(Test_enWires[70]),
    .Test_en_E_in(Test_enWires[69]),
    .SC_OUT_TOP(scff_Wires[33]),
    .SC_IN_BOT(scff_Wires[32]),
    .top_width_0_height_0__pin_0_(cbx_1__1__13_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__13_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__13_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__13_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__13_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__13_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__13_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__13_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__13_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__13_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__13_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__13_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__13_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__13_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__13_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__13_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[13]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[13]),
    .right_width_0_height_0__pin_16_(cby_1__1__14_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__14_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__14_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__14_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__14_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__14_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__14_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__14_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__14_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__14_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__14_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__14_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__14_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__14_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__14_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__14_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__2_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_14_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_14_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_14_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_14_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_14_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_14_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_14_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_14_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_14_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_14_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_14_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_14_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_14_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_14_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_14_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_14_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_14_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_14_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_14_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_14_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_14_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_14_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_14_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_14_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_14_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_14_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_14_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_14_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_14_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_14_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_14_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_14_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[12]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[12]),
    .ccff_tail(grid_clb_14_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__4_
  (
    .clk_0_S_in(clk_1_wires[12]),
    .prog_clk_0_S_in(prog_clk_1_wires[12]),
    .prog_clk_0_E_out(prog_clk_0_wires[73]),
    .prog_clk_0_S_out(prog_clk_0_wires[72]),
    .Reset_W_out(ResetWires[92]),
    .Reset_E_in(ResetWires[91]),
    .pReset_N_in(pResetWires[215]),
    .Test_en_W_out(Test_enWires[92]),
    .Test_en_E_in(Test_enWires[91]),
    .SC_OUT_TOP(scff_Wires[35]),
    .SC_IN_BOT(scff_Wires[34]),
    .top_width_0_height_0__pin_0_(cbx_1__1__14_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__14_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__14_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__14_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__14_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__14_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__14_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__14_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__14_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__14_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__14_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__14_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__14_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__14_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__14_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__14_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[14]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[14]),
    .right_width_0_height_0__pin_16_(cby_1__1__15_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__15_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__15_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__15_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__15_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__15_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__15_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__15_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__15_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__15_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__15_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__15_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__15_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__15_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__15_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__15_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__3_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_15_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_15_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_15_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_15_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_15_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_15_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_15_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_15_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_15_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_15_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_15_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_15_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_15_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_15_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_15_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_15_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_15_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_15_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_15_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_15_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_15_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_15_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_15_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_15_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_15_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_15_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_15_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_15_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_15_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_15_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_15_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_15_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[13]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[13]),
    .ccff_tail(grid_clb_15_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__5_
  (
    .clk_0_N_in(clk_1_wires[20]),
    .prog_clk_0_N_in(prog_clk_1_wires[20]),
    .prog_clk_0_E_out(prog_clk_0_wires[76]),
    .prog_clk_0_S_out(prog_clk_0_wires[75]),
    .Reset_W_out(ResetWires[114]),
    .Reset_E_in(ResetWires[113]),
    .pReset_N_in(pResetWires[264]),
    .Test_en_W_out(Test_enWires[114]),
    .Test_en_E_in(Test_enWires[113]),
    .SC_OUT_TOP(scff_Wires[37]),
    .SC_IN_BOT(scff_Wires[36]),
    .top_width_0_height_0__pin_0_(cbx_1__1__15_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__15_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__15_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__15_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__15_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__15_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__15_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__15_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__15_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__15_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__15_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__15_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__15_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__15_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__15_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__15_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[15]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[15]),
    .right_width_0_height_0__pin_16_(cby_1__1__16_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__16_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__16_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__16_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__16_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__16_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__16_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__16_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__16_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__16_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__16_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__16_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__16_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__16_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__16_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__16_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__4_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_16_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_16_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_16_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_16_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_16_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_16_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_16_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_16_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_16_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_16_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_16_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_16_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_16_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_16_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_16_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_16_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_16_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_16_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_16_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_16_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_16_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_16_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_16_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_16_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_16_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_16_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_16_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_16_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_16_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_16_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_16_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_16_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[14]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[14]),
    .ccff_tail(grid_clb_16_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__6_
  (
    .clk_0_S_in(clk_1_wires[19]),
    .prog_clk_0_S_in(prog_clk_1_wires[19]),
    .prog_clk_0_E_out(prog_clk_0_wires[79]),
    .prog_clk_0_S_out(prog_clk_0_wires[78]),
    .Reset_W_out(ResetWires[136]),
    .Reset_E_in(ResetWires[135]),
    .pReset_N_in(pResetWires[313]),
    .Test_en_W_out(Test_enWires[136]),
    .Test_en_E_in(Test_enWires[135]),
    .SC_OUT_TOP(scff_Wires[39]),
    .SC_IN_BOT(scff_Wires[38]),
    .top_width_0_height_0__pin_0_(cbx_1__1__16_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__16_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__16_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__16_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__16_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__16_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__16_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__16_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__16_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__16_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__16_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__16_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__16_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__16_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__16_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__16_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[16]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[16]),
    .right_width_0_height_0__pin_16_(cby_1__1__17_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__17_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__17_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__17_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__17_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__17_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__17_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__17_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__17_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__17_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__17_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__17_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__17_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__17_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__17_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__17_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__5_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_17_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_17_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_17_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_17_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_17_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_17_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_17_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_17_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_17_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_17_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_17_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_17_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_17_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_17_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_17_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_17_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_17_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_17_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_17_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_17_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_17_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_17_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_17_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_17_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_17_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_17_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_17_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_17_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_17_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_17_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_17_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_17_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[15]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[15]),
    .ccff_tail(grid_clb_17_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__7_
  (
    .clk_0_N_in(clk_1_wires[27]),
    .prog_clk_0_N_in(prog_clk_1_wires[27]),
    .prog_clk_0_E_out(prog_clk_0_wires[82]),
    .prog_clk_0_S_out(prog_clk_0_wires[81]),
    .Reset_W_out(ResetWires[158]),
    .Reset_E_in(ResetWires[157]),
    .pReset_N_in(pResetWires[362]),
    .Test_en_W_out(Test_enWires[158]),
    .Test_en_E_in(Test_enWires[157]),
    .SC_OUT_TOP(scff_Wires[41]),
    .SC_IN_BOT(scff_Wires[40]),
    .top_width_0_height_0__pin_0_(cbx_1__1__17_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__17_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__17_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__17_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__17_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__17_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__17_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__17_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__17_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__17_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__17_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__17_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__17_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__17_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__17_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__17_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[17]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[17]),
    .right_width_0_height_0__pin_16_(cby_1__1__18_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__18_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__18_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__18_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__18_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__18_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__18_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__18_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__18_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__18_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__18_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__18_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__18_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__18_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__18_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__18_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__6_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_18_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_18_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_18_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_18_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_18_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_18_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_18_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_18_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_18_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_18_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_18_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_18_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_18_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_18_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_18_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_18_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_18_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_18_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_18_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_18_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_18_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_18_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_18_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_18_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_18_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_18_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_18_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_18_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_18_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_18_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_18_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_18_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[16]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[16]),
    .ccff_tail(grid_clb_18_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__8_
  (
    .clk_0_S_in(clk_1_wires[26]),
    .prog_clk_0_S_in(prog_clk_1_wires[26]),
    .prog_clk_0_E_out(prog_clk_0_wires[85]),
    .prog_clk_0_S_out(prog_clk_0_wires[84]),
    .Reset_W_out(ResetWires[180]),
    .Reset_E_in(ResetWires[179]),
    .pReset_N_in(pResetWires[411]),
    .Test_en_W_out(Test_enWires[180]),
    .Test_en_E_in(Test_enWires[179]),
    .SC_OUT_TOP(scff_Wires[43]),
    .SC_IN_BOT(scff_Wires[42]),
    .top_width_0_height_0__pin_0_(cbx_1__1__18_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__18_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__18_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__18_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__18_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__18_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__18_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__18_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__18_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__18_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__18_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__18_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__18_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__18_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__18_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__18_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[18]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[18]),
    .right_width_0_height_0__pin_16_(cby_1__1__19_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__19_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__19_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__19_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__19_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__19_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__19_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__19_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__19_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__19_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__19_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__19_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__19_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__19_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__19_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__19_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__7_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_19_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_19_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_19_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_19_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_19_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_19_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_19_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_19_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_19_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_19_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_19_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_19_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_19_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_19_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_19_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_19_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_19_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_19_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_19_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_19_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_19_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_19_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_19_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_19_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_19_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_19_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_19_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_19_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_19_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_19_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_19_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_19_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[17]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[17]),
    .ccff_tail(grid_clb_19_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__9_
  (
    .clk_0_N_in(clk_1_wires[34]),
    .prog_clk_0_N_in(prog_clk_1_wires[34]),
    .prog_clk_0_E_out(prog_clk_0_wires[88]),
    .prog_clk_0_S_out(prog_clk_0_wires[87]),
    .Reset_W_out(ResetWires[202]),
    .Reset_E_in(ResetWires[201]),
    .pReset_N_in(pResetWires[460]),
    .Test_en_W_out(Test_enWires[202]),
    .Test_en_E_in(Test_enWires[201]),
    .SC_OUT_TOP(scff_Wires[45]),
    .SC_IN_BOT(scff_Wires[44]),
    .top_width_0_height_0__pin_0_(cbx_1__1__19_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__19_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__19_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__19_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__19_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__19_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__19_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__19_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__19_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__19_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__19_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__19_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__19_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__19_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__19_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__19_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[19]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[19]),
    .right_width_0_height_0__pin_16_(cby_1__1__20_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__20_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__20_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__20_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__20_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__20_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__20_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__20_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__20_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__20_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__20_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__20_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__20_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__20_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__20_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__20_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__8_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_20_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_20_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_20_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_20_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_20_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_20_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_20_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_20_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_20_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_20_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_20_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_20_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_20_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_20_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_20_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_20_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_20_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_20_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_20_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_20_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_20_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_20_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_20_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_20_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_20_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_20_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_20_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_20_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_20_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_20_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_20_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_20_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[18]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[18]),
    .ccff_tail(grid_clb_20_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__10_
  (
    .clk_0_S_in(clk_1_wires[33]),
    .prog_clk_0_S_in(prog_clk_1_wires[33]),
    .prog_clk_0_E_out(prog_clk_0_wires[91]),
    .prog_clk_0_S_out(prog_clk_0_wires[90]),
    .Reset_W_out(ResetWires[224]),
    .Reset_E_in(ResetWires[223]),
    .pReset_N_in(pResetWires[509]),
    .Test_en_W_out(Test_enWires[224]),
    .Test_en_E_in(Test_enWires[223]),
    .SC_OUT_TOP(scff_Wires[47]),
    .SC_IN_BOT(scff_Wires[46]),
    .top_width_0_height_0__pin_0_(cbx_1__1__20_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__20_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__20_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__20_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__20_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__20_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__20_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__20_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__20_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__20_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__20_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__20_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__20_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__20_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__20_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__20_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[20]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[20]),
    .right_width_0_height_0__pin_16_(cby_1__1__21_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__21_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__21_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__21_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__21_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__21_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__21_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__21_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__21_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__21_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__21_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__21_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__21_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__21_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__21_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__21_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__9_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_21_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_21_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_21_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_21_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_21_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_21_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_21_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_21_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_21_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_21_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_21_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_21_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_21_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_21_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_21_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_21_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_21_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_21_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_21_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_21_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_21_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_21_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_21_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_21_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_21_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_21_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_21_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_21_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_21_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_21_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_21_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_21_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[19]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[19]),
    .ccff_tail(grid_clb_21_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__11_
  (
    .clk_0_N_in(clk_1_wires[41]),
    .prog_clk_0_N_in(prog_clk_1_wires[41]),
    .prog_clk_0_E_out(prog_clk_0_wires[94]),
    .prog_clk_0_S_out(prog_clk_0_wires[93]),
    .Reset_W_out(ResetWires[246]),
    .Reset_E_in(ResetWires[245]),
    .pReset_N_in(pResetWires[558]),
    .Test_en_W_out(Test_enWires[246]),
    .Test_en_E_in(Test_enWires[245]),
    .SC_OUT_TOP(scff_Wires[49]),
    .SC_IN_BOT(scff_Wires[48]),
    .top_width_0_height_0__pin_0_(cbx_1__1__21_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__21_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__21_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__21_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__21_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__21_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__21_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__21_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__21_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__21_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__21_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__21_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__21_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__21_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__21_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__21_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[21]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[21]),
    .right_width_0_height_0__pin_16_(cby_1__1__22_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__22_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__22_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__22_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__22_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__22_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__22_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__22_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__22_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__22_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__22_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__22_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__22_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__22_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__22_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__22_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__10_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_22_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_22_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_22_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_22_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_22_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_22_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_22_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_22_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_22_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_22_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_22_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_22_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_22_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_22_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_22_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_22_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_22_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_22_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_22_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_22_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_22_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_22_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_22_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_22_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_22_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_22_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_22_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_22_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_22_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_22_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_22_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_22_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[20]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[20]),
    .ccff_tail(grid_clb_22_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__12_
  (
    .clk_0_S_in(clk_1_wires[40]),
    .prog_clk_0_S_in(prog_clk_1_wires[40]),
    .prog_clk_0_N_out(prog_clk_0_wires[99]),
    .prog_clk_0_E_out(prog_clk_0_wires[97]),
    .prog_clk_0_S_out(prog_clk_0_wires[96]),
    .Reset_W_out(ResetWires[268]),
    .Reset_E_in(ResetWires[267]),
    .pReset_N_in(pResetWires[606]),
    .Test_en_W_out(Test_enWires[268]),
    .Test_en_E_in(Test_enWires[267]),
    .SC_OUT_TOP(scff_Wires[51]),
    .SC_IN_BOT(scff_Wires[50]),
    .top_width_0_height_0__pin_0_(cbx_1__12__1_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__1_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__1_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__1_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__1_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__1_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__1_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__1_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__1_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__1_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__1_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__1_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__1_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__1_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__1_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__1_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_2__12__undriven_top_width_0_height_0__pin_32_[0]),
    .top_width_0_height_0__pin_34_(grid_clb_2__12__undriven_top_width_0_height_0__pin_34_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__23_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__23_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__23_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__23_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__23_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__23_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__23_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__23_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__23_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__23_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__23_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__23_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__23_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__23_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__23_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__23_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__11_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_23_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_23_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_23_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_23_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_23_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_23_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_23_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_23_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_23_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_23_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_23_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_23_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_23_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_23_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_23_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_23_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_23_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_23_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_23_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_23_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_23_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_23_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_23_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_23_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_23_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_23_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_23_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_23_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_23_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_23_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_23_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_23_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[21]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[21]),
    .ccff_tail(grid_clb_23_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__1_
  (
    .clk_0_N_in(clk_1_wires[46]),
    .prog_clk_0_N_in(prog_clk_1_wires[46]),
    .prog_clk_0_E_out(prog_clk_0_wires[102]),
    .prog_clk_0_S_out(prog_clk_0_wires[101]),
    .Reset_W_out(ResetWires[28]),
    .Reset_E_in(ResetWires[27]),
    .pReset_N_in(pResetWires[72]),
    .Test_en_W_out(Test_enWires[28]),
    .Test_en_E_in(Test_enWires[27]),
    .SC_OUT_BOT(scff_Wires[78]),
    .SC_IN_TOP(scff_Wires[76]),
    .top_width_0_height_0__pin_0_(cbx_1__1__22_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__22_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__22_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__22_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__22_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__22_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__22_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__22_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__22_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__22_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__22_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__22_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__22_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__22_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__22_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__22_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[22]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[22]),
    .right_width_0_height_0__pin_16_(cby_1__1__24_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__24_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__24_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__24_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__24_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__24_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__24_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__24_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__24_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__24_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__24_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__24_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__24_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__24_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__24_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__24_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__12_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_24_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_24_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_24_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_24_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_24_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_24_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_24_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_24_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_24_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_24_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_24_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_24_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_24_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_24_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_24_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_24_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_24_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_24_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_24_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_24_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_24_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_24_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_24_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_24_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_24_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_24_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_24_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_24_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_24_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_24_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_24_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_24_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(grid_clb_3__1__undriven_bottom_width_0_height_0__pin_52_[0]),
    .bottom_width_0_height_0__pin_54_(grid_clb_3__1__undriven_bottom_width_0_height_0__pin_54_[0]),
    .ccff_tail(grid_clb_24_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__2_
  (
    .clk_0_S_in(clk_1_wires[45]),
    .prog_clk_0_S_in(prog_clk_1_wires[45]),
    .prog_clk_0_E_out(prog_clk_0_wires[105]),
    .prog_clk_0_S_out(prog_clk_0_wires[104]),
    .Reset_W_out(ResetWires[50]),
    .Reset_E_in(ResetWires[49]),
    .pReset_N_in(pResetWires[121]),
    .Test_en_W_out(Test_enWires[50]),
    .Test_en_E_in(Test_enWires[49]),
    .SC_OUT_BOT(scff_Wires[75]),
    .SC_IN_TOP(scff_Wires[74]),
    .top_width_0_height_0__pin_0_(cbx_1__1__23_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__23_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__23_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__23_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__23_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__23_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__23_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__23_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__23_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__23_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__23_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__23_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__23_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__23_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__23_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__23_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[23]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[23]),
    .right_width_0_height_0__pin_16_(cby_1__1__25_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__25_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__25_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__25_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__25_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__25_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__25_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__25_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__25_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__25_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__25_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__25_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__25_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__25_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__25_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__25_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__13_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_25_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_25_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_25_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_25_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_25_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_25_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_25_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_25_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_25_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_25_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_25_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_25_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_25_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_25_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_25_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_25_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_25_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_25_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_25_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_25_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_25_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_25_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_25_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_25_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_25_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_25_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_25_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_25_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_25_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_25_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_25_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_25_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[22]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[22]),
    .ccff_tail(grid_clb_25_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__3_
  (
    .clk_0_N_in(clk_1_wires[53]),
    .prog_clk_0_N_in(prog_clk_1_wires[53]),
    .prog_clk_0_E_out(prog_clk_0_wires[108]),
    .prog_clk_0_S_out(prog_clk_0_wires[107]),
    .Reset_W_out(ResetWires[72]),
    .Reset_E_in(ResetWires[71]),
    .pReset_N_in(pResetWires[170]),
    .Test_en_W_out(Test_enWires[72]),
    .Test_en_E_in(Test_enWires[71]),
    .SC_OUT_BOT(scff_Wires[73]),
    .SC_IN_TOP(scff_Wires[72]),
    .top_width_0_height_0__pin_0_(cbx_1__1__24_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__24_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__24_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__24_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__24_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__24_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__24_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__24_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__24_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__24_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__24_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__24_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__24_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__24_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__24_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__24_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[24]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[24]),
    .right_width_0_height_0__pin_16_(cby_1__1__26_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__26_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__26_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__26_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__26_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__26_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__26_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__26_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__26_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__26_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__26_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__26_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__26_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__26_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__26_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__26_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__14_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_26_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_26_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_26_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_26_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_26_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_26_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_26_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_26_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_26_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_26_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_26_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_26_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_26_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_26_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_26_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_26_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_26_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_26_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_26_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_26_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_26_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_26_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_26_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_26_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_26_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_26_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_26_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_26_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_26_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_26_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_26_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_26_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[23]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[23]),
    .ccff_tail(grid_clb_26_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__4_
  (
    .clk_0_S_in(clk_1_wires[52]),
    .prog_clk_0_S_in(prog_clk_1_wires[52]),
    .prog_clk_0_E_out(prog_clk_0_wires[111]),
    .prog_clk_0_S_out(prog_clk_0_wires[110]),
    .Reset_W_out(ResetWires[94]),
    .Reset_E_in(ResetWires[93]),
    .pReset_N_in(pResetWires[219]),
    .Test_en_W_out(Test_enWires[94]),
    .Test_en_E_in(Test_enWires[93]),
    .SC_OUT_BOT(scff_Wires[71]),
    .SC_IN_TOP(scff_Wires[70]),
    .top_width_0_height_0__pin_0_(cbx_1__1__25_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__25_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__25_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__25_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__25_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__25_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__25_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__25_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__25_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__25_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__25_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__25_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__25_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__25_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__25_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__25_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[25]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[25]),
    .right_width_0_height_0__pin_16_(cby_1__1__27_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__27_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__27_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__27_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__27_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__27_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__27_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__27_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__27_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__27_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__27_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__27_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__27_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__27_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__27_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__27_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__15_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_27_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_27_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_27_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_27_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_27_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_27_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_27_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_27_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_27_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_27_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_27_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_27_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_27_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_27_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_27_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_27_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_27_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_27_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_27_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_27_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_27_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_27_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_27_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_27_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_27_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_27_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_27_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_27_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_27_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_27_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_27_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_27_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[24]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[24]),
    .ccff_tail(grid_clb_27_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__5_
  (
    .clk_0_N_in(clk_1_wires[60]),
    .prog_clk_0_N_in(prog_clk_1_wires[60]),
    .prog_clk_0_E_out(prog_clk_0_wires[114]),
    .prog_clk_0_S_out(prog_clk_0_wires[113]),
    .Reset_W_out(ResetWires[116]),
    .Reset_E_in(ResetWires[115]),
    .pReset_N_in(pResetWires[268]),
    .Test_en_W_out(Test_enWires[116]),
    .Test_en_E_in(Test_enWires[115]),
    .SC_OUT_BOT(scff_Wires[69]),
    .SC_IN_TOP(scff_Wires[68]),
    .top_width_0_height_0__pin_0_(cbx_1__1__26_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__26_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__26_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__26_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__26_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__26_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__26_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__26_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__26_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__26_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__26_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__26_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__26_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__26_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__26_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__26_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[26]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[26]),
    .right_width_0_height_0__pin_16_(cby_1__1__28_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__28_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__28_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__28_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__28_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__28_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__28_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__28_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__28_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__28_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__28_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__28_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__28_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__28_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__28_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__28_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__16_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_28_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_28_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_28_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_28_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_28_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_28_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_28_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_28_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_28_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_28_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_28_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_28_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_28_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_28_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_28_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_28_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_28_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_28_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_28_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_28_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_28_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_28_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_28_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_28_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_28_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_28_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_28_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_28_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_28_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_28_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_28_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_28_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[25]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[25]),
    .ccff_tail(grid_clb_28_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__6_
  (
    .clk_0_S_in(clk_1_wires[59]),
    .prog_clk_0_S_in(prog_clk_1_wires[59]),
    .prog_clk_0_E_out(prog_clk_0_wires[117]),
    .prog_clk_0_S_out(prog_clk_0_wires[116]),
    .Reset_W_out(ResetWires[138]),
    .Reset_E_in(ResetWires[137]),
    .pReset_N_in(pResetWires[317]),
    .Test_en_W_out(Test_enWires[138]),
    .Test_en_E_in(Test_enWires[137]),
    .SC_OUT_BOT(scff_Wires[67]),
    .SC_IN_TOP(scff_Wires[66]),
    .top_width_0_height_0__pin_0_(cbx_1__1__27_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__27_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__27_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__27_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__27_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__27_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__27_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__27_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__27_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__27_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__27_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__27_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__27_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__27_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__27_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__27_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[27]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[27]),
    .right_width_0_height_0__pin_16_(cby_1__1__29_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__29_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__29_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__29_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__29_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__29_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__29_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__29_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__29_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__29_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__29_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__29_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__29_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__29_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__29_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__29_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__17_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_29_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_29_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_29_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_29_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_29_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_29_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_29_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_29_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_29_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_29_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_29_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_29_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_29_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_29_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_29_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_29_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_29_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_29_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_29_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_29_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_29_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_29_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_29_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_29_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_29_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_29_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_29_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_29_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_29_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_29_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_29_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_29_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[26]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[26]),
    .ccff_tail(grid_clb_29_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__7_
  (
    .clk_0_N_in(clk_1_wires[67]),
    .prog_clk_0_N_in(prog_clk_1_wires[67]),
    .prog_clk_0_E_out(prog_clk_0_wires[120]),
    .prog_clk_0_S_out(prog_clk_0_wires[119]),
    .Reset_W_out(ResetWires[160]),
    .Reset_E_in(ResetWires[159]),
    .pReset_N_in(pResetWires[366]),
    .Test_en_W_out(Test_enWires[160]),
    .Test_en_E_in(Test_enWires[159]),
    .SC_OUT_BOT(scff_Wires[65]),
    .SC_IN_TOP(scff_Wires[64]),
    .top_width_0_height_0__pin_0_(cbx_1__1__28_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__28_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__28_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__28_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__28_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__28_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__28_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__28_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__28_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__28_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__28_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__28_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__28_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__28_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__28_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__28_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[28]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[28]),
    .right_width_0_height_0__pin_16_(cby_1__1__30_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__30_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__30_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__30_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__30_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__30_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__30_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__30_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__30_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__30_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__30_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__30_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__30_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__30_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__30_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__30_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__18_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_30_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_30_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_30_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_30_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_30_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_30_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_30_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_30_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_30_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_30_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_30_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_30_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_30_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_30_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_30_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_30_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_30_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_30_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_30_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_30_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_30_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_30_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_30_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_30_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_30_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_30_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_30_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_30_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_30_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_30_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_30_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_30_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[27]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[27]),
    .ccff_tail(grid_clb_30_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__8_
  (
    .clk_0_S_in(clk_1_wires[66]),
    .prog_clk_0_S_in(prog_clk_1_wires[66]),
    .prog_clk_0_E_out(prog_clk_0_wires[123]),
    .prog_clk_0_S_out(prog_clk_0_wires[122]),
    .Reset_W_out(ResetWires[182]),
    .Reset_E_in(ResetWires[181]),
    .pReset_N_in(pResetWires[415]),
    .Test_en_W_out(Test_enWires[182]),
    .Test_en_E_in(Test_enWires[181]),
    .SC_OUT_BOT(scff_Wires[63]),
    .SC_IN_TOP(scff_Wires[62]),
    .top_width_0_height_0__pin_0_(cbx_1__1__29_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__29_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__29_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__29_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__29_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__29_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__29_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__29_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__29_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__29_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__29_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__29_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__29_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__29_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__29_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__29_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[29]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[29]),
    .right_width_0_height_0__pin_16_(cby_1__1__31_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__31_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__31_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__31_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__31_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__31_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__31_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__31_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__31_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__31_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__31_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__31_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__31_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__31_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__31_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__31_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__19_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_31_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_31_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_31_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_31_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_31_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_31_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_31_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_31_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_31_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_31_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_31_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_31_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_31_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_31_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_31_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_31_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_31_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_31_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_31_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_31_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_31_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_31_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_31_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_31_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_31_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_31_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_31_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_31_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_31_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_31_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_31_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_31_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[28]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[28]),
    .ccff_tail(grid_clb_31_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__9_
  (
    .clk_0_N_in(clk_1_wires[74]),
    .prog_clk_0_N_in(prog_clk_1_wires[74]),
    .prog_clk_0_E_out(prog_clk_0_wires[126]),
    .prog_clk_0_S_out(prog_clk_0_wires[125]),
    .Reset_W_out(ResetWires[204]),
    .Reset_E_in(ResetWires[203]),
    .pReset_N_in(pResetWires[464]),
    .Test_en_W_out(Test_enWires[204]),
    .Test_en_E_in(Test_enWires[203]),
    .SC_OUT_BOT(scff_Wires[61]),
    .SC_IN_TOP(scff_Wires[60]),
    .top_width_0_height_0__pin_0_(cbx_1__1__30_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__30_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__30_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__30_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__30_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__30_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__30_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__30_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__30_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__30_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__30_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__30_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__30_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__30_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__30_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__30_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[30]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[30]),
    .right_width_0_height_0__pin_16_(cby_1__1__32_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__32_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__32_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__32_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__32_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__32_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__32_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__32_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__32_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__32_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__32_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__32_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__32_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__32_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__32_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__32_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__20_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_32_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_32_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_32_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_32_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_32_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_32_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_32_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_32_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_32_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_32_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_32_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_32_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_32_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_32_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_32_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_32_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_32_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_32_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_32_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_32_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_32_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_32_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_32_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_32_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_32_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_32_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_32_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_32_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_32_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_32_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_32_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_32_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[29]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[29]),
    .ccff_tail(grid_clb_32_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__10_
  (
    .clk_0_S_in(clk_1_wires[73]),
    .prog_clk_0_S_in(prog_clk_1_wires[73]),
    .prog_clk_0_E_out(prog_clk_0_wires[129]),
    .prog_clk_0_S_out(prog_clk_0_wires[128]),
    .Reset_W_out(ResetWires[226]),
    .Reset_E_in(ResetWires[225]),
    .pReset_N_in(pResetWires[513]),
    .Test_en_W_out(Test_enWires[226]),
    .Test_en_E_in(Test_enWires[225]),
    .SC_OUT_BOT(scff_Wires[59]),
    .SC_IN_TOP(scff_Wires[58]),
    .top_width_0_height_0__pin_0_(cbx_1__1__31_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__31_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__31_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__31_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__31_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__31_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__31_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__31_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__31_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__31_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__31_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__31_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__31_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__31_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__31_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__31_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[31]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[31]),
    .right_width_0_height_0__pin_16_(cby_1__1__33_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__33_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__33_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__33_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__33_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__33_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__33_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__33_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__33_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__33_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__33_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__33_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__33_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__33_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__33_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__33_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__21_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_33_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_33_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_33_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_33_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_33_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_33_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_33_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_33_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_33_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_33_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_33_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_33_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_33_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_33_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_33_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_33_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_33_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_33_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_33_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_33_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_33_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_33_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_33_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_33_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_33_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_33_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_33_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_33_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_33_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_33_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_33_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_33_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[30]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[30]),
    .ccff_tail(grid_clb_33_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__11_
  (
    .clk_0_N_in(clk_1_wires[81]),
    .prog_clk_0_N_in(prog_clk_1_wires[81]),
    .prog_clk_0_E_out(prog_clk_0_wires[132]),
    .prog_clk_0_S_out(prog_clk_0_wires[131]),
    .Reset_W_out(ResetWires[248]),
    .Reset_E_in(ResetWires[247]),
    .pReset_N_in(pResetWires[562]),
    .Test_en_W_out(Test_enWires[248]),
    .Test_en_E_in(Test_enWires[247]),
    .SC_OUT_BOT(scff_Wires[57]),
    .SC_IN_TOP(scff_Wires[56]),
    .top_width_0_height_0__pin_0_(cbx_1__1__32_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__32_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__32_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__32_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__32_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__32_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__32_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__32_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__32_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__32_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__32_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__32_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__32_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__32_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__32_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__32_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[32]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[32]),
    .right_width_0_height_0__pin_16_(cby_1__1__34_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__34_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__34_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__34_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__34_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__34_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__34_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__34_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__34_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__34_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__34_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__34_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__34_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__34_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__34_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__34_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__22_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_34_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_34_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_34_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_34_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_34_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_34_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_34_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_34_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_34_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_34_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_34_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_34_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_34_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_34_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_34_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_34_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_34_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_34_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_34_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_34_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_34_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_34_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_34_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_34_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_34_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_34_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_34_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_34_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_34_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_34_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_34_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_34_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[31]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[31]),
    .ccff_tail(grid_clb_34_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__12_
  (
    .clk_0_S_in(clk_1_wires[80]),
    .prog_clk_0_S_in(prog_clk_1_wires[80]),
    .prog_clk_0_N_out(prog_clk_0_wires[137]),
    .prog_clk_0_E_out(prog_clk_0_wires[135]),
    .prog_clk_0_S_out(prog_clk_0_wires[134]),
    .Reset_W_out(ResetWires[270]),
    .Reset_E_in(ResetWires[269]),
    .pReset_N_in(pResetWires[609]),
    .Test_en_W_out(Test_enWires[270]),
    .Test_en_E_in(Test_enWires[269]),
    .SC_OUT_BOT(scff_Wires[55]),
    .SC_IN_TOP(scff_Wires[54]),
    .top_width_0_height_0__pin_0_(cbx_1__12__2_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__2_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__2_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__2_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__2_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__2_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__2_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__2_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__2_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__2_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__2_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__2_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__2_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__2_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__2_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__2_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_3__12__undriven_top_width_0_height_0__pin_32_[0]),
    .top_width_0_height_0__pin_34_(grid_clb_3__12__undriven_top_width_0_height_0__pin_34_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__35_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__35_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__35_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__35_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__35_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__35_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__35_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__35_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__35_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__35_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__35_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__35_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__35_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__35_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__35_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__35_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__23_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_35_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_35_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_35_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_35_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_35_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_35_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_35_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_35_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_35_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_35_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_35_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_35_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_35_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_35_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_35_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_35_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_35_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_35_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_35_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_35_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_35_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_35_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_35_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_35_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_35_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_35_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_35_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_35_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_35_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_35_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_35_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_35_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[32]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[32]),
    .ccff_tail(grid_clb_35_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__1_
  (
    .clk_0_N_in(clk_1_wires[48]),
    .prog_clk_0_N_in(prog_clk_1_wires[48]),
    .prog_clk_0_E_out(prog_clk_0_wires[140]),
    .prog_clk_0_S_out(prog_clk_0_wires[139]),
    .Reset_W_out(ResetWires[30]),
    .Reset_E_in(ResetWires[29]),
    .pReset_N_in(pResetWires[76]),
    .Test_en_W_out(Test_enWires[30]),
    .Test_en_E_in(Test_enWires[29]),
    .SC_OUT_TOP(scff_Wires[82]),
    .SC_IN_BOT(scff_Wires[81]),
    .top_width_0_height_0__pin_0_(cbx_1__1__33_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__33_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__33_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__33_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__33_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__33_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__33_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__33_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__33_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__33_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__33_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__33_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__33_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__33_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__33_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__33_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[33]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[33]),
    .right_width_0_height_0__pin_16_(cby_1__1__36_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__36_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__36_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__36_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__36_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__36_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__36_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__36_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__36_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__36_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__36_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__36_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__36_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__36_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__36_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__36_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__24_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_36_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_36_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_36_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_36_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_36_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_36_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_36_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_36_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_36_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_36_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_36_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_36_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_36_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_36_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_36_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_36_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_36_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_36_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_36_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_36_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_36_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_36_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_36_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_36_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_36_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_36_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_36_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_36_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_36_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_36_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_36_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_36_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(grid_clb_4__1__undriven_bottom_width_0_height_0__pin_52_[0]),
    .bottom_width_0_height_0__pin_54_(grid_clb_4__1__undriven_bottom_width_0_height_0__pin_54_[0]),
    .ccff_tail(grid_clb_36_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__2_
  (
    .clk_0_S_in(clk_1_wires[47]),
    .prog_clk_0_S_in(prog_clk_1_wires[47]),
    .prog_clk_0_E_out(prog_clk_0_wires[143]),
    .prog_clk_0_S_out(prog_clk_0_wires[142]),
    .Reset_W_out(ResetWires[52]),
    .Reset_E_in(ResetWires[51]),
    .pReset_N_in(pResetWires[125]),
    .Test_en_W_out(Test_enWires[52]),
    .Test_en_E_in(Test_enWires[51]),
    .SC_OUT_TOP(scff_Wires[84]),
    .SC_IN_BOT(scff_Wires[83]),
    .top_width_0_height_0__pin_0_(cbx_1__1__34_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__34_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__34_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__34_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__34_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__34_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__34_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__34_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__34_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__34_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__34_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__34_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__34_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__34_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__34_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__34_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[34]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[34]),
    .right_width_0_height_0__pin_16_(cby_1__1__37_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__37_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__37_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__37_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__37_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__37_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__37_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__37_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__37_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__37_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__37_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__37_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__37_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__37_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__37_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__37_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__25_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_37_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_37_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_37_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_37_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_37_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_37_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_37_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_37_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_37_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_37_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_37_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_37_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_37_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_37_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_37_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_37_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_37_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_37_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_37_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_37_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_37_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_37_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_37_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_37_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_37_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_37_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_37_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_37_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_37_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_37_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_37_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_37_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[33]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[33]),
    .ccff_tail(grid_clb_37_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__3_
  (
    .clk_0_N_in(clk_1_wires[55]),
    .prog_clk_0_N_in(prog_clk_1_wires[55]),
    .prog_clk_0_E_out(prog_clk_0_wires[146]),
    .prog_clk_0_S_out(prog_clk_0_wires[145]),
    .Reset_W_out(ResetWires[74]),
    .Reset_E_in(ResetWires[73]),
    .pReset_N_in(pResetWires[174]),
    .Test_en_W_out(Test_enWires[74]),
    .Test_en_E_in(Test_enWires[73]),
    .SC_OUT_TOP(scff_Wires[86]),
    .SC_IN_BOT(scff_Wires[85]),
    .top_width_0_height_0__pin_0_(cbx_1__1__35_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__35_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__35_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__35_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__35_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__35_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__35_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__35_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__35_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__35_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__35_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__35_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__35_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__35_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__35_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__35_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[35]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[35]),
    .right_width_0_height_0__pin_16_(cby_1__1__38_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__38_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__38_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__38_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__38_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__38_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__38_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__38_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__38_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__38_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__38_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__38_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__38_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__38_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__38_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__38_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__26_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_38_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_38_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_38_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_38_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_38_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_38_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_38_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_38_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_38_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_38_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_38_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_38_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_38_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_38_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_38_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_38_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_38_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_38_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_38_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_38_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_38_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_38_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_38_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_38_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_38_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_38_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_38_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_38_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_38_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_38_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_38_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_38_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[34]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[34]),
    .ccff_tail(grid_clb_38_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__4_
  (
    .clk_0_S_in(clk_1_wires[54]),
    .prog_clk_0_S_in(prog_clk_1_wires[54]),
    .prog_clk_0_E_out(prog_clk_0_wires[149]),
    .prog_clk_0_S_out(prog_clk_0_wires[148]),
    .Reset_W_out(ResetWires[96]),
    .Reset_E_in(ResetWires[95]),
    .pReset_N_in(pResetWires[223]),
    .Test_en_W_out(Test_enWires[96]),
    .Test_en_E_in(Test_enWires[95]),
    .SC_OUT_TOP(scff_Wires[88]),
    .SC_IN_BOT(scff_Wires[87]),
    .top_width_0_height_0__pin_0_(cbx_1__1__36_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__36_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__36_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__36_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__36_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__36_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__36_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__36_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__36_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__36_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__36_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__36_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__36_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__36_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__36_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__36_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[36]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[36]),
    .right_width_0_height_0__pin_16_(cby_1__1__39_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__39_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__39_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__39_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__39_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__39_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__39_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__39_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__39_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__39_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__39_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__39_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__39_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__39_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__39_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__39_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__27_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_39_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_39_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_39_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_39_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_39_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_39_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_39_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_39_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_39_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_39_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_39_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_39_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_39_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_39_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_39_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_39_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_39_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_39_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_39_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_39_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_39_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_39_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_39_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_39_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_39_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_39_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_39_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_39_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_39_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_39_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_39_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_39_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[35]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[35]),
    .ccff_tail(grid_clb_39_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__5_
  (
    .clk_0_N_in(clk_1_wires[62]),
    .prog_clk_0_N_in(prog_clk_1_wires[62]),
    .prog_clk_0_E_out(prog_clk_0_wires[152]),
    .prog_clk_0_S_out(prog_clk_0_wires[151]),
    .Reset_W_out(ResetWires[118]),
    .Reset_E_in(ResetWires[117]),
    .pReset_N_in(pResetWires[272]),
    .Test_en_W_out(Test_enWires[118]),
    .Test_en_E_in(Test_enWires[117]),
    .SC_OUT_TOP(scff_Wires[90]),
    .SC_IN_BOT(scff_Wires[89]),
    .top_width_0_height_0__pin_0_(cbx_1__1__37_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__37_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__37_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__37_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__37_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__37_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__37_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__37_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__37_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__37_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__37_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__37_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__37_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__37_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__37_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__37_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[37]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[37]),
    .right_width_0_height_0__pin_16_(cby_1__1__40_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__40_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__40_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__40_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__40_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__40_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__40_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__40_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__40_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__40_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__40_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__40_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__40_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__40_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__40_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__40_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__28_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_40_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_40_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_40_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_40_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_40_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_40_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_40_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_40_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_40_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_40_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_40_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_40_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_40_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_40_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_40_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_40_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_40_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_40_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_40_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_40_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_40_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_40_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_40_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_40_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_40_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_40_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_40_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_40_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_40_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_40_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_40_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_40_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[36]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[36]),
    .ccff_tail(grid_clb_40_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__6_
  (
    .clk_0_S_in(clk_1_wires[61]),
    .prog_clk_0_S_in(prog_clk_1_wires[61]),
    .prog_clk_0_E_out(prog_clk_0_wires[155]),
    .prog_clk_0_S_out(prog_clk_0_wires[154]),
    .Reset_W_out(ResetWires[140]),
    .Reset_E_in(ResetWires[139]),
    .pReset_N_in(pResetWires[321]),
    .Test_en_W_out(Test_enWires[140]),
    .Test_en_E_in(Test_enWires[139]),
    .SC_OUT_TOP(scff_Wires[92]),
    .SC_IN_BOT(scff_Wires[91]),
    .top_width_0_height_0__pin_0_(cbx_1__1__38_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__38_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__38_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__38_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__38_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__38_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__38_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__38_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__38_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__38_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__38_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__38_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__38_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__38_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__38_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__38_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[38]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[38]),
    .right_width_0_height_0__pin_16_(cby_1__1__41_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__41_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__41_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__41_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__41_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__41_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__41_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__41_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__41_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__41_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__41_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__41_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__41_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__41_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__41_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__41_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__29_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_41_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_41_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_41_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_41_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_41_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_41_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_41_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_41_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_41_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_41_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_41_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_41_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_41_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_41_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_41_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_41_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_41_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_41_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_41_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_41_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_41_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_41_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_41_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_41_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_41_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_41_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_41_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_41_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_41_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_41_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_41_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_41_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[37]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[37]),
    .ccff_tail(grid_clb_41_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__7_
  (
    .clk_0_N_in(clk_1_wires[69]),
    .prog_clk_0_N_in(prog_clk_1_wires[69]),
    .prog_clk_0_E_out(prog_clk_0_wires[158]),
    .prog_clk_0_S_out(prog_clk_0_wires[157]),
    .Reset_W_out(ResetWires[162]),
    .Reset_E_in(ResetWires[161]),
    .pReset_N_in(pResetWires[370]),
    .Test_en_W_out(Test_enWires[162]),
    .Test_en_E_in(Test_enWires[161]),
    .SC_OUT_TOP(scff_Wires[94]),
    .SC_IN_BOT(scff_Wires[93]),
    .top_width_0_height_0__pin_0_(cbx_1__1__39_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__39_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__39_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__39_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__39_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__39_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__39_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__39_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__39_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__39_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__39_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__39_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__39_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__39_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__39_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__39_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[39]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[39]),
    .right_width_0_height_0__pin_16_(cby_1__1__42_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__42_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__42_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__42_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__42_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__42_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__42_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__42_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__42_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__42_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__42_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__42_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__42_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__42_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__42_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__42_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__30_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_42_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_42_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_42_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_42_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_42_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_42_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_42_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_42_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_42_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_42_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_42_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_42_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_42_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_42_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_42_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_42_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_42_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_42_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_42_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_42_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_42_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_42_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_42_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_42_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_42_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_42_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_42_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_42_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_42_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_42_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_42_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_42_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[38]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[38]),
    .ccff_tail(grid_clb_42_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__8_
  (
    .clk_0_S_in(clk_1_wires[68]),
    .prog_clk_0_S_in(prog_clk_1_wires[68]),
    .prog_clk_0_E_out(prog_clk_0_wires[161]),
    .prog_clk_0_S_out(prog_clk_0_wires[160]),
    .Reset_W_out(ResetWires[184]),
    .Reset_E_in(ResetWires[183]),
    .pReset_N_in(pResetWires[419]),
    .Test_en_W_out(Test_enWires[184]),
    .Test_en_E_in(Test_enWires[183]),
    .SC_OUT_TOP(scff_Wires[96]),
    .SC_IN_BOT(scff_Wires[95]),
    .top_width_0_height_0__pin_0_(cbx_1__1__40_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__40_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__40_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__40_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__40_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__40_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__40_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__40_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__40_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__40_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__40_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__40_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__40_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__40_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__40_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__40_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[40]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[40]),
    .right_width_0_height_0__pin_16_(cby_1__1__43_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__43_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__43_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__43_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__43_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__43_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__43_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__43_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__43_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__43_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__43_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__43_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__43_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__43_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__43_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__43_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__31_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_43_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_43_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_43_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_43_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_43_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_43_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_43_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_43_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_43_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_43_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_43_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_43_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_43_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_43_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_43_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_43_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_43_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_43_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_43_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_43_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_43_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_43_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_43_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_43_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_43_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_43_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_43_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_43_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_43_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_43_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_43_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_43_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[39]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[39]),
    .ccff_tail(grid_clb_43_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__9_
  (
    .clk_0_N_in(clk_1_wires[76]),
    .prog_clk_0_N_in(prog_clk_1_wires[76]),
    .prog_clk_0_E_out(prog_clk_0_wires[164]),
    .prog_clk_0_S_out(prog_clk_0_wires[163]),
    .Reset_W_out(ResetWires[206]),
    .Reset_E_in(ResetWires[205]),
    .pReset_N_in(pResetWires[468]),
    .Test_en_W_out(Test_enWires[206]),
    .Test_en_E_in(Test_enWires[205]),
    .SC_OUT_TOP(scff_Wires[98]),
    .SC_IN_BOT(scff_Wires[97]),
    .top_width_0_height_0__pin_0_(cbx_1__1__41_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__41_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__41_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__41_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__41_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__41_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__41_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__41_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__41_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__41_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__41_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__41_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__41_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__41_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__41_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__41_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[41]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[41]),
    .right_width_0_height_0__pin_16_(cby_1__1__44_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__44_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__44_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__44_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__44_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__44_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__44_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__44_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__44_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__44_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__44_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__44_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__44_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__44_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__44_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__44_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__32_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_44_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_44_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_44_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_44_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_44_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_44_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_44_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_44_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_44_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_44_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_44_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_44_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_44_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_44_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_44_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_44_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_44_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_44_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_44_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_44_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_44_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_44_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_44_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_44_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_44_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_44_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_44_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_44_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_44_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_44_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_44_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_44_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[40]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[40]),
    .ccff_tail(grid_clb_44_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__10_
  (
    .clk_0_S_in(clk_1_wires[75]),
    .prog_clk_0_S_in(prog_clk_1_wires[75]),
    .prog_clk_0_E_out(prog_clk_0_wires[167]),
    .prog_clk_0_S_out(prog_clk_0_wires[166]),
    .Reset_W_out(ResetWires[228]),
    .Reset_E_in(ResetWires[227]),
    .pReset_N_in(pResetWires[517]),
    .Test_en_W_out(Test_enWires[228]),
    .Test_en_E_in(Test_enWires[227]),
    .SC_OUT_TOP(scff_Wires[100]),
    .SC_IN_BOT(scff_Wires[99]),
    .top_width_0_height_0__pin_0_(cbx_1__1__42_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__42_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__42_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__42_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__42_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__42_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__42_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__42_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__42_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__42_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__42_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__42_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__42_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__42_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__42_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__42_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[42]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[42]),
    .right_width_0_height_0__pin_16_(cby_1__1__45_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__45_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__45_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__45_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__45_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__45_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__45_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__45_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__45_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__45_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__45_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__45_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__45_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__45_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__45_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__45_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__33_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_45_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_45_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_45_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_45_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_45_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_45_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_45_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_45_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_45_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_45_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_45_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_45_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_45_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_45_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_45_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_45_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_45_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_45_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_45_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_45_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_45_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_45_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_45_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_45_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_45_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_45_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_45_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_45_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_45_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_45_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_45_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_45_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[41]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[41]),
    .ccff_tail(grid_clb_45_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__11_
  (
    .clk_0_N_in(clk_1_wires[83]),
    .prog_clk_0_N_in(prog_clk_1_wires[83]),
    .prog_clk_0_E_out(prog_clk_0_wires[170]),
    .prog_clk_0_S_out(prog_clk_0_wires[169]),
    .Reset_W_out(ResetWires[250]),
    .Reset_E_in(ResetWires[249]),
    .pReset_N_in(pResetWires[566]),
    .Test_en_W_out(Test_enWires[250]),
    .Test_en_E_in(Test_enWires[249]),
    .SC_OUT_TOP(scff_Wires[102]),
    .SC_IN_BOT(scff_Wires[101]),
    .top_width_0_height_0__pin_0_(cbx_1__1__43_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__43_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__43_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__43_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__43_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__43_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__43_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__43_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__43_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__43_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__43_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__43_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__43_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__43_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__43_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__43_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[43]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[43]),
    .right_width_0_height_0__pin_16_(cby_1__1__46_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__46_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__46_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__46_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__46_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__46_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__46_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__46_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__46_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__46_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__46_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__46_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__46_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__46_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__46_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__46_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__34_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_46_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_46_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_46_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_46_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_46_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_46_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_46_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_46_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_46_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_46_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_46_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_46_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_46_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_46_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_46_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_46_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_46_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_46_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_46_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_46_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_46_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_46_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_46_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_46_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_46_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_46_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_46_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_46_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_46_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_46_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_46_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_46_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[42]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[42]),
    .ccff_tail(grid_clb_46_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__12_
  (
    .clk_0_S_in(clk_1_wires[82]),
    .prog_clk_0_S_in(prog_clk_1_wires[82]),
    .prog_clk_0_N_out(prog_clk_0_wires[175]),
    .prog_clk_0_E_out(prog_clk_0_wires[173]),
    .prog_clk_0_S_out(prog_clk_0_wires[172]),
    .Reset_W_out(ResetWires[272]),
    .Reset_E_in(ResetWires[271]),
    .pReset_N_in(pResetWires[612]),
    .Test_en_W_out(Test_enWires[272]),
    .Test_en_E_in(Test_enWires[271]),
    .SC_OUT_TOP(scff_Wires[104]),
    .SC_IN_BOT(scff_Wires[103]),
    .top_width_0_height_0__pin_0_(cbx_1__12__3_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__3_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__3_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__3_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__3_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__3_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__3_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__3_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__3_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__3_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__3_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__3_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__3_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__3_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__3_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__3_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_4__12__undriven_top_width_0_height_0__pin_32_[0]),
    .top_width_0_height_0__pin_34_(grid_clb_4__12__undriven_top_width_0_height_0__pin_34_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__47_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__47_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__47_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__47_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__47_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__47_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__47_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__47_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__47_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__47_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__47_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__47_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__47_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__47_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__47_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__47_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__35_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_47_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_47_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_47_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_47_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_47_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_47_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_47_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_47_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_47_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_47_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_47_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_47_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_47_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_47_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_47_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_47_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_47_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_47_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_47_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_47_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_47_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_47_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_47_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_47_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_47_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_47_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_47_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_47_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_47_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_47_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_47_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_47_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[43]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[43]),
    .ccff_tail(grid_clb_47_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__1_
  (
    .clk_0_N_in(clk_1_wires[88]),
    .prog_clk_0_N_in(prog_clk_1_wires[88]),
    .prog_clk_0_E_out(prog_clk_0_wires[178]),
    .prog_clk_0_S_out(prog_clk_0_wires[177]),
    .Reset_W_out(ResetWires[32]),
    .Reset_E_in(ResetWires[31]),
    .pReset_N_in(pResetWires[80]),
    .Test_en_W_out(Test_enWires[32]),
    .Test_en_E_in(Test_enWires[31]),
    .SC_OUT_BOT(scff_Wires[131]),
    .SC_IN_TOP(scff_Wires[129]),
    .top_width_0_height_0__pin_0_(cbx_1__1__44_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__44_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__44_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__44_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__44_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__44_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__44_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__44_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__44_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__44_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__44_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__44_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__44_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__44_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__44_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__44_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[44]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[44]),
    .right_width_0_height_0__pin_16_(cby_1__1__48_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__48_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__48_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__48_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__48_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__48_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__48_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__48_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__48_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__48_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__48_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__48_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__48_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__48_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__48_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__48_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__36_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_48_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_48_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_48_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_48_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_48_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_48_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_48_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_48_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_48_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_48_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_48_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_48_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_48_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_48_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_48_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_48_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_48_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_48_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_48_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_48_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_48_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_48_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_48_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_48_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_48_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_48_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_48_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_48_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_48_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_48_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_48_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_48_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(grid_clb_5__1__undriven_bottom_width_0_height_0__pin_52_[0]),
    .bottom_width_0_height_0__pin_54_(grid_clb_5__1__undriven_bottom_width_0_height_0__pin_54_[0]),
    .ccff_tail(grid_clb_48_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__2_
  (
    .clk_0_S_in(clk_1_wires[87]),
    .prog_clk_0_S_in(prog_clk_1_wires[87]),
    .prog_clk_0_E_out(prog_clk_0_wires[181]),
    .prog_clk_0_S_out(prog_clk_0_wires[180]),
    .Reset_W_out(ResetWires[54]),
    .Reset_E_in(ResetWires[53]),
    .pReset_N_in(pResetWires[129]),
    .Test_en_W_out(Test_enWires[54]),
    .Test_en_E_in(Test_enWires[53]),
    .SC_OUT_BOT(scff_Wires[128]),
    .SC_IN_TOP(scff_Wires[127]),
    .top_width_0_height_0__pin_0_(cbx_1__1__45_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__45_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__45_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__45_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__45_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__45_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__45_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__45_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__45_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__45_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__45_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__45_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__45_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__45_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__45_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__45_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[45]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[45]),
    .right_width_0_height_0__pin_16_(cby_1__1__49_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__49_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__49_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__49_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__49_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__49_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__49_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__49_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__49_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__49_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__49_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__49_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__49_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__49_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__49_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__49_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__37_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_49_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_49_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_49_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_49_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_49_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_49_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_49_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_49_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_49_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_49_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_49_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_49_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_49_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_49_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_49_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_49_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_49_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_49_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_49_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_49_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_49_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_49_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_49_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_49_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_49_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_49_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_49_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_49_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_49_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_49_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_49_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_49_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[44]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[44]),
    .ccff_tail(grid_clb_49_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__3_
  (
    .clk_0_N_in(clk_1_wires[95]),
    .prog_clk_0_N_in(prog_clk_1_wires[95]),
    .prog_clk_0_E_out(prog_clk_0_wires[184]),
    .prog_clk_0_S_out(prog_clk_0_wires[183]),
    .Reset_W_out(ResetWires[76]),
    .Reset_E_in(ResetWires[75]),
    .pReset_N_in(pResetWires[178]),
    .Test_en_W_out(Test_enWires[76]),
    .Test_en_E_in(Test_enWires[75]),
    .SC_OUT_BOT(scff_Wires[126]),
    .SC_IN_TOP(scff_Wires[125]),
    .top_width_0_height_0__pin_0_(cbx_1__1__46_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__46_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__46_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__46_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__46_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__46_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__46_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__46_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__46_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__46_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__46_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__46_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__46_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__46_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__46_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__46_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[46]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[46]),
    .right_width_0_height_0__pin_16_(cby_1__1__50_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__50_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__50_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__50_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__50_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__50_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__50_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__50_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__50_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__50_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__50_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__50_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__50_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__50_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__50_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__50_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__38_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_50_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_50_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_50_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_50_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_50_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_50_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_50_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_50_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_50_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_50_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_50_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_50_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_50_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_50_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_50_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_50_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_50_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_50_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_50_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_50_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_50_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_50_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_50_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_50_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_50_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_50_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_50_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_50_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_50_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_50_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_50_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_50_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[45]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[45]),
    .ccff_tail(grid_clb_50_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__4_
  (
    .clk_0_S_in(clk_1_wires[94]),
    .prog_clk_0_S_in(prog_clk_1_wires[94]),
    .prog_clk_0_E_out(prog_clk_0_wires[187]),
    .prog_clk_0_S_out(prog_clk_0_wires[186]),
    .Reset_W_out(ResetWires[98]),
    .Reset_E_in(ResetWires[97]),
    .pReset_N_in(pResetWires[227]),
    .Test_en_W_out(Test_enWires[98]),
    .Test_en_E_in(Test_enWires[97]),
    .SC_OUT_BOT(scff_Wires[124]),
    .SC_IN_TOP(scff_Wires[123]),
    .top_width_0_height_0__pin_0_(cbx_1__1__47_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__47_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__47_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__47_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__47_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__47_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__47_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__47_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__47_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__47_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__47_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__47_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__47_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__47_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__47_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__47_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[47]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[47]),
    .right_width_0_height_0__pin_16_(cby_1__1__51_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__51_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__51_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__51_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__51_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__51_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__51_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__51_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__51_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__51_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__51_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__51_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__51_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__51_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__51_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__51_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__39_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_51_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_51_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_51_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_51_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_51_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_51_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_51_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_51_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_51_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_51_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_51_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_51_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_51_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_51_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_51_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_51_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_51_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_51_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_51_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_51_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_51_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_51_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_51_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_51_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_51_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_51_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_51_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_51_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_51_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_51_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_51_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_51_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[46]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[46]),
    .ccff_tail(grid_clb_51_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__5_
  (
    .clk_0_N_in(clk_1_wires[102]),
    .prog_clk_0_N_in(prog_clk_1_wires[102]),
    .prog_clk_0_E_out(prog_clk_0_wires[190]),
    .prog_clk_0_S_out(prog_clk_0_wires[189]),
    .Reset_W_out(ResetWires[120]),
    .Reset_E_in(ResetWires[119]),
    .pReset_N_in(pResetWires[276]),
    .Test_en_W_out(Test_enWires[120]),
    .Test_en_E_in(Test_enWires[119]),
    .SC_OUT_BOT(scff_Wires[122]),
    .SC_IN_TOP(scff_Wires[121]),
    .top_width_0_height_0__pin_0_(cbx_1__1__48_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__48_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__48_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__48_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__48_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__48_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__48_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__48_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__48_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__48_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__48_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__48_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__48_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__48_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__48_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__48_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[48]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[48]),
    .right_width_0_height_0__pin_16_(cby_1__1__52_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__52_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__52_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__52_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__52_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__52_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__52_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__52_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__52_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__52_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__52_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__52_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__52_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__52_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__52_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__52_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__40_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_52_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_52_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_52_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_52_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_52_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_52_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_52_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_52_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_52_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_52_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_52_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_52_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_52_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_52_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_52_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_52_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_52_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_52_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_52_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_52_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_52_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_52_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_52_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_52_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_52_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_52_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_52_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_52_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_52_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_52_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_52_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_52_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[47]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[47]),
    .ccff_tail(grid_clb_52_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__6_
  (
    .clk_0_S_in(clk_1_wires[101]),
    .prog_clk_0_S_in(prog_clk_1_wires[101]),
    .prog_clk_0_E_out(prog_clk_0_wires[193]),
    .prog_clk_0_S_out(prog_clk_0_wires[192]),
    .Reset_W_out(ResetWires[142]),
    .Reset_E_in(ResetWires[141]),
    .pReset_N_in(pResetWires[325]),
    .Test_en_W_out(Test_enWires[142]),
    .Test_en_E_in(Test_enWires[141]),
    .SC_OUT_BOT(scff_Wires[120]),
    .SC_IN_TOP(scff_Wires[119]),
    .top_width_0_height_0__pin_0_(cbx_1__1__49_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__49_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__49_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__49_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__49_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__49_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__49_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__49_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__49_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__49_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__49_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__49_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__49_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__49_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__49_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__49_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[49]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[49]),
    .right_width_0_height_0__pin_16_(cby_1__1__53_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__53_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__53_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__53_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__53_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__53_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__53_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__53_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__53_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__53_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__53_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__53_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__53_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__53_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__53_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__53_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__41_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_53_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_53_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_53_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_53_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_53_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_53_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_53_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_53_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_53_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_53_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_53_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_53_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_53_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_53_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_53_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_53_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_53_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_53_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_53_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_53_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_53_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_53_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_53_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_53_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_53_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_53_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_53_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_53_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_53_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_53_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_53_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_53_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[48]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[48]),
    .ccff_tail(grid_clb_53_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__7_
  (
    .clk_0_N_in(clk_1_wires[109]),
    .prog_clk_0_N_in(prog_clk_1_wires[109]),
    .prog_clk_0_E_out(prog_clk_0_wires[196]),
    .prog_clk_0_S_out(prog_clk_0_wires[195]),
    .Reset_W_out(ResetWires[164]),
    .Reset_E_in(ResetWires[163]),
    .pReset_N_in(pResetWires[374]),
    .Test_en_W_out(Test_enWires[164]),
    .Test_en_E_in(Test_enWires[163]),
    .SC_OUT_BOT(scff_Wires[118]),
    .SC_IN_TOP(scff_Wires[117]),
    .top_width_0_height_0__pin_0_(cbx_1__1__50_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__50_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__50_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__50_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__50_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__50_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__50_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__50_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__50_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__50_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__50_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__50_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__50_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__50_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__50_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__50_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[50]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[50]),
    .right_width_0_height_0__pin_16_(cby_1__1__54_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__54_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__54_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__54_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__54_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__54_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__54_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__54_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__54_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__54_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__54_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__54_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__54_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__54_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__54_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__54_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__42_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_54_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_54_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_54_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_54_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_54_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_54_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_54_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_54_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_54_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_54_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_54_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_54_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_54_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_54_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_54_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_54_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_54_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_54_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_54_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_54_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_54_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_54_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_54_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_54_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_54_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_54_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_54_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_54_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_54_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_54_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_54_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_54_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[49]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[49]),
    .ccff_tail(grid_clb_54_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__8_
  (
    .clk_0_S_in(clk_1_wires[108]),
    .prog_clk_0_S_in(prog_clk_1_wires[108]),
    .prog_clk_0_E_out(prog_clk_0_wires[199]),
    .prog_clk_0_S_out(prog_clk_0_wires[198]),
    .Reset_W_out(ResetWires[186]),
    .Reset_E_in(ResetWires[185]),
    .pReset_N_in(pResetWires[423]),
    .Test_en_W_out(Test_enWires[186]),
    .Test_en_E_in(Test_enWires[185]),
    .SC_OUT_BOT(scff_Wires[116]),
    .SC_IN_TOP(scff_Wires[115]),
    .top_width_0_height_0__pin_0_(cbx_1__1__51_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__51_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__51_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__51_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__51_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__51_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__51_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__51_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__51_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__51_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__51_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__51_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__51_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__51_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__51_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__51_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[51]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[51]),
    .right_width_0_height_0__pin_16_(cby_1__1__55_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__55_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__55_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__55_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__55_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__55_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__55_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__55_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__55_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__55_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__55_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__55_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__55_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__55_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__55_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__55_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__43_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_55_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_55_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_55_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_55_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_55_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_55_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_55_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_55_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_55_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_55_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_55_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_55_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_55_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_55_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_55_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_55_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_55_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_55_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_55_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_55_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_55_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_55_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_55_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_55_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_55_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_55_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_55_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_55_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_55_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_55_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_55_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_55_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[50]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[50]),
    .ccff_tail(grid_clb_55_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__9_
  (
    .clk_0_N_in(clk_1_wires[116]),
    .prog_clk_0_N_in(prog_clk_1_wires[116]),
    .prog_clk_0_E_out(prog_clk_0_wires[202]),
    .prog_clk_0_S_out(prog_clk_0_wires[201]),
    .Reset_W_out(ResetWires[208]),
    .Reset_E_in(ResetWires[207]),
    .pReset_N_in(pResetWires[472]),
    .Test_en_W_out(Test_enWires[208]),
    .Test_en_E_in(Test_enWires[207]),
    .SC_OUT_BOT(scff_Wires[114]),
    .SC_IN_TOP(scff_Wires[113]),
    .top_width_0_height_0__pin_0_(cbx_1__1__52_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__52_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__52_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__52_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__52_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__52_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__52_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__52_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__52_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__52_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__52_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__52_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__52_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__52_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__52_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__52_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[52]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[52]),
    .right_width_0_height_0__pin_16_(cby_1__1__56_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__56_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__56_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__56_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__56_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__56_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__56_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__56_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__56_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__56_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__56_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__56_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__56_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__56_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__56_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__56_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__44_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_56_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_56_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_56_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_56_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_56_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_56_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_56_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_56_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_56_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_56_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_56_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_56_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_56_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_56_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_56_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_56_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_56_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_56_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_56_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_56_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_56_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_56_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_56_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_56_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_56_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_56_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_56_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_56_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_56_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_56_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_56_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_56_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[51]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[51]),
    .ccff_tail(grid_clb_56_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__10_
  (
    .clk_0_S_in(clk_1_wires[115]),
    .prog_clk_0_S_in(prog_clk_1_wires[115]),
    .prog_clk_0_E_out(prog_clk_0_wires[205]),
    .prog_clk_0_S_out(prog_clk_0_wires[204]),
    .Reset_W_out(ResetWires[230]),
    .Reset_E_in(ResetWires[229]),
    .pReset_N_in(pResetWires[521]),
    .Test_en_W_out(Test_enWires[230]),
    .Test_en_E_in(Test_enWires[229]),
    .SC_OUT_BOT(scff_Wires[112]),
    .SC_IN_TOP(scff_Wires[111]),
    .top_width_0_height_0__pin_0_(cbx_1__1__53_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__53_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__53_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__53_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__53_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__53_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__53_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__53_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__53_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__53_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__53_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__53_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__53_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__53_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__53_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__53_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[53]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[53]),
    .right_width_0_height_0__pin_16_(cby_1__1__57_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__57_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__57_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__57_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__57_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__57_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__57_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__57_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__57_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__57_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__57_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__57_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__57_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__57_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__57_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__57_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__45_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_57_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_57_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_57_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_57_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_57_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_57_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_57_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_57_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_57_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_57_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_57_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_57_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_57_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_57_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_57_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_57_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_57_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_57_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_57_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_57_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_57_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_57_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_57_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_57_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_57_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_57_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_57_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_57_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_57_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_57_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_57_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_57_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[52]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[52]),
    .ccff_tail(grid_clb_57_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__11_
  (
    .clk_0_N_in(clk_1_wires[123]),
    .prog_clk_0_N_in(prog_clk_1_wires[123]),
    .prog_clk_0_E_out(prog_clk_0_wires[208]),
    .prog_clk_0_S_out(prog_clk_0_wires[207]),
    .Reset_W_out(ResetWires[252]),
    .Reset_E_in(ResetWires[251]),
    .pReset_N_in(pResetWires[570]),
    .Test_en_W_out(Test_enWires[252]),
    .Test_en_E_in(Test_enWires[251]),
    .SC_OUT_BOT(scff_Wires[110]),
    .SC_IN_TOP(scff_Wires[109]),
    .top_width_0_height_0__pin_0_(cbx_1__1__54_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__54_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__54_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__54_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__54_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__54_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__54_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__54_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__54_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__54_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__54_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__54_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__54_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__54_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__54_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__54_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[54]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[54]),
    .right_width_0_height_0__pin_16_(cby_1__1__58_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__58_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__58_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__58_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__58_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__58_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__58_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__58_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__58_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__58_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__58_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__58_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__58_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__58_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__58_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__58_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__46_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_58_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_58_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_58_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_58_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_58_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_58_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_58_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_58_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_58_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_58_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_58_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_58_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_58_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_58_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_58_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_58_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_58_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_58_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_58_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_58_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_58_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_58_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_58_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_58_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_58_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_58_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_58_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_58_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_58_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_58_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_58_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_58_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[53]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[53]),
    .ccff_tail(grid_clb_58_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__12_
  (
    .clk_0_S_in(clk_1_wires[122]),
    .prog_clk_0_S_in(prog_clk_1_wires[122]),
    .prog_clk_0_N_out(prog_clk_0_wires[213]),
    .prog_clk_0_E_out(prog_clk_0_wires[211]),
    .prog_clk_0_S_out(prog_clk_0_wires[210]),
    .Reset_W_out(ResetWires[274]),
    .Reset_E_in(ResetWires[273]),
    .pReset_N_in(pResetWires[615]),
    .Test_en_W_out(Test_enWires[274]),
    .Test_en_E_in(Test_enWires[273]),
    .SC_OUT_BOT(scff_Wires[108]),
    .SC_IN_TOP(scff_Wires[107]),
    .top_width_0_height_0__pin_0_(cbx_1__12__4_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__4_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__4_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__4_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__4_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__4_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__4_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__4_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__4_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__4_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__4_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__4_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__4_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__4_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__4_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__4_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_5__12__undriven_top_width_0_height_0__pin_32_[0]),
    .top_width_0_height_0__pin_34_(grid_clb_5__12__undriven_top_width_0_height_0__pin_34_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__59_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__59_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__59_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__59_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__59_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__59_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__59_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__59_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__59_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__59_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__59_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__59_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__59_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__59_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__59_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__59_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__47_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_59_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_59_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_59_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_59_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_59_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_59_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_59_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_59_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_59_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_59_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_59_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_59_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_59_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_59_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_59_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_59_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_59_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_59_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_59_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_59_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_59_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_59_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_59_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_59_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_59_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_59_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_59_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_59_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_59_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_59_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_59_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_59_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[54]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[54]),
    .ccff_tail(grid_clb_59_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__1_
  (
    .clk_0_N_in(clk_1_wires[90]),
    .prog_clk_0_N_in(prog_clk_1_wires[90]),
    .prog_clk_0_E_out(prog_clk_0_wires[216]),
    .prog_clk_0_S_out(prog_clk_0_wires[215]),
    .Reset_W_out(ResetWires[34]),
    .Reset_E_in(ResetWires[33]),
    .pReset_N_in(pResetWires[84]),
    .Test_en_W_out(Test_enWires[34]),
    .Test_en_E_in(Test_enWires[33]),
    .SC_OUT_TOP(scff_Wires[135]),
    .SC_IN_BOT(scff_Wires[134]),
    .top_width_0_height_0__pin_0_(cbx_1__1__55_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__55_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__55_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__55_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__55_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__55_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__55_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__55_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__55_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__55_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__55_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__55_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__55_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__55_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__55_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__55_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[55]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[55]),
    .right_width_0_height_0__pin_16_(cby_1__1__60_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__60_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__60_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__60_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__60_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__60_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__60_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__60_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__60_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__60_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__60_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__60_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__60_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__60_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__60_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__60_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__48_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_60_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_60_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_60_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_60_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_60_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_60_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_60_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_60_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_60_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_60_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_60_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_60_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_60_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_60_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_60_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_60_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_60_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_60_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_60_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_60_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_60_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_60_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_60_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_60_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_60_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_60_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_60_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_60_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_60_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_60_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_60_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_60_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(grid_clb_6__1__undriven_bottom_width_0_height_0__pin_52_[0]),
    .bottom_width_0_height_0__pin_54_(grid_clb_6__1__undriven_bottom_width_0_height_0__pin_54_[0]),
    .ccff_tail(grid_clb_60_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__2_
  (
    .clk_0_S_in(clk_1_wires[89]),
    .prog_clk_0_S_in(prog_clk_1_wires[89]),
    .prog_clk_0_E_out(prog_clk_0_wires[219]),
    .prog_clk_0_S_out(prog_clk_0_wires[218]),
    .Reset_W_out(ResetWires[56]),
    .Reset_E_in(ResetWires[55]),
    .pReset_N_in(pResetWires[133]),
    .Test_en_W_out(Test_enWires[56]),
    .Test_en_E_in(Test_enWires[55]),
    .SC_OUT_TOP(scff_Wires[137]),
    .SC_IN_BOT(scff_Wires[136]),
    .top_width_0_height_0__pin_0_(cbx_1__1__56_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__56_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__56_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__56_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__56_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__56_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__56_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__56_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__56_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__56_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__56_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__56_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__56_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__56_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__56_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__56_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[56]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[56]),
    .right_width_0_height_0__pin_16_(cby_1__1__61_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__61_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__61_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__61_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__61_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__61_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__61_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__61_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__61_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__61_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__61_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__61_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__61_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__61_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__61_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__61_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__49_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_61_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_61_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_61_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_61_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_61_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_61_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_61_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_61_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_61_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_61_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_61_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_61_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_61_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_61_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_61_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_61_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_61_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_61_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_61_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_61_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_61_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_61_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_61_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_61_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_61_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_61_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_61_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_61_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_61_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_61_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_61_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_61_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[55]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[55]),
    .ccff_tail(grid_clb_61_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__3_
  (
    .clk_0_N_in(clk_1_wires[97]),
    .prog_clk_0_N_in(prog_clk_1_wires[97]),
    .prog_clk_0_E_out(prog_clk_0_wires[222]),
    .prog_clk_0_S_out(prog_clk_0_wires[221]),
    .Reset_W_out(ResetWires[78]),
    .Reset_E_in(ResetWires[77]),
    .pReset_N_in(pResetWires[182]),
    .Test_en_W_out(Test_enWires[78]),
    .Test_en_E_in(Test_enWires[77]),
    .SC_OUT_TOP(scff_Wires[139]),
    .SC_IN_BOT(scff_Wires[138]),
    .top_width_0_height_0__pin_0_(cbx_1__1__57_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__57_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__57_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__57_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__57_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__57_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__57_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__57_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__57_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__57_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__57_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__57_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__57_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__57_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__57_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__57_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[57]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[57]),
    .right_width_0_height_0__pin_16_(cby_1__1__62_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__62_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__62_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__62_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__62_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__62_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__62_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__62_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__62_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__62_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__62_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__62_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__62_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__62_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__62_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__62_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__50_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_62_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_62_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_62_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_62_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_62_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_62_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_62_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_62_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_62_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_62_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_62_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_62_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_62_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_62_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_62_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_62_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_62_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_62_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_62_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_62_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_62_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_62_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_62_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_62_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_62_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_62_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_62_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_62_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_62_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_62_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_62_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_62_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[56]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[56]),
    .ccff_tail(grid_clb_62_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__4_
  (
    .clk_0_S_in(clk_1_wires[96]),
    .prog_clk_0_S_in(prog_clk_1_wires[96]),
    .prog_clk_0_E_out(prog_clk_0_wires[225]),
    .prog_clk_0_S_out(prog_clk_0_wires[224]),
    .Reset_W_out(ResetWires[100]),
    .Reset_E_in(ResetWires[99]),
    .pReset_N_in(pResetWires[231]),
    .Test_en_W_out(Test_enWires[100]),
    .Test_en_E_in(Test_enWires[99]),
    .SC_OUT_TOP(scff_Wires[141]),
    .SC_IN_BOT(scff_Wires[140]),
    .top_width_0_height_0__pin_0_(cbx_1__1__58_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__58_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__58_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__58_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__58_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__58_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__58_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__58_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__58_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__58_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__58_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__58_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__58_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__58_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__58_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__58_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[58]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[58]),
    .right_width_0_height_0__pin_16_(cby_1__1__63_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__63_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__63_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__63_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__63_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__63_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__63_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__63_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__63_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__63_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__63_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__63_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__63_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__63_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__63_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__63_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__51_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_63_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_63_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_63_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_63_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_63_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_63_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_63_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_63_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_63_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_63_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_63_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_63_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_63_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_63_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_63_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_63_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_63_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_63_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_63_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_63_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_63_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_63_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_63_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_63_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_63_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_63_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_63_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_63_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_63_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_63_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_63_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_63_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[57]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[57]),
    .ccff_tail(grid_clb_63_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__5_
  (
    .clk_0_N_in(clk_1_wires[104]),
    .prog_clk_0_N_in(prog_clk_1_wires[104]),
    .prog_clk_0_E_out(prog_clk_0_wires[228]),
    .prog_clk_0_S_out(prog_clk_0_wires[227]),
    .Reset_W_out(ResetWires[122]),
    .Reset_E_in(ResetWires[121]),
    .pReset_N_in(pResetWires[280]),
    .Test_en_W_out(Test_enWires[122]),
    .Test_en_E_in(Test_enWires[121]),
    .SC_OUT_TOP(scff_Wires[143]),
    .SC_IN_BOT(scff_Wires[142]),
    .top_width_0_height_0__pin_0_(cbx_1__1__59_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__59_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__59_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__59_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__59_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__59_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__59_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__59_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__59_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__59_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__59_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__59_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__59_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__59_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__59_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__59_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[59]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[59]),
    .right_width_0_height_0__pin_16_(cby_1__1__64_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__64_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__64_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__64_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__64_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__64_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__64_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__64_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__64_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__64_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__64_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__64_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__64_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__64_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__64_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__64_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__52_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_64_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_64_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_64_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_64_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_64_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_64_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_64_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_64_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_64_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_64_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_64_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_64_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_64_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_64_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_64_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_64_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_64_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_64_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_64_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_64_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_64_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_64_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_64_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_64_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_64_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_64_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_64_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_64_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_64_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_64_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_64_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_64_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[58]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[58]),
    .ccff_tail(grid_clb_64_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__6_
  (
    .clk_0_S_in(clk_1_wires[103]),
    .prog_clk_0_S_in(prog_clk_1_wires[103]),
    .prog_clk_0_E_out(prog_clk_0_wires[231]),
    .prog_clk_0_S_out(prog_clk_0_wires[230]),
    .Reset_W_out(ResetWires[144]),
    .Reset_E_in(ResetWires[143]),
    .pReset_N_in(pResetWires[329]),
    .Test_en_W_out(Test_enWires[144]),
    .Test_en_E_in(Test_enWires[143]),
    .SC_OUT_TOP(scff_Wires[145]),
    .SC_IN_BOT(scff_Wires[144]),
    .top_width_0_height_0__pin_0_(cbx_1__1__60_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__60_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__60_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__60_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__60_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__60_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__60_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__60_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__60_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__60_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__60_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__60_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__60_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__60_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__60_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__60_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[60]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[60]),
    .right_width_0_height_0__pin_16_(cby_1__1__65_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__65_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__65_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__65_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__65_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__65_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__65_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__65_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__65_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__65_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__65_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__65_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__65_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__65_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__65_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__65_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__53_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_65_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_65_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_65_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_65_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_65_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_65_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_65_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_65_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_65_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_65_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_65_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_65_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_65_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_65_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_65_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_65_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_65_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_65_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_65_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_65_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_65_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_65_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_65_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_65_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_65_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_65_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_65_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_65_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_65_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_65_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_65_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_65_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[59]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[59]),
    .ccff_tail(grid_clb_65_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__7_
  (
    .clk_0_N_in(clk_1_wires[111]),
    .prog_clk_0_N_in(prog_clk_1_wires[111]),
    .prog_clk_0_E_out(prog_clk_0_wires[234]),
    .prog_clk_0_S_out(prog_clk_0_wires[233]),
    .Reset_W_out(ResetWires[166]),
    .Reset_E_in(ResetWires[165]),
    .pReset_N_in(pResetWires[378]),
    .Test_en_W_out(Test_enWires[166]),
    .Test_en_E_in(Test_enWires[165]),
    .SC_OUT_TOP(scff_Wires[147]),
    .SC_IN_BOT(scff_Wires[146]),
    .top_width_0_height_0__pin_0_(cbx_1__1__61_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__61_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__61_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__61_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__61_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__61_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__61_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__61_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__61_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__61_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__61_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__61_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__61_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__61_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__61_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__61_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[61]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[61]),
    .right_width_0_height_0__pin_16_(cby_1__1__66_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__66_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__66_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__66_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__66_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__66_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__66_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__66_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__66_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__66_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__66_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__66_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__66_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__66_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__66_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__66_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__54_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_66_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_66_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_66_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_66_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_66_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_66_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_66_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_66_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_66_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_66_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_66_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_66_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_66_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_66_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_66_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_66_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_66_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_66_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_66_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_66_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_66_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_66_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_66_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_66_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_66_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_66_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_66_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_66_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_66_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_66_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_66_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_66_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[60]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[60]),
    .ccff_tail(grid_clb_66_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__8_
  (
    .clk_0_S_in(clk_1_wires[110]),
    .prog_clk_0_S_in(prog_clk_1_wires[110]),
    .prog_clk_0_E_out(prog_clk_0_wires[237]),
    .prog_clk_0_S_out(prog_clk_0_wires[236]),
    .Reset_W_out(ResetWires[188]),
    .Reset_E_in(ResetWires[187]),
    .pReset_N_in(pResetWires[427]),
    .Test_en_W_out(Test_enWires[188]),
    .Test_en_E_in(Test_enWires[187]),
    .SC_OUT_TOP(scff_Wires[149]),
    .SC_IN_BOT(scff_Wires[148]),
    .top_width_0_height_0__pin_0_(cbx_1__1__62_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__62_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__62_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__62_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__62_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__62_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__62_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__62_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__62_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__62_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__62_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__62_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__62_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__62_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__62_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__62_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[62]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[62]),
    .right_width_0_height_0__pin_16_(cby_1__1__67_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__67_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__67_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__67_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__67_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__67_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__67_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__67_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__67_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__67_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__67_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__67_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__67_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__67_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__67_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__67_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__55_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_67_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_67_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_67_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_67_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_67_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_67_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_67_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_67_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_67_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_67_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_67_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_67_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_67_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_67_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_67_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_67_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_67_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_67_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_67_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_67_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_67_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_67_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_67_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_67_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_67_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_67_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_67_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_67_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_67_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_67_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_67_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_67_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[61]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[61]),
    .ccff_tail(grid_clb_67_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__9_
  (
    .clk_0_N_in(clk_1_wires[118]),
    .prog_clk_0_N_in(prog_clk_1_wires[118]),
    .prog_clk_0_E_out(prog_clk_0_wires[240]),
    .prog_clk_0_S_out(prog_clk_0_wires[239]),
    .Reset_W_out(ResetWires[210]),
    .Reset_E_in(ResetWires[209]),
    .pReset_N_in(pResetWires[476]),
    .Test_en_W_out(Test_enWires[210]),
    .Test_en_E_in(Test_enWires[209]),
    .SC_OUT_TOP(scff_Wires[151]),
    .SC_IN_BOT(scff_Wires[150]),
    .top_width_0_height_0__pin_0_(cbx_1__1__63_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__63_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__63_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__63_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__63_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__63_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__63_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__63_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__63_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__63_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__63_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__63_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__63_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__63_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__63_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__63_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[63]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[63]),
    .right_width_0_height_0__pin_16_(cby_1__1__68_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__68_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__68_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__68_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__68_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__68_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__68_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__68_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__68_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__68_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__68_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__68_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__68_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__68_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__68_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__68_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__56_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_68_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_68_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_68_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_68_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_68_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_68_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_68_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_68_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_68_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_68_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_68_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_68_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_68_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_68_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_68_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_68_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_68_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_68_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_68_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_68_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_68_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_68_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_68_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_68_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_68_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_68_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_68_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_68_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_68_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_68_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_68_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_68_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[62]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[62]),
    .ccff_tail(grid_clb_68_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__10_
  (
    .clk_0_S_in(clk_1_wires[117]),
    .prog_clk_0_S_in(prog_clk_1_wires[117]),
    .prog_clk_0_E_out(prog_clk_0_wires[243]),
    .prog_clk_0_S_out(prog_clk_0_wires[242]),
    .Reset_W_out(ResetWires[232]),
    .Reset_E_in(ResetWires[231]),
    .pReset_N_in(pResetWires[525]),
    .Test_en_W_out(Test_enWires[232]),
    .Test_en_E_in(Test_enWires[231]),
    .SC_OUT_TOP(scff_Wires[153]),
    .SC_IN_BOT(scff_Wires[152]),
    .top_width_0_height_0__pin_0_(cbx_1__1__64_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__64_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__64_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__64_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__64_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__64_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__64_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__64_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__64_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__64_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__64_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__64_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__64_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__64_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__64_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__64_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[64]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[64]),
    .right_width_0_height_0__pin_16_(cby_1__1__69_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__69_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__69_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__69_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__69_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__69_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__69_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__69_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__69_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__69_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__69_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__69_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__69_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__69_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__69_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__69_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__57_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_69_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_69_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_69_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_69_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_69_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_69_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_69_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_69_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_69_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_69_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_69_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_69_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_69_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_69_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_69_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_69_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_69_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_69_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_69_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_69_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_69_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_69_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_69_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_69_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_69_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_69_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_69_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_69_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_69_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_69_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_69_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_69_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[63]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[63]),
    .ccff_tail(grid_clb_69_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__11_
  (
    .clk_0_N_in(clk_1_wires[125]),
    .prog_clk_0_N_in(prog_clk_1_wires[125]),
    .prog_clk_0_E_out(prog_clk_0_wires[246]),
    .prog_clk_0_S_out(prog_clk_0_wires[245]),
    .Reset_W_out(ResetWires[254]),
    .Reset_E_in(ResetWires[253]),
    .pReset_N_in(pResetWires[574]),
    .Test_en_W_out(Test_enWires[254]),
    .Test_en_E_in(Test_enWires[253]),
    .SC_OUT_TOP(scff_Wires[155]),
    .SC_IN_BOT(scff_Wires[154]),
    .top_width_0_height_0__pin_0_(cbx_1__1__65_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__65_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__65_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__65_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__65_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__65_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__65_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__65_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__65_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__65_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__65_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__65_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__65_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__65_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__65_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__65_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[65]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[65]),
    .right_width_0_height_0__pin_16_(cby_1__1__70_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__70_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__70_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__70_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__70_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__70_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__70_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__70_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__70_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__70_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__70_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__70_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__70_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__70_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__70_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__70_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__58_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_70_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_70_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_70_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_70_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_70_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_70_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_70_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_70_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_70_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_70_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_70_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_70_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_70_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_70_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_70_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_70_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_70_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_70_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_70_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_70_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_70_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_70_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_70_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_70_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_70_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_70_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_70_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_70_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_70_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_70_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_70_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_70_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[64]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[64]),
    .ccff_tail(grid_clb_70_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__12_
  (
    .clk_0_S_in(clk_1_wires[124]),
    .prog_clk_0_S_in(prog_clk_1_wires[124]),
    .prog_clk_0_N_out(prog_clk_0_wires[251]),
    .prog_clk_0_E_out(prog_clk_0_wires[249]),
    .prog_clk_0_S_out(prog_clk_0_wires[248]),
    .Reset_W_out(ResetWires[276]),
    .Reset_E_in(ResetWires[275]),
    .pReset_N_in(pResetWires[618]),
    .Test_en_W_out(Test_enWires[276]),
    .Test_en_E_in(Test_enWires[275]),
    .SC_OUT_TOP(scff_Wires[157]),
    .SC_IN_BOT(scff_Wires[156]),
    .top_width_0_height_0__pin_0_(cbx_1__12__5_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__5_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__5_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__5_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__5_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__5_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__5_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__5_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__5_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__5_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__5_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__5_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__5_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__5_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__5_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__5_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_6__12__undriven_top_width_0_height_0__pin_32_[0]),
    .top_width_0_height_0__pin_34_(grid_clb_6__12__undriven_top_width_0_height_0__pin_34_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__71_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__71_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__71_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__71_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__71_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__71_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__71_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__71_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__71_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__71_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__71_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__71_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__71_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__71_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__71_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__71_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__59_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_71_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_71_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_71_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_71_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_71_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_71_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_71_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_71_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_71_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_71_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_71_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_71_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_71_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_71_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_71_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_71_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_71_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_71_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_71_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_71_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_71_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_71_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_71_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_71_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_71_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_71_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_71_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_71_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_71_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_71_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_71_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_71_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[65]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[65]),
    .ccff_tail(grid_clb_71_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__1_
  (
    .clk_0_N_in(clk_1_wires[130]),
    .prog_clk_0_N_in(prog_clk_1_wires[130]),
    .prog_clk_0_E_out(prog_clk_0_wires[254]),
    .prog_clk_0_S_out(prog_clk_0_wires[253]),
    .Reset_E_out(ResetWires[36]),
    .Reset_W_in(ResetWires[35]),
    .pReset_N_in(pResetWires[88]),
    .Test_en_E_out(Test_enWires[36]),
    .Test_en_W_in(Test_enWires[35]),
    .SC_OUT_BOT(scff_Wires[184]),
    .SC_IN_TOP(scff_Wires[182]),
    .top_width_0_height_0__pin_0_(cbx_1__1__66_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__66_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__66_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__66_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__66_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__66_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__66_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__66_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__66_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__66_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__66_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__66_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__66_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__66_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__66_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__66_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[66]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[66]),
    .right_width_0_height_0__pin_16_(cby_1__1__72_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__72_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__72_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__72_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__72_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__72_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__72_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__72_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__72_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__72_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__72_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__72_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__72_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__72_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__72_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__72_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__60_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_72_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_72_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_72_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_72_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_72_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_72_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_72_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_72_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_72_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_72_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_72_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_72_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_72_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_72_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_72_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_72_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_72_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_72_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_72_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_72_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_72_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_72_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_72_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_72_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_72_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_72_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_72_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_72_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_72_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_72_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_72_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_72_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(grid_clb_7__1__undriven_bottom_width_0_height_0__pin_52_[0]),
    .bottom_width_0_height_0__pin_54_(grid_clb_7__1__undriven_bottom_width_0_height_0__pin_54_[0]),
    .ccff_tail(grid_clb_72_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__2_
  (
    .clk_0_S_in(clk_1_wires[129]),
    .prog_clk_0_S_in(prog_clk_1_wires[129]),
    .prog_clk_0_E_out(prog_clk_0_wires[257]),
    .prog_clk_0_S_out(prog_clk_0_wires[256]),
    .Reset_E_out(ResetWires[58]),
    .Reset_W_in(ResetWires[57]),
    .pReset_N_in(pResetWires[137]),
    .Test_en_E_out(Test_enWires[58]),
    .Test_en_W_in(Test_enWires[57]),
    .SC_OUT_BOT(scff_Wires[181]),
    .SC_IN_TOP(scff_Wires[180]),
    .top_width_0_height_0__pin_0_(cbx_1__1__67_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__67_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__67_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__67_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__67_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__67_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__67_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__67_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__67_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__67_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__67_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__67_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__67_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__67_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__67_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__67_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[67]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[67]),
    .right_width_0_height_0__pin_16_(cby_1__1__73_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__73_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__73_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__73_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__73_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__73_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__73_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__73_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__73_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__73_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__73_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__73_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__73_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__73_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__73_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__73_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__61_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_73_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_73_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_73_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_73_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_73_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_73_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_73_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_73_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_73_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_73_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_73_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_73_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_73_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_73_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_73_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_73_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_73_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_73_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_73_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_73_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_73_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_73_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_73_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_73_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_73_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_73_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_73_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_73_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_73_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_73_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_73_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_73_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[66]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[66]),
    .ccff_tail(grid_clb_73_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__3_
  (
    .clk_0_N_in(clk_1_wires[137]),
    .prog_clk_0_N_in(prog_clk_1_wires[137]),
    .prog_clk_0_E_out(prog_clk_0_wires[260]),
    .prog_clk_0_S_out(prog_clk_0_wires[259]),
    .Reset_E_out(ResetWires[80]),
    .Reset_W_in(ResetWires[79]),
    .pReset_N_in(pResetWires[186]),
    .Test_en_E_out(Test_enWires[80]),
    .Test_en_W_in(Test_enWires[79]),
    .SC_OUT_BOT(scff_Wires[179]),
    .SC_IN_TOP(scff_Wires[178]),
    .top_width_0_height_0__pin_0_(cbx_1__1__68_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__68_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__68_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__68_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__68_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__68_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__68_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__68_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__68_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__68_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__68_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__68_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__68_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__68_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__68_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__68_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[68]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[68]),
    .right_width_0_height_0__pin_16_(cby_1__1__74_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__74_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__74_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__74_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__74_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__74_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__74_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__74_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__74_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__74_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__74_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__74_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__74_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__74_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__74_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__74_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__62_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_74_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_74_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_74_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_74_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_74_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_74_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_74_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_74_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_74_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_74_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_74_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_74_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_74_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_74_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_74_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_74_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_74_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_74_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_74_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_74_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_74_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_74_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_74_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_74_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_74_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_74_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_74_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_74_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_74_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_74_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_74_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_74_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[67]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[67]),
    .ccff_tail(grid_clb_74_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__4_
  (
    .clk_0_S_in(clk_1_wires[136]),
    .prog_clk_0_S_in(prog_clk_1_wires[136]),
    .prog_clk_0_E_out(prog_clk_0_wires[263]),
    .prog_clk_0_S_out(prog_clk_0_wires[262]),
    .Reset_E_out(ResetWires[102]),
    .Reset_W_in(ResetWires[101]),
    .pReset_N_in(pResetWires[235]),
    .Test_en_E_out(Test_enWires[102]),
    .Test_en_W_in(Test_enWires[101]),
    .SC_OUT_BOT(scff_Wires[177]),
    .SC_IN_TOP(scff_Wires[176]),
    .top_width_0_height_0__pin_0_(cbx_1__1__69_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__69_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__69_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__69_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__69_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__69_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__69_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__69_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__69_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__69_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__69_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__69_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__69_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__69_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__69_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__69_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[69]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[69]),
    .right_width_0_height_0__pin_16_(cby_1__1__75_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__75_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__75_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__75_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__75_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__75_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__75_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__75_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__75_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__75_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__75_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__75_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__75_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__75_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__75_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__75_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__63_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_75_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_75_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_75_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_75_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_75_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_75_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_75_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_75_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_75_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_75_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_75_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_75_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_75_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_75_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_75_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_75_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_75_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_75_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_75_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_75_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_75_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_75_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_75_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_75_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_75_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_75_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_75_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_75_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_75_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_75_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_75_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_75_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[68]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[68]),
    .ccff_tail(grid_clb_75_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__5_
  (
    .clk_0_N_in(clk_1_wires[144]),
    .prog_clk_0_N_in(prog_clk_1_wires[144]),
    .prog_clk_0_E_out(prog_clk_0_wires[266]),
    .prog_clk_0_S_out(prog_clk_0_wires[265]),
    .Reset_E_out(ResetWires[124]),
    .Reset_W_in(ResetWires[123]),
    .pReset_N_in(pResetWires[284]),
    .Test_en_E_out(Test_enWires[124]),
    .Test_en_W_in(Test_enWires[123]),
    .SC_OUT_BOT(scff_Wires[175]),
    .SC_IN_TOP(scff_Wires[174]),
    .top_width_0_height_0__pin_0_(cbx_1__1__70_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__70_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__70_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__70_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__70_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__70_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__70_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__70_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__70_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__70_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__70_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__70_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__70_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__70_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__70_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__70_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[70]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[70]),
    .right_width_0_height_0__pin_16_(cby_1__1__76_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__76_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__76_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__76_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__76_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__76_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__76_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__76_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__76_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__76_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__76_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__76_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__76_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__76_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__76_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__76_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__64_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_76_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_76_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_76_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_76_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_76_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_76_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_76_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_76_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_76_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_76_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_76_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_76_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_76_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_76_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_76_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_76_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_76_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_76_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_76_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_76_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_76_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_76_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_76_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_76_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_76_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_76_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_76_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_76_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_76_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_76_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_76_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_76_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[69]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[69]),
    .ccff_tail(grid_clb_76_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__6_
  (
    .clk_0_S_in(clk_1_wires[143]),
    .prog_clk_0_S_in(prog_clk_1_wires[143]),
    .prog_clk_0_E_out(prog_clk_0_wires[269]),
    .prog_clk_0_S_out(prog_clk_0_wires[268]),
    .Reset_E_out(ResetWires[146]),
    .Reset_W_in(ResetWires[145]),
    .pReset_N_in(pResetWires[333]),
    .Test_en_E_out(Test_enWires[146]),
    .Test_en_W_in(Test_enWires[145]),
    .SC_OUT_BOT(scff_Wires[173]),
    .SC_IN_TOP(scff_Wires[172]),
    .top_width_0_height_0__pin_0_(cbx_1__1__71_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__71_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__71_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__71_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__71_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__71_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__71_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__71_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__71_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__71_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__71_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__71_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__71_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__71_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__71_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__71_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[71]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[71]),
    .right_width_0_height_0__pin_16_(cby_1__1__77_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__77_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__77_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__77_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__77_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__77_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__77_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__77_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__77_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__77_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__77_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__77_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__77_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__77_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__77_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__77_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__65_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_77_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_77_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_77_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_77_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_77_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_77_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_77_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_77_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_77_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_77_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_77_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_77_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_77_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_77_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_77_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_77_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_77_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_77_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_77_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_77_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_77_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_77_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_77_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_77_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_77_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_77_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_77_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_77_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_77_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_77_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_77_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_77_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[70]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[70]),
    .ccff_tail(grid_clb_77_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__7_
  (
    .clk_0_N_in(clk_1_wires[151]),
    .prog_clk_0_N_in(prog_clk_1_wires[151]),
    .prog_clk_0_E_out(prog_clk_0_wires[272]),
    .prog_clk_0_S_out(prog_clk_0_wires[271]),
    .Reset_E_out(ResetWires[168]),
    .Reset_W_in(ResetWires[167]),
    .pReset_N_in(pResetWires[382]),
    .Test_en_E_out(Test_enWires[168]),
    .Test_en_W_in(Test_enWires[167]),
    .SC_OUT_BOT(scff_Wires[171]),
    .SC_IN_TOP(scff_Wires[170]),
    .top_width_0_height_0__pin_0_(cbx_1__1__72_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__72_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__72_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__72_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__72_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__72_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__72_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__72_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__72_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__72_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__72_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__72_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__72_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__72_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__72_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__72_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[72]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[72]),
    .right_width_0_height_0__pin_16_(cby_1__1__78_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__78_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__78_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__78_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__78_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__78_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__78_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__78_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__78_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__78_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__78_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__78_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__78_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__78_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__78_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__78_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__66_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_78_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_78_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_78_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_78_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_78_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_78_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_78_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_78_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_78_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_78_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_78_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_78_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_78_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_78_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_78_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_78_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_78_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_78_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_78_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_78_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_78_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_78_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_78_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_78_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_78_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_78_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_78_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_78_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_78_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_78_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_78_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_78_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[71]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[71]),
    .ccff_tail(grid_clb_78_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__8_
  (
    .clk_0_S_in(clk_1_wires[150]),
    .prog_clk_0_S_in(prog_clk_1_wires[150]),
    .prog_clk_0_E_out(prog_clk_0_wires[275]),
    .prog_clk_0_S_out(prog_clk_0_wires[274]),
    .Reset_E_out(ResetWires[190]),
    .Reset_W_in(ResetWires[189]),
    .pReset_N_in(pResetWires[431]),
    .Test_en_E_out(Test_enWires[190]),
    .Test_en_W_in(Test_enWires[189]),
    .SC_OUT_BOT(scff_Wires[169]),
    .SC_IN_TOP(scff_Wires[168]),
    .top_width_0_height_0__pin_0_(cbx_1__1__73_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__73_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__73_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__73_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__73_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__73_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__73_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__73_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__73_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__73_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__73_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__73_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__73_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__73_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__73_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__73_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[73]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[73]),
    .right_width_0_height_0__pin_16_(cby_1__1__79_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__79_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__79_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__79_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__79_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__79_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__79_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__79_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__79_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__79_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__79_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__79_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__79_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__79_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__79_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__79_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__67_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_79_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_79_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_79_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_79_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_79_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_79_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_79_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_79_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_79_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_79_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_79_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_79_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_79_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_79_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_79_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_79_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_79_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_79_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_79_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_79_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_79_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_79_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_79_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_79_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_79_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_79_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_79_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_79_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_79_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_79_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_79_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_79_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[72]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[72]),
    .ccff_tail(grid_clb_79_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__9_
  (
    .clk_0_N_in(clk_1_wires[158]),
    .prog_clk_0_N_in(prog_clk_1_wires[158]),
    .prog_clk_0_E_out(prog_clk_0_wires[278]),
    .prog_clk_0_S_out(prog_clk_0_wires[277]),
    .Reset_E_out(ResetWires[212]),
    .Reset_W_in(ResetWires[211]),
    .pReset_N_in(pResetWires[480]),
    .Test_en_E_out(Test_enWires[212]),
    .Test_en_W_in(Test_enWires[211]),
    .SC_OUT_BOT(scff_Wires[167]),
    .SC_IN_TOP(scff_Wires[166]),
    .top_width_0_height_0__pin_0_(cbx_1__1__74_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__74_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__74_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__74_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__74_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__74_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__74_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__74_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__74_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__74_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__74_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__74_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__74_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__74_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__74_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__74_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[74]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[74]),
    .right_width_0_height_0__pin_16_(cby_1__1__80_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__80_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__80_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__80_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__80_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__80_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__80_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__80_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__80_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__80_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__80_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__80_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__80_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__80_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__80_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__80_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__68_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_80_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_80_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_80_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_80_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_80_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_80_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_80_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_80_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_80_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_80_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_80_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_80_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_80_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_80_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_80_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_80_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_80_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_80_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_80_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_80_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_80_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_80_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_80_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_80_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_80_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_80_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_80_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_80_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_80_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_80_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_80_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_80_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[73]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[73]),
    .ccff_tail(grid_clb_80_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__10_
  (
    .clk_0_S_in(clk_1_wires[157]),
    .prog_clk_0_S_in(prog_clk_1_wires[157]),
    .prog_clk_0_E_out(prog_clk_0_wires[281]),
    .prog_clk_0_S_out(prog_clk_0_wires[280]),
    .Reset_E_out(ResetWires[234]),
    .Reset_W_in(ResetWires[233]),
    .pReset_N_in(pResetWires[529]),
    .Test_en_E_out(Test_enWires[234]),
    .Test_en_W_in(Test_enWires[233]),
    .SC_OUT_BOT(scff_Wires[165]),
    .SC_IN_TOP(scff_Wires[164]),
    .top_width_0_height_0__pin_0_(cbx_1__1__75_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__75_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__75_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__75_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__75_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__75_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__75_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__75_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__75_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__75_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__75_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__75_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__75_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__75_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__75_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__75_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[75]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[75]),
    .right_width_0_height_0__pin_16_(cby_1__1__81_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__81_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__81_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__81_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__81_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__81_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__81_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__81_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__81_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__81_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__81_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__81_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__81_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__81_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__81_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__81_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__69_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_81_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_81_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_81_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_81_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_81_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_81_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_81_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_81_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_81_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_81_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_81_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_81_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_81_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_81_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_81_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_81_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_81_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_81_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_81_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_81_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_81_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_81_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_81_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_81_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_81_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_81_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_81_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_81_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_81_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_81_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_81_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_81_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[74]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[74]),
    .ccff_tail(grid_clb_81_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__11_
  (
    .clk_0_N_in(clk_1_wires[165]),
    .prog_clk_0_N_in(prog_clk_1_wires[165]),
    .prog_clk_0_E_out(prog_clk_0_wires[284]),
    .prog_clk_0_S_out(prog_clk_0_wires[283]),
    .Reset_E_out(ResetWires[256]),
    .Reset_W_in(ResetWires[255]),
    .pReset_N_in(pResetWires[578]),
    .Test_en_E_out(Test_enWires[256]),
    .Test_en_W_in(Test_enWires[255]),
    .SC_OUT_BOT(scff_Wires[163]),
    .SC_IN_TOP(scff_Wires[162]),
    .top_width_0_height_0__pin_0_(cbx_1__1__76_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__76_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__76_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__76_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__76_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__76_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__76_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__76_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__76_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__76_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__76_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__76_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__76_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__76_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__76_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__76_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[76]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[76]),
    .right_width_0_height_0__pin_16_(cby_1__1__82_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__82_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__82_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__82_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__82_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__82_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__82_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__82_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__82_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__82_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__82_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__82_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__82_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__82_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__82_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__82_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__70_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_82_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_82_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_82_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_82_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_82_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_82_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_82_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_82_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_82_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_82_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_82_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_82_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_82_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_82_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_82_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_82_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_82_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_82_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_82_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_82_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_82_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_82_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_82_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_82_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_82_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_82_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_82_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_82_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_82_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_82_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_82_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_82_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[75]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[75]),
    .ccff_tail(grid_clb_82_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__12_
  (
    .clk_0_S_in(clk_1_wires[164]),
    .prog_clk_0_S_in(prog_clk_1_wires[164]),
    .prog_clk_0_N_out(prog_clk_0_wires[289]),
    .prog_clk_0_E_out(prog_clk_0_wires[287]),
    .prog_clk_0_S_out(prog_clk_0_wires[286]),
    .Reset_E_out(ResetWires[278]),
    .Reset_W_in(ResetWires[277]),
    .pReset_N_in(pResetWires[621]),
    .Test_en_E_out(Test_enWires[278]),
    .Test_en_W_in(Test_enWires[277]),
    .SC_OUT_BOT(scff_Wires[161]),
    .SC_IN_TOP(scff_Wires[160]),
    .top_width_0_height_0__pin_0_(cbx_1__12__6_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__6_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__6_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__6_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__6_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__6_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__6_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__6_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__6_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__6_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__6_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__6_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__6_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__6_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__6_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__6_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_7__12__undriven_top_width_0_height_0__pin_32_[0]),
    .top_width_0_height_0__pin_34_(grid_clb_7__12__undriven_top_width_0_height_0__pin_34_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__83_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__83_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__83_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__83_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__83_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__83_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__83_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__83_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__83_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__83_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__83_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__83_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__83_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__83_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__83_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__83_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__71_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_83_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_83_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_83_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_83_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_83_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_83_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_83_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_83_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_83_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_83_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_83_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_83_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_83_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_83_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_83_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_83_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_83_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_83_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_83_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_83_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_83_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_83_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_83_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_83_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_83_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_83_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_83_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_83_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_83_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_83_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_83_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_83_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[76]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[76]),
    .ccff_tail(grid_clb_83_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__1_
  (
    .clk_0_N_in(clk_1_wires[132]),
    .prog_clk_0_N_in(prog_clk_1_wires[132]),
    .prog_clk_0_E_out(prog_clk_0_wires[292]),
    .prog_clk_0_S_out(prog_clk_0_wires[291]),
    .Reset_E_out(ResetWires[38]),
    .Reset_W_in(ResetWires[37]),
    .pReset_N_in(pResetWires[92]),
    .Test_en_E_out(Test_enWires[38]),
    .Test_en_W_in(Test_enWires[37]),
    .SC_OUT_TOP(scff_Wires[188]),
    .SC_IN_BOT(scff_Wires[187]),
    .top_width_0_height_0__pin_0_(cbx_1__1__77_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__77_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__77_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__77_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__77_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__77_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__77_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__77_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__77_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__77_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__77_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__77_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__77_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__77_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__77_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__77_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[77]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[77]),
    .right_width_0_height_0__pin_16_(cby_1__1__84_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__84_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__84_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__84_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__84_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__84_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__84_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__84_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__84_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__84_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__84_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__84_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__84_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__84_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__84_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__84_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__72_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_84_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_84_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_84_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_84_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_84_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_84_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_84_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_84_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_84_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_84_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_84_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_84_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_84_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_84_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_84_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_84_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_84_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_84_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_84_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_84_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_84_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_84_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_84_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_84_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_84_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_84_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_84_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_84_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_84_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_84_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_84_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_84_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(grid_clb_8__1__undriven_bottom_width_0_height_0__pin_52_[0]),
    .bottom_width_0_height_0__pin_54_(grid_clb_8__1__undriven_bottom_width_0_height_0__pin_54_[0]),
    .ccff_tail(grid_clb_84_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__2_
  (
    .clk_0_S_in(clk_1_wires[131]),
    .prog_clk_0_S_in(prog_clk_1_wires[131]),
    .prog_clk_0_E_out(prog_clk_0_wires[295]),
    .prog_clk_0_S_out(prog_clk_0_wires[294]),
    .Reset_E_out(ResetWires[60]),
    .Reset_W_in(ResetWires[59]),
    .pReset_N_in(pResetWires[141]),
    .Test_en_E_out(Test_enWires[60]),
    .Test_en_W_in(Test_enWires[59]),
    .SC_OUT_TOP(scff_Wires[190]),
    .SC_IN_BOT(scff_Wires[189]),
    .top_width_0_height_0__pin_0_(cbx_1__1__78_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__78_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__78_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__78_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__78_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__78_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__78_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__78_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__78_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__78_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__78_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__78_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__78_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__78_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__78_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__78_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[78]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[78]),
    .right_width_0_height_0__pin_16_(cby_1__1__85_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__85_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__85_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__85_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__85_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__85_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__85_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__85_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__85_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__85_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__85_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__85_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__85_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__85_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__85_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__85_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__73_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_85_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_85_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_85_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_85_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_85_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_85_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_85_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_85_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_85_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_85_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_85_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_85_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_85_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_85_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_85_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_85_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_85_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_85_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_85_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_85_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_85_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_85_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_85_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_85_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_85_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_85_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_85_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_85_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_85_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_85_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_85_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_85_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[77]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[77]),
    .ccff_tail(grid_clb_85_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__3_
  (
    .clk_0_N_in(clk_1_wires[139]),
    .prog_clk_0_N_in(prog_clk_1_wires[139]),
    .prog_clk_0_E_out(prog_clk_0_wires[298]),
    .prog_clk_0_S_out(prog_clk_0_wires[297]),
    .Reset_E_out(ResetWires[82]),
    .Reset_W_in(ResetWires[81]),
    .pReset_N_in(pResetWires[190]),
    .Test_en_E_out(Test_enWires[82]),
    .Test_en_W_in(Test_enWires[81]),
    .SC_OUT_TOP(scff_Wires[192]),
    .SC_IN_BOT(scff_Wires[191]),
    .top_width_0_height_0__pin_0_(cbx_1__1__79_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__79_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__79_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__79_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__79_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__79_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__79_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__79_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__79_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__79_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__79_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__79_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__79_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__79_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__79_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__79_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[79]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[79]),
    .right_width_0_height_0__pin_16_(cby_1__1__86_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__86_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__86_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__86_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__86_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__86_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__86_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__86_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__86_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__86_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__86_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__86_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__86_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__86_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__86_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__86_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__74_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_86_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_86_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_86_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_86_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_86_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_86_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_86_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_86_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_86_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_86_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_86_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_86_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_86_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_86_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_86_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_86_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_86_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_86_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_86_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_86_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_86_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_86_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_86_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_86_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_86_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_86_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_86_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_86_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_86_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_86_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_86_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_86_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[78]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[78]),
    .ccff_tail(grid_clb_86_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__4_
  (
    .clk_0_S_in(clk_1_wires[138]),
    .prog_clk_0_S_in(prog_clk_1_wires[138]),
    .prog_clk_0_E_out(prog_clk_0_wires[301]),
    .prog_clk_0_S_out(prog_clk_0_wires[300]),
    .Reset_E_out(ResetWires[104]),
    .Reset_W_in(ResetWires[103]),
    .pReset_N_in(pResetWires[239]),
    .Test_en_E_out(Test_enWires[104]),
    .Test_en_W_in(Test_enWires[103]),
    .SC_OUT_TOP(scff_Wires[194]),
    .SC_IN_BOT(scff_Wires[193]),
    .top_width_0_height_0__pin_0_(cbx_1__1__80_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__80_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__80_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__80_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__80_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__80_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__80_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__80_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__80_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__80_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__80_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__80_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__80_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__80_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__80_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__80_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[80]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[80]),
    .right_width_0_height_0__pin_16_(cby_1__1__87_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__87_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__87_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__87_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__87_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__87_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__87_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__87_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__87_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__87_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__87_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__87_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__87_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__87_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__87_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__87_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__75_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_87_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_87_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_87_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_87_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_87_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_87_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_87_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_87_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_87_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_87_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_87_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_87_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_87_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_87_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_87_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_87_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_87_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_87_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_87_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_87_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_87_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_87_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_87_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_87_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_87_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_87_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_87_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_87_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_87_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_87_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_87_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_87_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[79]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[79]),
    .ccff_tail(grid_clb_87_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__5_
  (
    .clk_0_N_in(clk_1_wires[146]),
    .prog_clk_0_N_in(prog_clk_1_wires[146]),
    .prog_clk_0_E_out(prog_clk_0_wires[304]),
    .prog_clk_0_S_out(prog_clk_0_wires[303]),
    .Reset_E_out(ResetWires[126]),
    .Reset_W_in(ResetWires[125]),
    .pReset_N_in(pResetWires[288]),
    .Test_en_E_out(Test_enWires[126]),
    .Test_en_W_in(Test_enWires[125]),
    .SC_OUT_TOP(scff_Wires[196]),
    .SC_IN_BOT(scff_Wires[195]),
    .top_width_0_height_0__pin_0_(cbx_1__1__81_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__81_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__81_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__81_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__81_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__81_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__81_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__81_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__81_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__81_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__81_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__81_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__81_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__81_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__81_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__81_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[81]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[81]),
    .right_width_0_height_0__pin_16_(cby_1__1__88_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__88_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__88_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__88_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__88_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__88_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__88_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__88_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__88_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__88_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__88_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__88_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__88_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__88_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__88_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__88_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__76_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_88_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_88_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_88_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_88_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_88_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_88_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_88_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_88_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_88_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_88_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_88_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_88_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_88_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_88_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_88_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_88_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_88_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_88_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_88_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_88_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_88_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_88_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_88_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_88_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_88_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_88_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_88_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_88_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_88_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_88_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_88_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_88_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[80]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[80]),
    .ccff_tail(grid_clb_88_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__6_
  (
    .clk_0_S_in(clk_1_wires[145]),
    .prog_clk_0_S_in(prog_clk_1_wires[145]),
    .prog_clk_0_E_out(prog_clk_0_wires[307]),
    .prog_clk_0_S_out(prog_clk_0_wires[306]),
    .Reset_E_out(ResetWires[148]),
    .Reset_W_in(ResetWires[147]),
    .pReset_N_in(pResetWires[337]),
    .Test_en_E_out(Test_enWires[148]),
    .Test_en_W_in(Test_enWires[147]),
    .SC_OUT_TOP(scff_Wires[198]),
    .SC_IN_BOT(scff_Wires[197]),
    .top_width_0_height_0__pin_0_(cbx_1__1__82_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__82_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__82_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__82_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__82_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__82_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__82_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__82_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__82_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__82_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__82_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__82_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__82_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__82_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__82_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__82_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[82]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[82]),
    .right_width_0_height_0__pin_16_(cby_1__1__89_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__89_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__89_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__89_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__89_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__89_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__89_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__89_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__89_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__89_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__89_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__89_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__89_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__89_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__89_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__89_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__77_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_89_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_89_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_89_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_89_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_89_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_89_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_89_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_89_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_89_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_89_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_89_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_89_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_89_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_89_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_89_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_89_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_89_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_89_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_89_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_89_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_89_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_89_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_89_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_89_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_89_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_89_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_89_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_89_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_89_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_89_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_89_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_89_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[81]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[81]),
    .ccff_tail(grid_clb_89_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__7_
  (
    .clk_0_N_in(clk_1_wires[153]),
    .prog_clk_0_N_in(prog_clk_1_wires[153]),
    .prog_clk_0_E_out(prog_clk_0_wires[310]),
    .prog_clk_0_S_out(prog_clk_0_wires[309]),
    .Reset_E_out(ResetWires[170]),
    .Reset_W_in(ResetWires[169]),
    .pReset_N_in(pResetWires[386]),
    .Test_en_E_out(Test_enWires[170]),
    .Test_en_W_in(Test_enWires[169]),
    .SC_OUT_TOP(scff_Wires[200]),
    .SC_IN_BOT(scff_Wires[199]),
    .top_width_0_height_0__pin_0_(cbx_1__1__83_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__83_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__83_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__83_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__83_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__83_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__83_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__83_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__83_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__83_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__83_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__83_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__83_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__83_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__83_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__83_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[83]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[83]),
    .right_width_0_height_0__pin_16_(cby_1__1__90_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__90_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__90_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__90_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__90_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__90_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__90_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__90_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__90_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__90_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__90_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__90_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__90_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__90_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__90_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__90_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__78_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_90_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_90_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_90_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_90_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_90_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_90_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_90_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_90_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_90_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_90_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_90_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_90_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_90_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_90_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_90_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_90_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_90_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_90_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_90_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_90_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_90_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_90_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_90_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_90_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_90_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_90_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_90_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_90_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_90_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_90_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_90_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_90_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[82]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[82]),
    .ccff_tail(grid_clb_90_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__8_
  (
    .clk_0_S_in(clk_1_wires[152]),
    .prog_clk_0_S_in(prog_clk_1_wires[152]),
    .prog_clk_0_E_out(prog_clk_0_wires[313]),
    .prog_clk_0_S_out(prog_clk_0_wires[312]),
    .Reset_E_out(ResetWires[192]),
    .Reset_W_in(ResetWires[191]),
    .pReset_N_in(pResetWires[435]),
    .Test_en_E_out(Test_enWires[192]),
    .Test_en_W_in(Test_enWires[191]),
    .SC_OUT_TOP(scff_Wires[202]),
    .SC_IN_BOT(scff_Wires[201]),
    .top_width_0_height_0__pin_0_(cbx_1__1__84_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__84_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__84_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__84_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__84_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__84_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__84_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__84_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__84_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__84_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__84_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__84_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__84_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__84_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__84_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__84_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[84]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[84]),
    .right_width_0_height_0__pin_16_(cby_1__1__91_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__91_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__91_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__91_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__91_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__91_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__91_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__91_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__91_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__91_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__91_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__91_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__91_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__91_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__91_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__91_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__79_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_91_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_91_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_91_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_91_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_91_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_91_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_91_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_91_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_91_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_91_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_91_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_91_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_91_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_91_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_91_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_91_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_91_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_91_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_91_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_91_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_91_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_91_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_91_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_91_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_91_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_91_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_91_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_91_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_91_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_91_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_91_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_91_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[83]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[83]),
    .ccff_tail(grid_clb_91_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__9_
  (
    .clk_0_N_in(clk_1_wires[160]),
    .prog_clk_0_N_in(prog_clk_1_wires[160]),
    .prog_clk_0_E_out(prog_clk_0_wires[316]),
    .prog_clk_0_S_out(prog_clk_0_wires[315]),
    .Reset_E_out(ResetWires[214]),
    .Reset_W_in(ResetWires[213]),
    .pReset_N_in(pResetWires[484]),
    .Test_en_E_out(Test_enWires[214]),
    .Test_en_W_in(Test_enWires[213]),
    .SC_OUT_TOP(scff_Wires[204]),
    .SC_IN_BOT(scff_Wires[203]),
    .top_width_0_height_0__pin_0_(cbx_1__1__85_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__85_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__85_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__85_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__85_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__85_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__85_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__85_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__85_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__85_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__85_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__85_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__85_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__85_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__85_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__85_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[85]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[85]),
    .right_width_0_height_0__pin_16_(cby_1__1__92_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__92_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__92_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__92_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__92_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__92_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__92_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__92_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__92_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__92_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__92_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__92_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__92_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__92_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__92_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__92_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__80_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_92_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_92_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_92_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_92_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_92_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_92_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_92_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_92_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_92_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_92_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_92_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_92_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_92_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_92_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_92_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_92_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_92_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_92_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_92_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_92_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_92_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_92_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_92_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_92_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_92_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_92_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_92_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_92_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_92_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_92_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_92_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_92_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[84]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[84]),
    .ccff_tail(grid_clb_92_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__10_
  (
    .clk_0_S_in(clk_1_wires[159]),
    .prog_clk_0_S_in(prog_clk_1_wires[159]),
    .prog_clk_0_E_out(prog_clk_0_wires[319]),
    .prog_clk_0_S_out(prog_clk_0_wires[318]),
    .Reset_E_out(ResetWires[236]),
    .Reset_W_in(ResetWires[235]),
    .pReset_N_in(pResetWires[533]),
    .Test_en_E_out(Test_enWires[236]),
    .Test_en_W_in(Test_enWires[235]),
    .SC_OUT_TOP(scff_Wires[206]),
    .SC_IN_BOT(scff_Wires[205]),
    .top_width_0_height_0__pin_0_(cbx_1__1__86_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__86_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__86_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__86_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__86_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__86_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__86_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__86_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__86_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__86_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__86_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__86_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__86_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__86_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__86_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__86_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[86]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[86]),
    .right_width_0_height_0__pin_16_(cby_1__1__93_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__93_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__93_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__93_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__93_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__93_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__93_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__93_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__93_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__93_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__93_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__93_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__93_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__93_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__93_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__93_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__81_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_93_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_93_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_93_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_93_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_93_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_93_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_93_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_93_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_93_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_93_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_93_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_93_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_93_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_93_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_93_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_93_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_93_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_93_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_93_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_93_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_93_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_93_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_93_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_93_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_93_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_93_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_93_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_93_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_93_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_93_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_93_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_93_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[85]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[85]),
    .ccff_tail(grid_clb_93_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__11_
  (
    .clk_0_N_in(clk_1_wires[167]),
    .prog_clk_0_N_in(prog_clk_1_wires[167]),
    .prog_clk_0_E_out(prog_clk_0_wires[322]),
    .prog_clk_0_S_out(prog_clk_0_wires[321]),
    .Reset_E_out(ResetWires[258]),
    .Reset_W_in(ResetWires[257]),
    .pReset_N_in(pResetWires[582]),
    .Test_en_E_out(Test_enWires[258]),
    .Test_en_W_in(Test_enWires[257]),
    .SC_OUT_TOP(scff_Wires[208]),
    .SC_IN_BOT(scff_Wires[207]),
    .top_width_0_height_0__pin_0_(cbx_1__1__87_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__87_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__87_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__87_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__87_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__87_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__87_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__87_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__87_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__87_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__87_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__87_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__87_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__87_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__87_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__87_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[87]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[87]),
    .right_width_0_height_0__pin_16_(cby_1__1__94_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__94_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__94_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__94_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__94_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__94_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__94_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__94_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__94_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__94_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__94_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__94_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__94_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__94_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__94_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__94_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__82_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_94_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_94_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_94_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_94_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_94_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_94_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_94_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_94_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_94_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_94_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_94_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_94_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_94_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_94_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_94_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_94_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_94_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_94_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_94_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_94_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_94_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_94_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_94_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_94_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_94_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_94_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_94_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_94_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_94_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_94_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_94_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_94_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[86]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[86]),
    .ccff_tail(grid_clb_94_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__12_
  (
    .clk_0_S_in(clk_1_wires[166]),
    .prog_clk_0_S_in(prog_clk_1_wires[166]),
    .prog_clk_0_N_out(prog_clk_0_wires[327]),
    .prog_clk_0_E_out(prog_clk_0_wires[325]),
    .prog_clk_0_S_out(prog_clk_0_wires[324]),
    .Reset_E_out(ResetWires[280]),
    .Reset_W_in(ResetWires[279]),
    .pReset_N_in(pResetWires[624]),
    .Test_en_E_out(Test_enWires[280]),
    .Test_en_W_in(Test_enWires[279]),
    .SC_OUT_TOP(scff_Wires[210]),
    .SC_IN_BOT(scff_Wires[209]),
    .top_width_0_height_0__pin_0_(cbx_1__12__7_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__7_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__7_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__7_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__7_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__7_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__7_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__7_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__7_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__7_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__7_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__7_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__7_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__7_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__7_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__7_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_8__12__undriven_top_width_0_height_0__pin_32_[0]),
    .top_width_0_height_0__pin_34_(grid_clb_8__12__undriven_top_width_0_height_0__pin_34_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__95_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__95_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__95_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__95_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__95_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__95_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__95_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__95_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__95_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__95_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__95_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__95_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__95_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__95_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__95_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__95_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__83_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_95_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_95_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_95_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_95_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_95_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_95_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_95_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_95_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_95_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_95_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_95_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_95_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_95_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_95_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_95_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_95_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_95_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_95_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_95_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_95_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_95_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_95_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_95_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_95_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_95_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_95_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_95_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_95_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_95_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_95_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_95_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_95_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[87]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[87]),
    .ccff_tail(grid_clb_95_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__1_
  (
    .clk_0_N_in(clk_1_wires[172]),
    .prog_clk_0_N_in(prog_clk_1_wires[172]),
    .prog_clk_0_E_out(prog_clk_0_wires[330]),
    .prog_clk_0_S_out(prog_clk_0_wires[329]),
    .Reset_E_out(ResetWires[40]),
    .Reset_W_in(ResetWires[39]),
    .pReset_N_in(pResetWires[96]),
    .Test_en_E_out(Test_enWires[40]),
    .Test_en_W_in(Test_enWires[39]),
    .SC_OUT_BOT(scff_Wires[237]),
    .SC_IN_TOP(scff_Wires[235]),
    .top_width_0_height_0__pin_0_(cbx_1__1__88_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__88_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__88_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__88_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__88_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__88_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__88_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__88_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__88_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__88_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__88_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__88_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__88_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__88_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__88_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__88_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[88]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[88]),
    .right_width_0_height_0__pin_16_(cby_1__1__96_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__96_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__96_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__96_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__96_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__96_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__96_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__96_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__96_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__96_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__96_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__96_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__96_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__96_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__96_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__96_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__84_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_96_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_96_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_96_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_96_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_96_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_96_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_96_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_96_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_96_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_96_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_96_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_96_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_96_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_96_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_96_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_96_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_96_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_96_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_96_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_96_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_96_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_96_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_96_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_96_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_96_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_96_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_96_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_96_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_96_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_96_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_96_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_96_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(grid_clb_9__1__undriven_bottom_width_0_height_0__pin_52_[0]),
    .bottom_width_0_height_0__pin_54_(grid_clb_9__1__undriven_bottom_width_0_height_0__pin_54_[0]),
    .ccff_tail(grid_clb_96_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__2_
  (
    .clk_0_S_in(clk_1_wires[171]),
    .prog_clk_0_S_in(prog_clk_1_wires[171]),
    .prog_clk_0_E_out(prog_clk_0_wires[333]),
    .prog_clk_0_S_out(prog_clk_0_wires[332]),
    .Reset_E_out(ResetWires[62]),
    .Reset_W_in(ResetWires[61]),
    .pReset_N_in(pResetWires[145]),
    .Test_en_E_out(Test_enWires[62]),
    .Test_en_W_in(Test_enWires[61]),
    .SC_OUT_BOT(scff_Wires[234]),
    .SC_IN_TOP(scff_Wires[233]),
    .top_width_0_height_0__pin_0_(cbx_1__1__89_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__89_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__89_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__89_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__89_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__89_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__89_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__89_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__89_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__89_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__89_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__89_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__89_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__89_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__89_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__89_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[89]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[89]),
    .right_width_0_height_0__pin_16_(cby_1__1__97_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__97_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__97_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__97_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__97_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__97_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__97_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__97_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__97_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__97_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__97_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__97_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__97_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__97_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__97_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__97_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__85_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_97_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_97_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_97_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_97_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_97_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_97_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_97_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_97_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_97_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_97_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_97_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_97_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_97_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_97_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_97_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_97_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_97_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_97_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_97_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_97_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_97_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_97_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_97_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_97_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_97_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_97_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_97_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_97_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_97_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_97_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_97_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_97_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[88]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[88]),
    .ccff_tail(grid_clb_97_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__3_
  (
    .clk_0_N_in(clk_1_wires[179]),
    .prog_clk_0_N_in(prog_clk_1_wires[179]),
    .prog_clk_0_E_out(prog_clk_0_wires[336]),
    .prog_clk_0_S_out(prog_clk_0_wires[335]),
    .Reset_E_out(ResetWires[84]),
    .Reset_W_in(ResetWires[83]),
    .pReset_N_in(pResetWires[194]),
    .Test_en_E_out(Test_enWires[84]),
    .Test_en_W_in(Test_enWires[83]),
    .SC_OUT_BOT(scff_Wires[232]),
    .SC_IN_TOP(scff_Wires[231]),
    .top_width_0_height_0__pin_0_(cbx_1__1__90_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__90_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__90_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__90_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__90_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__90_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__90_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__90_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__90_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__90_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__90_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__90_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__90_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__90_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__90_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__90_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[90]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[90]),
    .right_width_0_height_0__pin_16_(cby_1__1__98_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__98_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__98_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__98_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__98_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__98_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__98_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__98_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__98_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__98_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__98_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__98_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__98_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__98_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__98_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__98_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__86_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_98_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_98_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_98_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_98_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_98_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_98_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_98_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_98_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_98_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_98_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_98_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_98_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_98_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_98_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_98_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_98_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_98_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_98_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_98_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_98_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_98_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_98_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_98_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_98_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_98_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_98_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_98_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_98_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_98_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_98_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_98_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_98_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[89]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[89]),
    .ccff_tail(grid_clb_98_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__4_
  (
    .clk_0_S_in(clk_1_wires[178]),
    .prog_clk_0_S_in(prog_clk_1_wires[178]),
    .prog_clk_0_E_out(prog_clk_0_wires[339]),
    .prog_clk_0_S_out(prog_clk_0_wires[338]),
    .Reset_E_out(ResetWires[106]),
    .Reset_W_in(ResetWires[105]),
    .pReset_N_in(pResetWires[243]),
    .Test_en_E_out(Test_enWires[106]),
    .Test_en_W_in(Test_enWires[105]),
    .SC_OUT_BOT(scff_Wires[230]),
    .SC_IN_TOP(scff_Wires[229]),
    .top_width_0_height_0__pin_0_(cbx_1__1__91_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__91_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__91_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__91_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__91_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__91_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__91_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__91_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__91_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__91_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__91_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__91_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__91_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__91_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__91_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__91_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[91]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[91]),
    .right_width_0_height_0__pin_16_(cby_1__1__99_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__99_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__99_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__99_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__99_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__99_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__99_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__99_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__99_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__99_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__99_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__99_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__99_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__99_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__99_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__99_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__87_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_99_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_99_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_99_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_99_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_99_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_99_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_99_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_99_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_99_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_99_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_99_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_99_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_99_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_99_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_99_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_99_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_99_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_99_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_99_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_99_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_99_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_99_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_99_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_99_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_99_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_99_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_99_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_99_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_99_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_99_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_99_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_99_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[90]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[90]),
    .ccff_tail(grid_clb_99_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__5_
  (
    .clk_0_N_in(clk_1_wires[186]),
    .prog_clk_0_N_in(prog_clk_1_wires[186]),
    .prog_clk_0_E_out(prog_clk_0_wires[342]),
    .prog_clk_0_S_out(prog_clk_0_wires[341]),
    .Reset_E_out(ResetWires[128]),
    .Reset_W_in(ResetWires[127]),
    .pReset_N_in(pResetWires[292]),
    .Test_en_E_out(Test_enWires[128]),
    .Test_en_W_in(Test_enWires[127]),
    .SC_OUT_BOT(scff_Wires[228]),
    .SC_IN_TOP(scff_Wires[227]),
    .top_width_0_height_0__pin_0_(cbx_1__1__92_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__92_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__92_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__92_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__92_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__92_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__92_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__92_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__92_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__92_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__92_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__92_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__92_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__92_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__92_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__92_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[92]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[92]),
    .right_width_0_height_0__pin_16_(cby_1__1__100_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__100_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__100_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__100_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__100_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__100_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__100_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__100_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__100_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__100_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__100_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__100_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__100_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__100_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__100_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__100_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__88_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_100_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_100_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_100_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_100_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_100_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_100_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_100_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_100_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_100_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_100_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_100_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_100_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_100_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_100_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_100_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_100_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_100_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_100_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_100_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_100_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_100_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_100_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_100_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_100_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_100_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_100_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_100_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_100_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_100_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_100_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_100_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_100_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[91]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[91]),
    .ccff_tail(grid_clb_100_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__6_
  (
    .clk_0_S_in(clk_1_wires[185]),
    .prog_clk_0_S_in(prog_clk_1_wires[185]),
    .prog_clk_0_E_out(prog_clk_0_wires[345]),
    .prog_clk_0_S_out(prog_clk_0_wires[344]),
    .Reset_E_out(ResetWires[150]),
    .Reset_W_in(ResetWires[149]),
    .pReset_N_in(pResetWires[341]),
    .Test_en_E_out(Test_enWires[150]),
    .Test_en_W_in(Test_enWires[149]),
    .SC_OUT_BOT(scff_Wires[226]),
    .SC_IN_TOP(scff_Wires[225]),
    .top_width_0_height_0__pin_0_(cbx_1__1__93_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__93_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__93_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__93_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__93_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__93_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__93_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__93_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__93_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__93_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__93_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__93_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__93_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__93_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__93_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__93_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[93]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[93]),
    .right_width_0_height_0__pin_16_(cby_1__1__101_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__101_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__101_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__101_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__101_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__101_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__101_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__101_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__101_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__101_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__101_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__101_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__101_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__101_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__101_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__101_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__89_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_101_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_101_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_101_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_101_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_101_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_101_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_101_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_101_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_101_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_101_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_101_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_101_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_101_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_101_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_101_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_101_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_101_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_101_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_101_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_101_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_101_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_101_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_101_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_101_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_101_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_101_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_101_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_101_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_101_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_101_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_101_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_101_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[92]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[92]),
    .ccff_tail(grid_clb_101_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__7_
  (
    .clk_0_N_in(clk_1_wires[193]),
    .prog_clk_0_N_in(prog_clk_1_wires[193]),
    .prog_clk_0_E_out(prog_clk_0_wires[348]),
    .prog_clk_0_S_out(prog_clk_0_wires[347]),
    .Reset_E_out(ResetWires[172]),
    .Reset_W_in(ResetWires[171]),
    .pReset_N_in(pResetWires[390]),
    .Test_en_E_out(Test_enWires[172]),
    .Test_en_W_in(Test_enWires[171]),
    .SC_OUT_BOT(scff_Wires[224]),
    .SC_IN_TOP(scff_Wires[223]),
    .top_width_0_height_0__pin_0_(cbx_1__1__94_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__94_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__94_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__94_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__94_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__94_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__94_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__94_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__94_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__94_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__94_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__94_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__94_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__94_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__94_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__94_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[94]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[94]),
    .right_width_0_height_0__pin_16_(cby_1__1__102_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__102_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__102_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__102_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__102_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__102_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__102_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__102_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__102_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__102_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__102_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__102_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__102_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__102_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__102_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__102_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__90_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_102_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_102_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_102_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_102_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_102_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_102_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_102_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_102_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_102_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_102_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_102_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_102_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_102_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_102_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_102_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_102_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_102_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_102_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_102_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_102_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_102_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_102_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_102_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_102_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_102_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_102_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_102_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_102_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_102_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_102_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_102_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_102_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[93]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[93]),
    .ccff_tail(grid_clb_102_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__8_
  (
    .clk_0_S_in(clk_1_wires[192]),
    .prog_clk_0_S_in(prog_clk_1_wires[192]),
    .prog_clk_0_E_out(prog_clk_0_wires[351]),
    .prog_clk_0_S_out(prog_clk_0_wires[350]),
    .Reset_E_out(ResetWires[194]),
    .Reset_W_in(ResetWires[193]),
    .pReset_N_in(pResetWires[439]),
    .Test_en_E_out(Test_enWires[194]),
    .Test_en_W_in(Test_enWires[193]),
    .SC_OUT_BOT(scff_Wires[222]),
    .SC_IN_TOP(scff_Wires[221]),
    .top_width_0_height_0__pin_0_(cbx_1__1__95_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__95_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__95_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__95_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__95_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__95_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__95_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__95_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__95_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__95_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__95_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__95_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__95_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__95_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__95_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__95_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[95]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[95]),
    .right_width_0_height_0__pin_16_(cby_1__1__103_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__103_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__103_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__103_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__103_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__103_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__103_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__103_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__103_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__103_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__103_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__103_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__103_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__103_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__103_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__103_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__91_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_103_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_103_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_103_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_103_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_103_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_103_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_103_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_103_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_103_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_103_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_103_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_103_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_103_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_103_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_103_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_103_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_103_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_103_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_103_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_103_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_103_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_103_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_103_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_103_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_103_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_103_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_103_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_103_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_103_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_103_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_103_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_103_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[94]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[94]),
    .ccff_tail(grid_clb_103_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__9_
  (
    .clk_0_N_in(clk_1_wires[200]),
    .prog_clk_0_N_in(prog_clk_1_wires[200]),
    .prog_clk_0_E_out(prog_clk_0_wires[354]),
    .prog_clk_0_S_out(prog_clk_0_wires[353]),
    .Reset_E_out(ResetWires[216]),
    .Reset_W_in(ResetWires[215]),
    .pReset_N_in(pResetWires[488]),
    .Test_en_E_out(Test_enWires[216]),
    .Test_en_W_in(Test_enWires[215]),
    .SC_OUT_BOT(scff_Wires[220]),
    .SC_IN_TOP(scff_Wires[219]),
    .top_width_0_height_0__pin_0_(cbx_1__1__96_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__96_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__96_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__96_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__96_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__96_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__96_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__96_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__96_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__96_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__96_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__96_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__96_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__96_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__96_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__96_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[96]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[96]),
    .right_width_0_height_0__pin_16_(cby_1__1__104_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__104_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__104_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__104_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__104_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__104_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__104_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__104_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__104_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__104_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__104_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__104_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__104_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__104_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__104_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__104_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__92_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_104_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_104_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_104_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_104_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_104_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_104_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_104_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_104_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_104_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_104_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_104_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_104_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_104_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_104_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_104_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_104_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_104_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_104_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_104_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_104_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_104_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_104_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_104_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_104_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_104_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_104_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_104_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_104_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_104_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_104_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_104_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_104_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[95]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[95]),
    .ccff_tail(grid_clb_104_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__10_
  (
    .clk_0_S_in(clk_1_wires[199]),
    .prog_clk_0_S_in(prog_clk_1_wires[199]),
    .prog_clk_0_E_out(prog_clk_0_wires[357]),
    .prog_clk_0_S_out(prog_clk_0_wires[356]),
    .Reset_E_out(ResetWires[238]),
    .Reset_W_in(ResetWires[237]),
    .pReset_N_in(pResetWires[537]),
    .Test_en_E_out(Test_enWires[238]),
    .Test_en_W_in(Test_enWires[237]),
    .SC_OUT_BOT(scff_Wires[218]),
    .SC_IN_TOP(scff_Wires[217]),
    .top_width_0_height_0__pin_0_(cbx_1__1__97_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__97_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__97_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__97_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__97_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__97_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__97_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__97_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__97_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__97_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__97_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__97_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__97_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__97_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__97_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__97_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[97]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[97]),
    .right_width_0_height_0__pin_16_(cby_1__1__105_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__105_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__105_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__105_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__105_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__105_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__105_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__105_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__105_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__105_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__105_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__105_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__105_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__105_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__105_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__105_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__93_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_105_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_105_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_105_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_105_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_105_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_105_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_105_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_105_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_105_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_105_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_105_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_105_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_105_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_105_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_105_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_105_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_105_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_105_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_105_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_105_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_105_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_105_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_105_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_105_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_105_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_105_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_105_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_105_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_105_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_105_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_105_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_105_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[96]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[96]),
    .ccff_tail(grid_clb_105_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__11_
  (
    .clk_0_N_in(clk_1_wires[207]),
    .prog_clk_0_N_in(prog_clk_1_wires[207]),
    .prog_clk_0_E_out(prog_clk_0_wires[360]),
    .prog_clk_0_S_out(prog_clk_0_wires[359]),
    .Reset_E_out(ResetWires[260]),
    .Reset_W_in(ResetWires[259]),
    .pReset_N_in(pResetWires[586]),
    .Test_en_E_out(Test_enWires[260]),
    .Test_en_W_in(Test_enWires[259]),
    .SC_OUT_BOT(scff_Wires[216]),
    .SC_IN_TOP(scff_Wires[215]),
    .top_width_0_height_0__pin_0_(cbx_1__1__98_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__98_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__98_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__98_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__98_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__98_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__98_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__98_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__98_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__98_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__98_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__98_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__98_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__98_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__98_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__98_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[98]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[98]),
    .right_width_0_height_0__pin_16_(cby_1__1__106_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__106_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__106_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__106_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__106_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__106_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__106_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__106_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__106_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__106_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__106_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__106_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__106_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__106_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__106_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__106_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__94_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_106_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_106_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_106_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_106_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_106_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_106_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_106_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_106_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_106_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_106_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_106_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_106_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_106_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_106_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_106_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_106_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_106_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_106_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_106_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_106_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_106_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_106_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_106_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_106_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_106_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_106_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_106_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_106_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_106_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_106_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_106_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_106_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[97]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[97]),
    .ccff_tail(grid_clb_106_ccff_tail[0])
  );


  grid_clb
  grid_clb_9__12_
  (
    .clk_0_S_in(clk_1_wires[206]),
    .prog_clk_0_S_in(prog_clk_1_wires[206]),
    .prog_clk_0_N_out(prog_clk_0_wires[365]),
    .prog_clk_0_E_out(prog_clk_0_wires[363]),
    .prog_clk_0_S_out(prog_clk_0_wires[362]),
    .Reset_E_out(ResetWires[282]),
    .Reset_W_in(ResetWires[281]),
    .pReset_N_in(pResetWires[627]),
    .Test_en_E_out(Test_enWires[282]),
    .Test_en_W_in(Test_enWires[281]),
    .SC_OUT_BOT(scff_Wires[214]),
    .SC_IN_TOP(scff_Wires[213]),
    .top_width_0_height_0__pin_0_(cbx_1__12__8_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__8_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__8_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__8_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__8_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__8_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__8_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__8_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__8_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__8_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__8_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__8_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__8_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__8_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__8_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__8_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_9__12__undriven_top_width_0_height_0__pin_32_[0]),
    .top_width_0_height_0__pin_34_(grid_clb_9__12__undriven_top_width_0_height_0__pin_34_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__107_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__107_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__107_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__107_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__107_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__107_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__107_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__107_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__107_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__107_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__107_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__107_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__107_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__107_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__107_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__107_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__95_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_107_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_107_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_107_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_107_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_107_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_107_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_107_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_107_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_107_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_107_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_107_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_107_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_107_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_107_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_107_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_107_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_107_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_107_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_107_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_107_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_107_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_107_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_107_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_107_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_107_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_107_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_107_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_107_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_107_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_107_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_107_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_107_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[98]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[98]),
    .ccff_tail(grid_clb_107_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__1_
  (
    .clk_0_N_in(clk_1_wires[174]),
    .prog_clk_0_N_in(prog_clk_1_wires[174]),
    .prog_clk_0_E_out(prog_clk_0_wires[368]),
    .prog_clk_0_S_out(prog_clk_0_wires[367]),
    .Reset_E_out(ResetWires[42]),
    .Reset_W_in(ResetWires[41]),
    .pReset_N_in(pResetWires[100]),
    .Test_en_E_out(Test_enWires[42]),
    .Test_en_W_in(Test_enWires[41]),
    .SC_OUT_TOP(scff_Wires[241]),
    .SC_IN_BOT(scff_Wires[240]),
    .top_width_0_height_0__pin_0_(cbx_1__1__99_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__99_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__99_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__99_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__99_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__99_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__99_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__99_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__99_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__99_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__99_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__99_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__99_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__99_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__99_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__99_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[99]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[99]),
    .right_width_0_height_0__pin_16_(cby_1__1__108_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__108_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__108_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__108_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__108_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__108_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__108_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__108_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__108_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__108_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__108_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__108_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__108_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__108_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__108_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__108_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__96_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_108_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_108_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_108_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_108_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_108_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_108_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_108_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_108_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_108_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_108_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_108_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_108_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_108_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_108_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_108_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_108_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_108_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_108_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_108_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_108_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_108_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_108_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_108_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_108_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_108_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_108_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_108_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_108_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_108_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_108_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_108_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_108_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(grid_clb_10__1__undriven_bottom_width_0_height_0__pin_52_[0]),
    .bottom_width_0_height_0__pin_54_(grid_clb_10__1__undriven_bottom_width_0_height_0__pin_54_[0]),
    .ccff_tail(grid_clb_108_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__2_
  (
    .clk_0_S_in(clk_1_wires[173]),
    .prog_clk_0_S_in(prog_clk_1_wires[173]),
    .prog_clk_0_E_out(prog_clk_0_wires[371]),
    .prog_clk_0_S_out(prog_clk_0_wires[370]),
    .Reset_E_out(ResetWires[64]),
    .Reset_W_in(ResetWires[63]),
    .pReset_N_in(pResetWires[149]),
    .Test_en_E_out(Test_enWires[64]),
    .Test_en_W_in(Test_enWires[63]),
    .SC_OUT_TOP(scff_Wires[243]),
    .SC_IN_BOT(scff_Wires[242]),
    .top_width_0_height_0__pin_0_(cbx_1__1__100_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__100_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__100_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__100_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__100_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__100_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__100_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__100_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__100_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__100_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__100_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__100_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__100_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__100_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__100_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__100_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[100]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[100]),
    .right_width_0_height_0__pin_16_(cby_1__1__109_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__109_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__109_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__109_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__109_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__109_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__109_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__109_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__109_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__109_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__109_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__109_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__109_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__109_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__109_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__109_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__97_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_109_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_109_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_109_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_109_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_109_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_109_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_109_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_109_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_109_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_109_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_109_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_109_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_109_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_109_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_109_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_109_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_109_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_109_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_109_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_109_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_109_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_109_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_109_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_109_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_109_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_109_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_109_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_109_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_109_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_109_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_109_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_109_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[99]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[99]),
    .ccff_tail(grid_clb_109_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__3_
  (
    .clk_0_N_in(clk_1_wires[181]),
    .prog_clk_0_N_in(prog_clk_1_wires[181]),
    .prog_clk_0_E_out(prog_clk_0_wires[374]),
    .prog_clk_0_S_out(prog_clk_0_wires[373]),
    .Reset_E_out(ResetWires[86]),
    .Reset_W_in(ResetWires[85]),
    .pReset_N_in(pResetWires[198]),
    .Test_en_E_out(Test_enWires[86]),
    .Test_en_W_in(Test_enWires[85]),
    .SC_OUT_TOP(scff_Wires[245]),
    .SC_IN_BOT(scff_Wires[244]),
    .top_width_0_height_0__pin_0_(cbx_1__1__101_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__101_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__101_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__101_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__101_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__101_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__101_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__101_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__101_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__101_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__101_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__101_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__101_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__101_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__101_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__101_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[101]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[101]),
    .right_width_0_height_0__pin_16_(cby_1__1__110_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__110_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__110_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__110_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__110_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__110_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__110_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__110_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__110_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__110_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__110_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__110_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__110_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__110_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__110_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__110_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__98_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_110_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_110_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_110_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_110_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_110_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_110_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_110_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_110_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_110_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_110_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_110_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_110_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_110_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_110_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_110_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_110_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_110_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_110_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_110_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_110_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_110_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_110_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_110_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_110_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_110_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_110_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_110_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_110_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_110_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_110_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_110_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_110_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[100]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[100]),
    .ccff_tail(grid_clb_110_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__4_
  (
    .clk_0_S_in(clk_1_wires[180]),
    .prog_clk_0_S_in(prog_clk_1_wires[180]),
    .prog_clk_0_E_out(prog_clk_0_wires[377]),
    .prog_clk_0_S_out(prog_clk_0_wires[376]),
    .Reset_E_out(ResetWires[108]),
    .Reset_W_in(ResetWires[107]),
    .pReset_N_in(pResetWires[247]),
    .Test_en_E_out(Test_enWires[108]),
    .Test_en_W_in(Test_enWires[107]),
    .SC_OUT_TOP(scff_Wires[247]),
    .SC_IN_BOT(scff_Wires[246]),
    .top_width_0_height_0__pin_0_(cbx_1__1__102_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__102_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__102_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__102_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__102_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__102_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__102_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__102_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__102_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__102_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__102_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__102_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__102_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__102_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__102_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__102_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[102]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[102]),
    .right_width_0_height_0__pin_16_(cby_1__1__111_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__111_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__111_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__111_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__111_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__111_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__111_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__111_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__111_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__111_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__111_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__111_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__111_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__111_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__111_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__111_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__99_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_111_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_111_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_111_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_111_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_111_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_111_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_111_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_111_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_111_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_111_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_111_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_111_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_111_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_111_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_111_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_111_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_111_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_111_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_111_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_111_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_111_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_111_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_111_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_111_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_111_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_111_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_111_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_111_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_111_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_111_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_111_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_111_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[101]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[101]),
    .ccff_tail(grid_clb_111_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__5_
  (
    .clk_0_N_in(clk_1_wires[188]),
    .prog_clk_0_N_in(prog_clk_1_wires[188]),
    .prog_clk_0_E_out(prog_clk_0_wires[380]),
    .prog_clk_0_S_out(prog_clk_0_wires[379]),
    .Reset_E_out(ResetWires[130]),
    .Reset_W_in(ResetWires[129]),
    .pReset_N_in(pResetWires[296]),
    .Test_en_E_out(Test_enWires[130]),
    .Test_en_W_in(Test_enWires[129]),
    .SC_OUT_TOP(scff_Wires[249]),
    .SC_IN_BOT(scff_Wires[248]),
    .top_width_0_height_0__pin_0_(cbx_1__1__103_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__103_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__103_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__103_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__103_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__103_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__103_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__103_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__103_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__103_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__103_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__103_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__103_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__103_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__103_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__103_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[103]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[103]),
    .right_width_0_height_0__pin_16_(cby_1__1__112_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__112_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__112_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__112_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__112_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__112_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__112_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__112_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__112_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__112_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__112_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__112_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__112_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__112_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__112_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__112_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__100_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_112_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_112_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_112_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_112_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_112_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_112_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_112_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_112_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_112_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_112_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_112_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_112_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_112_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_112_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_112_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_112_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_112_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_112_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_112_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_112_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_112_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_112_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_112_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_112_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_112_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_112_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_112_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_112_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_112_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_112_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_112_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_112_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[102]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[102]),
    .ccff_tail(grid_clb_112_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__6_
  (
    .clk_0_S_in(clk_1_wires[187]),
    .prog_clk_0_S_in(prog_clk_1_wires[187]),
    .prog_clk_0_E_out(prog_clk_0_wires[383]),
    .prog_clk_0_S_out(prog_clk_0_wires[382]),
    .Reset_E_out(ResetWires[152]),
    .Reset_W_in(ResetWires[151]),
    .pReset_N_in(pResetWires[345]),
    .Test_en_E_out(Test_enWires[152]),
    .Test_en_W_in(Test_enWires[151]),
    .SC_OUT_TOP(scff_Wires[251]),
    .SC_IN_BOT(scff_Wires[250]),
    .top_width_0_height_0__pin_0_(cbx_1__1__104_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__104_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__104_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__104_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__104_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__104_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__104_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__104_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__104_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__104_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__104_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__104_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__104_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__104_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__104_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__104_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[104]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[104]),
    .right_width_0_height_0__pin_16_(cby_1__1__113_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__113_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__113_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__113_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__113_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__113_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__113_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__113_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__113_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__113_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__113_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__113_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__113_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__113_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__113_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__113_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__101_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_113_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_113_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_113_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_113_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_113_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_113_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_113_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_113_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_113_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_113_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_113_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_113_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_113_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_113_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_113_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_113_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_113_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_113_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_113_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_113_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_113_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_113_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_113_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_113_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_113_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_113_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_113_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_113_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_113_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_113_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_113_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_113_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[103]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[103]),
    .ccff_tail(grid_clb_113_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__7_
  (
    .clk_0_N_in(clk_1_wires[195]),
    .prog_clk_0_N_in(prog_clk_1_wires[195]),
    .prog_clk_0_E_out(prog_clk_0_wires[386]),
    .prog_clk_0_S_out(prog_clk_0_wires[385]),
    .Reset_E_out(ResetWires[174]),
    .Reset_W_in(ResetWires[173]),
    .pReset_N_in(pResetWires[394]),
    .Test_en_E_out(Test_enWires[174]),
    .Test_en_W_in(Test_enWires[173]),
    .SC_OUT_TOP(scff_Wires[253]),
    .SC_IN_BOT(scff_Wires[252]),
    .top_width_0_height_0__pin_0_(cbx_1__1__105_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__105_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__105_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__105_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__105_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__105_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__105_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__105_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__105_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__105_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__105_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__105_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__105_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__105_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__105_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__105_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[105]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[105]),
    .right_width_0_height_0__pin_16_(cby_1__1__114_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__114_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__114_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__114_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__114_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__114_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__114_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__114_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__114_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__114_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__114_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__114_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__114_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__114_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__114_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__114_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__102_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_114_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_114_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_114_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_114_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_114_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_114_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_114_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_114_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_114_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_114_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_114_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_114_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_114_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_114_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_114_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_114_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_114_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_114_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_114_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_114_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_114_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_114_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_114_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_114_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_114_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_114_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_114_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_114_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_114_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_114_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_114_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_114_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[104]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[104]),
    .ccff_tail(grid_clb_114_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__8_
  (
    .clk_0_S_in(clk_1_wires[194]),
    .prog_clk_0_S_in(prog_clk_1_wires[194]),
    .prog_clk_0_E_out(prog_clk_0_wires[389]),
    .prog_clk_0_S_out(prog_clk_0_wires[388]),
    .Reset_E_out(ResetWires[196]),
    .Reset_W_in(ResetWires[195]),
    .pReset_N_in(pResetWires[443]),
    .Test_en_E_out(Test_enWires[196]),
    .Test_en_W_in(Test_enWires[195]),
    .SC_OUT_TOP(scff_Wires[255]),
    .SC_IN_BOT(scff_Wires[254]),
    .top_width_0_height_0__pin_0_(cbx_1__1__106_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__106_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__106_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__106_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__106_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__106_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__106_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__106_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__106_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__106_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__106_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__106_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__106_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__106_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__106_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__106_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[106]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[106]),
    .right_width_0_height_0__pin_16_(cby_1__1__115_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__115_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__115_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__115_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__115_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__115_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__115_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__115_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__115_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__115_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__115_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__115_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__115_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__115_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__115_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__115_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__103_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_115_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_115_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_115_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_115_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_115_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_115_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_115_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_115_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_115_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_115_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_115_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_115_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_115_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_115_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_115_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_115_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_115_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_115_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_115_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_115_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_115_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_115_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_115_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_115_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_115_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_115_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_115_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_115_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_115_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_115_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_115_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_115_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[105]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[105]),
    .ccff_tail(grid_clb_115_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__9_
  (
    .clk_0_N_in(clk_1_wires[202]),
    .prog_clk_0_N_in(prog_clk_1_wires[202]),
    .prog_clk_0_E_out(prog_clk_0_wires[392]),
    .prog_clk_0_S_out(prog_clk_0_wires[391]),
    .Reset_E_out(ResetWires[218]),
    .Reset_W_in(ResetWires[217]),
    .pReset_N_in(pResetWires[492]),
    .Test_en_E_out(Test_enWires[218]),
    .Test_en_W_in(Test_enWires[217]),
    .SC_OUT_TOP(scff_Wires[257]),
    .SC_IN_BOT(scff_Wires[256]),
    .top_width_0_height_0__pin_0_(cbx_1__1__107_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__107_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__107_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__107_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__107_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__107_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__107_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__107_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__107_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__107_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__107_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__107_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__107_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__107_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__107_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__107_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[107]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[107]),
    .right_width_0_height_0__pin_16_(cby_1__1__116_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__116_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__116_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__116_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__116_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__116_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__116_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__116_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__116_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__116_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__116_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__116_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__116_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__116_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__116_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__116_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__104_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_116_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_116_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_116_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_116_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_116_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_116_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_116_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_116_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_116_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_116_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_116_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_116_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_116_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_116_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_116_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_116_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_116_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_116_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_116_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_116_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_116_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_116_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_116_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_116_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_116_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_116_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_116_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_116_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_116_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_116_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_116_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_116_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[106]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[106]),
    .ccff_tail(grid_clb_116_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__10_
  (
    .clk_0_S_in(clk_1_wires[201]),
    .prog_clk_0_S_in(prog_clk_1_wires[201]),
    .prog_clk_0_E_out(prog_clk_0_wires[395]),
    .prog_clk_0_S_out(prog_clk_0_wires[394]),
    .Reset_E_out(ResetWires[240]),
    .Reset_W_in(ResetWires[239]),
    .pReset_N_in(pResetWires[541]),
    .Test_en_E_out(Test_enWires[240]),
    .Test_en_W_in(Test_enWires[239]),
    .SC_OUT_TOP(scff_Wires[259]),
    .SC_IN_BOT(scff_Wires[258]),
    .top_width_0_height_0__pin_0_(cbx_1__1__108_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__108_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__108_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__108_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__108_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__108_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__108_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__108_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__108_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__108_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__108_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__108_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__108_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__108_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__108_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__108_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[108]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[108]),
    .right_width_0_height_0__pin_16_(cby_1__1__117_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__117_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__117_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__117_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__117_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__117_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__117_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__117_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__117_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__117_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__117_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__117_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__117_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__117_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__117_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__117_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__105_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_117_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_117_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_117_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_117_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_117_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_117_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_117_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_117_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_117_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_117_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_117_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_117_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_117_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_117_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_117_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_117_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_117_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_117_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_117_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_117_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_117_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_117_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_117_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_117_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_117_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_117_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_117_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_117_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_117_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_117_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_117_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_117_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[107]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[107]),
    .ccff_tail(grid_clb_117_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__11_
  (
    .clk_0_N_in(clk_1_wires[209]),
    .prog_clk_0_N_in(prog_clk_1_wires[209]),
    .prog_clk_0_E_out(prog_clk_0_wires[398]),
    .prog_clk_0_S_out(prog_clk_0_wires[397]),
    .Reset_E_out(ResetWires[262]),
    .Reset_W_in(ResetWires[261]),
    .pReset_N_in(pResetWires[590]),
    .Test_en_E_out(Test_enWires[262]),
    .Test_en_W_in(Test_enWires[261]),
    .SC_OUT_TOP(scff_Wires[261]),
    .SC_IN_BOT(scff_Wires[260]),
    .top_width_0_height_0__pin_0_(cbx_1__1__109_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__109_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__109_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__109_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__109_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__109_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__109_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__109_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__109_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__109_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__109_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__109_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__109_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__109_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__109_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__109_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[109]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[109]),
    .right_width_0_height_0__pin_16_(cby_1__1__118_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__118_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__118_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__118_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__118_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__118_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__118_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__118_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__118_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__118_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__118_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__118_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__118_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__118_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__118_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__118_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__106_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_118_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_118_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_118_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_118_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_118_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_118_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_118_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_118_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_118_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_118_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_118_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_118_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_118_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_118_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_118_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_118_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_118_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_118_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_118_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_118_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_118_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_118_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_118_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_118_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_118_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_118_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_118_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_118_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_118_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_118_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_118_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_118_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[108]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[108]),
    .ccff_tail(grid_clb_118_ccff_tail[0])
  );


  grid_clb
  grid_clb_10__12_
  (
    .clk_0_S_in(clk_1_wires[208]),
    .prog_clk_0_S_in(prog_clk_1_wires[208]),
    .prog_clk_0_N_out(prog_clk_0_wires[403]),
    .prog_clk_0_E_out(prog_clk_0_wires[401]),
    .prog_clk_0_S_out(prog_clk_0_wires[400]),
    .Reset_E_out(ResetWires[284]),
    .Reset_W_in(ResetWires[283]),
    .pReset_N_in(pResetWires[630]),
    .Test_en_E_out(Test_enWires[284]),
    .Test_en_W_in(Test_enWires[283]),
    .SC_OUT_TOP(scff_Wires[263]),
    .SC_IN_BOT(scff_Wires[262]),
    .top_width_0_height_0__pin_0_(cbx_1__12__9_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__9_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__9_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__9_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__9_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__9_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__9_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__9_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__9_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__9_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__9_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__9_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__9_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__9_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__9_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__9_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_10__12__undriven_top_width_0_height_0__pin_32_[0]),
    .top_width_0_height_0__pin_34_(grid_clb_10__12__undriven_top_width_0_height_0__pin_34_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__119_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__119_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__119_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__119_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__119_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__119_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__119_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__119_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__119_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__119_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__119_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__119_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__119_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__119_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__119_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__119_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__107_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_119_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_119_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_119_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_119_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_119_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_119_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_119_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_119_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_119_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_119_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_119_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_119_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_119_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_119_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_119_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_119_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_119_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_119_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_119_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_119_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_119_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_119_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_119_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_119_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_119_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_119_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_119_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_119_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_119_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_119_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_119_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_119_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[109]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[109]),
    .ccff_tail(grid_clb_119_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__1_
  (
    .clk_0_N_in(clk_1_wires[214]),
    .prog_clk_0_N_in(prog_clk_1_wires[214]),
    .prog_clk_0_E_out(prog_clk_0_wires[406]),
    .prog_clk_0_S_out(prog_clk_0_wires[405]),
    .Reset_E_out(ResetWires[44]),
    .Reset_W_in(ResetWires[43]),
    .pReset_N_in(pResetWires[104]),
    .Test_en_E_out(Test_enWires[44]),
    .Test_en_W_in(Test_enWires[43]),
    .SC_OUT_BOT(scff_Wires[290]),
    .SC_IN_TOP(scff_Wires[288]),
    .top_width_0_height_0__pin_0_(cbx_1__1__110_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__110_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__110_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__110_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__110_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__110_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__110_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__110_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__110_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__110_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__110_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__110_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__110_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__110_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__110_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__110_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[110]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[110]),
    .right_width_0_height_0__pin_16_(cby_1__1__120_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__120_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__120_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__120_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__120_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__120_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__120_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__120_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__120_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__120_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__120_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__120_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__120_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__120_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__120_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__120_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__108_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_120_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_120_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_120_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_120_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_120_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_120_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_120_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_120_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_120_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_120_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_120_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_120_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_120_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_120_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_120_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_120_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_120_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_120_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_120_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_120_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_120_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_120_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_120_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_120_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_120_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_120_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_120_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_120_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_120_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_120_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_120_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_120_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(grid_clb_11__1__undriven_bottom_width_0_height_0__pin_52_[0]),
    .bottom_width_0_height_0__pin_54_(grid_clb_11__1__undriven_bottom_width_0_height_0__pin_54_[0]),
    .ccff_tail(grid_clb_120_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__2_
  (
    .clk_0_S_in(clk_1_wires[213]),
    .prog_clk_0_S_in(prog_clk_1_wires[213]),
    .prog_clk_0_E_out(prog_clk_0_wires[409]),
    .prog_clk_0_S_out(prog_clk_0_wires[408]),
    .Reset_E_out(ResetWires[66]),
    .Reset_W_in(ResetWires[65]),
    .pReset_N_in(pResetWires[153]),
    .Test_en_E_out(Test_enWires[66]),
    .Test_en_W_in(Test_enWires[65]),
    .SC_OUT_BOT(scff_Wires[287]),
    .SC_IN_TOP(scff_Wires[286]),
    .top_width_0_height_0__pin_0_(cbx_1__1__111_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__111_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__111_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__111_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__111_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__111_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__111_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__111_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__111_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__111_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__111_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__111_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__111_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__111_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__111_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__111_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[111]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[111]),
    .right_width_0_height_0__pin_16_(cby_1__1__121_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__121_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__121_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__121_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__121_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__121_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__121_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__121_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__121_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__121_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__121_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__121_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__121_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__121_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__121_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__121_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__109_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_121_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_121_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_121_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_121_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_121_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_121_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_121_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_121_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_121_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_121_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_121_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_121_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_121_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_121_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_121_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_121_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_121_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_121_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_121_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_121_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_121_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_121_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_121_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_121_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_121_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_121_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_121_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_121_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_121_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_121_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_121_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_121_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[110]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[110]),
    .ccff_tail(grid_clb_121_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__3_
  (
    .clk_0_N_in(clk_1_wires[221]),
    .prog_clk_0_N_in(prog_clk_1_wires[221]),
    .prog_clk_0_E_out(prog_clk_0_wires[412]),
    .prog_clk_0_S_out(prog_clk_0_wires[411]),
    .Reset_E_out(ResetWires[88]),
    .Reset_W_in(ResetWires[87]),
    .pReset_N_in(pResetWires[202]),
    .Test_en_E_out(Test_enWires[88]),
    .Test_en_W_in(Test_enWires[87]),
    .SC_OUT_BOT(scff_Wires[285]),
    .SC_IN_TOP(scff_Wires[284]),
    .top_width_0_height_0__pin_0_(cbx_1__1__112_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__112_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__112_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__112_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__112_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__112_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__112_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__112_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__112_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__112_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__112_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__112_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__112_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__112_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__112_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__112_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[112]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[112]),
    .right_width_0_height_0__pin_16_(cby_1__1__122_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__122_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__122_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__122_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__122_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__122_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__122_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__122_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__122_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__122_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__122_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__122_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__122_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__122_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__122_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__122_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__110_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_122_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_122_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_122_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_122_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_122_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_122_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_122_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_122_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_122_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_122_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_122_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_122_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_122_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_122_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_122_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_122_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_122_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_122_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_122_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_122_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_122_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_122_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_122_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_122_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_122_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_122_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_122_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_122_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_122_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_122_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_122_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_122_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[111]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[111]),
    .ccff_tail(grid_clb_122_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__4_
  (
    .clk_0_S_in(clk_1_wires[220]),
    .prog_clk_0_S_in(prog_clk_1_wires[220]),
    .prog_clk_0_E_out(prog_clk_0_wires[415]),
    .prog_clk_0_S_out(prog_clk_0_wires[414]),
    .Reset_E_out(ResetWires[110]),
    .Reset_W_in(ResetWires[109]),
    .pReset_N_in(pResetWires[251]),
    .Test_en_E_out(Test_enWires[110]),
    .Test_en_W_in(Test_enWires[109]),
    .SC_OUT_BOT(scff_Wires[283]),
    .SC_IN_TOP(scff_Wires[282]),
    .top_width_0_height_0__pin_0_(cbx_1__1__113_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__113_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__113_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__113_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__113_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__113_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__113_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__113_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__113_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__113_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__113_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__113_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__113_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__113_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__113_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__113_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[113]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[113]),
    .right_width_0_height_0__pin_16_(cby_1__1__123_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__123_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__123_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__123_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__123_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__123_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__123_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__123_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__123_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__123_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__123_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__123_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__123_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__123_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__123_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__123_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__111_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_123_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_123_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_123_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_123_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_123_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_123_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_123_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_123_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_123_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_123_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_123_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_123_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_123_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_123_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_123_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_123_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_123_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_123_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_123_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_123_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_123_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_123_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_123_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_123_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_123_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_123_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_123_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_123_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_123_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_123_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_123_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_123_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[112]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[112]),
    .ccff_tail(grid_clb_123_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__5_
  (
    .clk_0_N_in(clk_1_wires[228]),
    .prog_clk_0_N_in(prog_clk_1_wires[228]),
    .prog_clk_0_E_out(prog_clk_0_wires[418]),
    .prog_clk_0_S_out(prog_clk_0_wires[417]),
    .Reset_E_out(ResetWires[132]),
    .Reset_W_in(ResetWires[131]),
    .pReset_N_in(pResetWires[300]),
    .Test_en_E_out(Test_enWires[132]),
    .Test_en_W_in(Test_enWires[131]),
    .SC_OUT_BOT(scff_Wires[281]),
    .SC_IN_TOP(scff_Wires[280]),
    .top_width_0_height_0__pin_0_(cbx_1__1__114_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__114_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__114_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__114_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__114_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__114_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__114_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__114_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__114_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__114_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__114_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__114_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__114_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__114_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__114_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__114_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[114]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[114]),
    .right_width_0_height_0__pin_16_(cby_1__1__124_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__124_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__124_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__124_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__124_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__124_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__124_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__124_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__124_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__124_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__124_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__124_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__124_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__124_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__124_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__124_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__112_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_124_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_124_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_124_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_124_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_124_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_124_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_124_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_124_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_124_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_124_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_124_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_124_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_124_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_124_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_124_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_124_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_124_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_124_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_124_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_124_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_124_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_124_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_124_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_124_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_124_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_124_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_124_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_124_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_124_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_124_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_124_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_124_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[113]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[113]),
    .ccff_tail(grid_clb_124_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__6_
  (
    .clk_0_S_in(clk_1_wires[227]),
    .prog_clk_0_S_in(prog_clk_1_wires[227]),
    .prog_clk_0_E_out(prog_clk_0_wires[421]),
    .prog_clk_0_S_out(prog_clk_0_wires[420]),
    .Reset_E_out(ResetWires[154]),
    .Reset_W_in(ResetWires[153]),
    .pReset_N_in(pResetWires[349]),
    .Test_en_E_out(Test_enWires[154]),
    .Test_en_W_in(Test_enWires[153]),
    .SC_OUT_BOT(scff_Wires[279]),
    .SC_IN_TOP(scff_Wires[278]),
    .top_width_0_height_0__pin_0_(cbx_1__1__115_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__115_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__115_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__115_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__115_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__115_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__115_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__115_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__115_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__115_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__115_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__115_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__115_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__115_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__115_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__115_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[115]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[115]),
    .right_width_0_height_0__pin_16_(cby_1__1__125_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__125_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__125_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__125_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__125_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__125_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__125_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__125_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__125_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__125_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__125_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__125_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__125_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__125_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__125_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__125_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__113_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_125_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_125_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_125_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_125_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_125_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_125_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_125_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_125_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_125_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_125_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_125_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_125_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_125_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_125_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_125_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_125_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_125_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_125_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_125_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_125_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_125_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_125_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_125_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_125_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_125_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_125_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_125_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_125_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_125_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_125_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_125_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_125_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[114]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[114]),
    .ccff_tail(grid_clb_125_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__7_
  (
    .clk_0_N_in(clk_1_wires[235]),
    .prog_clk_0_N_in(prog_clk_1_wires[235]),
    .prog_clk_0_E_out(prog_clk_0_wires[424]),
    .prog_clk_0_S_out(prog_clk_0_wires[423]),
    .Reset_E_out(ResetWires[176]),
    .Reset_W_in(ResetWires[175]),
    .pReset_N_in(pResetWires[398]),
    .Test_en_E_out(Test_enWires[176]),
    .Test_en_W_in(Test_enWires[175]),
    .SC_OUT_BOT(scff_Wires[277]),
    .SC_IN_TOP(scff_Wires[276]),
    .top_width_0_height_0__pin_0_(cbx_1__1__116_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__116_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__116_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__116_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__116_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__116_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__116_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__116_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__116_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__116_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__116_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__116_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__116_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__116_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__116_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__116_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[116]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[116]),
    .right_width_0_height_0__pin_16_(cby_1__1__126_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__126_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__126_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__126_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__126_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__126_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__126_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__126_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__126_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__126_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__126_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__126_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__126_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__126_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__126_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__126_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__114_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_126_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_126_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_126_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_126_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_126_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_126_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_126_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_126_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_126_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_126_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_126_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_126_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_126_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_126_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_126_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_126_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_126_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_126_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_126_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_126_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_126_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_126_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_126_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_126_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_126_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_126_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_126_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_126_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_126_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_126_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_126_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_126_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[115]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[115]),
    .ccff_tail(grid_clb_126_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__8_
  (
    .clk_0_S_in(clk_1_wires[234]),
    .prog_clk_0_S_in(prog_clk_1_wires[234]),
    .prog_clk_0_E_out(prog_clk_0_wires[427]),
    .prog_clk_0_S_out(prog_clk_0_wires[426]),
    .Reset_E_out(ResetWires[198]),
    .Reset_W_in(ResetWires[197]),
    .pReset_N_in(pResetWires[447]),
    .Test_en_E_out(Test_enWires[198]),
    .Test_en_W_in(Test_enWires[197]),
    .SC_OUT_BOT(scff_Wires[275]),
    .SC_IN_TOP(scff_Wires[274]),
    .top_width_0_height_0__pin_0_(cbx_1__1__117_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__117_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__117_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__117_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__117_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__117_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__117_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__117_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__117_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__117_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__117_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__117_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__117_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__117_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__117_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__117_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[117]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[117]),
    .right_width_0_height_0__pin_16_(cby_1__1__127_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__127_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__127_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__127_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__127_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__127_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__127_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__127_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__127_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__127_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__127_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__127_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__127_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__127_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__127_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__127_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__115_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_127_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_127_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_127_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_127_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_127_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_127_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_127_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_127_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_127_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_127_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_127_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_127_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_127_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_127_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_127_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_127_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_127_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_127_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_127_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_127_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_127_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_127_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_127_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_127_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_127_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_127_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_127_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_127_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_127_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_127_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_127_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_127_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[116]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[116]),
    .ccff_tail(grid_clb_127_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__9_
  (
    .clk_0_N_in(clk_1_wires[242]),
    .prog_clk_0_N_in(prog_clk_1_wires[242]),
    .prog_clk_0_E_out(prog_clk_0_wires[430]),
    .prog_clk_0_S_out(prog_clk_0_wires[429]),
    .Reset_E_out(ResetWires[220]),
    .Reset_W_in(ResetWires[219]),
    .pReset_N_in(pResetWires[496]),
    .Test_en_E_out(Test_enWires[220]),
    .Test_en_W_in(Test_enWires[219]),
    .SC_OUT_BOT(scff_Wires[273]),
    .SC_IN_TOP(scff_Wires[272]),
    .top_width_0_height_0__pin_0_(cbx_1__1__118_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__118_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__118_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__118_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__118_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__118_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__118_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__118_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__118_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__118_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__118_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__118_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__118_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__118_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__118_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__118_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[118]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[118]),
    .right_width_0_height_0__pin_16_(cby_1__1__128_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__128_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__128_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__128_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__128_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__128_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__128_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__128_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__128_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__128_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__128_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__128_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__128_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__128_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__128_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__128_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__116_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_128_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_128_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_128_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_128_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_128_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_128_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_128_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_128_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_128_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_128_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_128_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_128_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_128_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_128_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_128_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_128_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_128_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_128_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_128_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_128_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_128_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_128_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_128_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_128_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_128_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_128_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_128_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_128_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_128_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_128_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_128_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_128_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[117]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[117]),
    .ccff_tail(grid_clb_128_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__10_
  (
    .clk_0_S_in(clk_1_wires[241]),
    .prog_clk_0_S_in(prog_clk_1_wires[241]),
    .prog_clk_0_E_out(prog_clk_0_wires[433]),
    .prog_clk_0_S_out(prog_clk_0_wires[432]),
    .Reset_E_out(ResetWires[242]),
    .Reset_W_in(ResetWires[241]),
    .pReset_N_in(pResetWires[545]),
    .Test_en_E_out(Test_enWires[242]),
    .Test_en_W_in(Test_enWires[241]),
    .SC_OUT_BOT(scff_Wires[271]),
    .SC_IN_TOP(scff_Wires[270]),
    .top_width_0_height_0__pin_0_(cbx_1__1__119_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__119_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__119_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__119_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__119_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__119_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__119_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__119_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__119_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__119_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__119_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__119_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__119_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__119_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__119_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__119_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[119]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[119]),
    .right_width_0_height_0__pin_16_(cby_1__1__129_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__129_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__129_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__129_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__129_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__129_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__129_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__129_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__129_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__129_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__129_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__129_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__129_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__129_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__129_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__129_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__117_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_129_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_129_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_129_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_129_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_129_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_129_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_129_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_129_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_129_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_129_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_129_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_129_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_129_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_129_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_129_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_129_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_129_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_129_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_129_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_129_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_129_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_129_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_129_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_129_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_129_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_129_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_129_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_129_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_129_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_129_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_129_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_129_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[118]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[118]),
    .ccff_tail(grid_clb_129_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__11_
  (
    .clk_0_N_in(clk_1_wires[249]),
    .prog_clk_0_N_in(prog_clk_1_wires[249]),
    .prog_clk_0_E_out(prog_clk_0_wires[436]),
    .prog_clk_0_S_out(prog_clk_0_wires[435]),
    .Reset_E_out(ResetWires[264]),
    .Reset_W_in(ResetWires[263]),
    .pReset_N_in(pResetWires[594]),
    .Test_en_E_out(Test_enWires[264]),
    .Test_en_W_in(Test_enWires[263]),
    .SC_OUT_BOT(scff_Wires[269]),
    .SC_IN_TOP(scff_Wires[268]),
    .top_width_0_height_0__pin_0_(cbx_1__1__120_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__120_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__120_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__120_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__120_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__120_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__120_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__120_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__120_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__120_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__120_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__120_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__120_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__120_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__120_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__120_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[120]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[120]),
    .right_width_0_height_0__pin_16_(cby_1__1__130_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__130_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__130_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__130_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__130_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__130_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__130_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__130_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__130_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__130_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__130_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__130_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__130_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__130_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__130_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__130_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__118_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_130_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_130_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_130_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_130_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_130_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_130_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_130_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_130_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_130_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_130_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_130_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_130_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_130_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_130_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_130_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_130_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_130_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_130_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_130_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_130_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_130_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_130_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_130_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_130_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_130_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_130_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_130_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_130_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_130_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_130_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_130_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_130_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[119]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[119]),
    .ccff_tail(grid_clb_130_ccff_tail[0])
  );


  grid_clb
  grid_clb_11__12_
  (
    .clk_0_S_in(clk_1_wires[248]),
    .prog_clk_0_S_in(prog_clk_1_wires[248]),
    .prog_clk_0_N_out(prog_clk_0_wires[441]),
    .prog_clk_0_E_out(prog_clk_0_wires[439]),
    .prog_clk_0_S_out(prog_clk_0_wires[438]),
    .Reset_E_out(ResetWires[286]),
    .Reset_W_in(ResetWires[285]),
    .pReset_N_in(pResetWires[633]),
    .Test_en_E_out(Test_enWires[286]),
    .Test_en_W_in(Test_enWires[285]),
    .SC_OUT_BOT(scff_Wires[267]),
    .SC_IN_TOP(scff_Wires[266]),
    .top_width_0_height_0__pin_0_(cbx_1__12__10_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__10_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__10_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__10_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__10_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__10_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__10_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__10_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__10_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__10_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__10_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__10_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__10_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__10_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__10_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__10_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_11__12__undriven_top_width_0_height_0__pin_32_[0]),
    .top_width_0_height_0__pin_34_(grid_clb_11__12__undriven_top_width_0_height_0__pin_34_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__131_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__131_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__131_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__131_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__131_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__131_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__131_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__131_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__131_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__131_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__131_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__131_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__131_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__131_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__131_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__131_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__119_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_131_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_131_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_131_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_131_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_131_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_131_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_131_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_131_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_131_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_131_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_131_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_131_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_131_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_131_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_131_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_131_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_131_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_131_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_131_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_131_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_131_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_131_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_131_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_131_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_131_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_131_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_131_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_131_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_131_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_131_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_131_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_131_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[120]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[120]),
    .ccff_tail(grid_clb_131_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__1_
  (
    .clk_0_N_in(clk_1_wires[216]),
    .prog_clk_0_N_in(prog_clk_1_wires[216]),
    .prog_clk_0_E_out(prog_clk_0_wires[444]),
    .prog_clk_0_S_out(prog_clk_0_wires[443]),
    .Reset_W_in(ResetWires[45]),
    .pReset_N_in(pResetWires[108]),
    .Test_en_W_in(Test_enWires[45]),
    .SC_OUT_TOP(scff_Wires[294]),
    .SC_IN_BOT(scff_Wires[293]),
    .top_width_0_height_0__pin_0_(cbx_1__1__121_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__121_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__121_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__121_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__121_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__121_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__121_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__121_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__121_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__121_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__121_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__121_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__121_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__121_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__121_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__121_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[121]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[121]),
    .right_width_0_height_0__pin_16_(cby_12__1__0_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__0_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__0_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__0_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__0_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__0_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__0_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__0_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__0_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__0_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__0_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__0_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__0_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__0_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__0_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__0_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__120_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_132_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_132_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_132_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_132_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_132_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_132_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_132_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_132_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_132_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_132_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_132_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_132_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_132_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_132_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_132_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_132_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_132_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_132_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_132_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_132_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_132_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_132_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_132_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_132_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_132_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_132_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_132_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_132_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_132_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_132_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_132_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_132_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(grid_clb_12__1__undriven_bottom_width_0_height_0__pin_52_[0]),
    .bottom_width_0_height_0__pin_54_(grid_clb_12__1__undriven_bottom_width_0_height_0__pin_54_[0]),
    .ccff_tail(grid_clb_132_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__2_
  (
    .clk_0_S_in(clk_1_wires[215]),
    .prog_clk_0_S_in(prog_clk_1_wires[215]),
    .prog_clk_0_E_out(prog_clk_0_wires[447]),
    .prog_clk_0_S_out(prog_clk_0_wires[446]),
    .Reset_W_in(ResetWires[67]),
    .pReset_N_in(pResetWires[157]),
    .Test_en_W_in(Test_enWires[67]),
    .SC_OUT_TOP(scff_Wires[296]),
    .SC_IN_BOT(scff_Wires[295]),
    .top_width_0_height_0__pin_0_(cbx_1__1__122_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__122_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__122_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__122_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__122_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__122_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__122_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__122_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__122_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__122_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__122_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__122_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__122_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__122_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__122_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__122_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[122]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[122]),
    .right_width_0_height_0__pin_16_(cby_12__1__1_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__1_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__1_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__1_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__1_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__1_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__1_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__1_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__1_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__1_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__1_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__1_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__1_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__1_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__1_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__1_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__121_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_133_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_133_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_133_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_133_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_133_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_133_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_133_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_133_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_133_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_133_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_133_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_133_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_133_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_133_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_133_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_133_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_133_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_133_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_133_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_133_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_133_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_133_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_133_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_133_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_133_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_133_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_133_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_133_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_133_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_133_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_133_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_133_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[121]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[121]),
    .ccff_tail(grid_clb_133_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__3_
  (
    .clk_0_N_in(clk_1_wires[223]),
    .prog_clk_0_N_in(prog_clk_1_wires[223]),
    .prog_clk_0_E_out(prog_clk_0_wires[450]),
    .prog_clk_0_S_out(prog_clk_0_wires[449]),
    .Reset_W_in(ResetWires[89]),
    .pReset_N_in(pResetWires[206]),
    .Test_en_W_in(Test_enWires[89]),
    .SC_OUT_TOP(scff_Wires[298]),
    .SC_IN_BOT(scff_Wires[297]),
    .top_width_0_height_0__pin_0_(cbx_1__1__123_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__123_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__123_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__123_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__123_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__123_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__123_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__123_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__123_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__123_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__123_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__123_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__123_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__123_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__123_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__123_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[123]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[123]),
    .right_width_0_height_0__pin_16_(cby_12__1__2_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__2_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__2_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__2_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__2_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__2_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__2_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__2_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__2_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__2_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__2_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__2_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__2_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__2_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__2_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__2_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__122_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_134_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_134_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_134_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_134_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_134_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_134_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_134_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_134_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_134_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_134_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_134_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_134_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_134_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_134_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_134_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_134_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_134_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_134_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_134_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_134_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_134_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_134_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_134_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_134_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_134_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_134_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_134_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_134_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_134_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_134_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_134_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_134_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[122]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[122]),
    .ccff_tail(grid_clb_134_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__4_
  (
    .clk_0_S_in(clk_1_wires[222]),
    .prog_clk_0_S_in(prog_clk_1_wires[222]),
    .prog_clk_0_E_out(prog_clk_0_wires[453]),
    .prog_clk_0_S_out(prog_clk_0_wires[452]),
    .Reset_W_in(ResetWires[111]),
    .pReset_N_in(pResetWires[255]),
    .Test_en_W_in(Test_enWires[111]),
    .SC_OUT_TOP(scff_Wires[300]),
    .SC_IN_BOT(scff_Wires[299]),
    .top_width_0_height_0__pin_0_(cbx_1__1__124_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__124_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__124_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__124_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__124_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__124_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__124_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__124_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__124_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__124_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__124_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__124_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__124_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__124_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__124_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__124_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[124]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[124]),
    .right_width_0_height_0__pin_16_(cby_12__1__3_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__3_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__3_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__3_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__3_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__3_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__3_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__3_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__3_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__3_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__3_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__3_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__3_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__3_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__3_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__3_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__123_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_135_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_135_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_135_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_135_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_135_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_135_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_135_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_135_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_135_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_135_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_135_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_135_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_135_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_135_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_135_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_135_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_135_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_135_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_135_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_135_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_135_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_135_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_135_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_135_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_135_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_135_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_135_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_135_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_135_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_135_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_135_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_135_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[123]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[123]),
    .ccff_tail(grid_clb_135_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__5_
  (
    .clk_0_N_in(clk_1_wires[230]),
    .prog_clk_0_N_in(prog_clk_1_wires[230]),
    .prog_clk_0_E_out(prog_clk_0_wires[456]),
    .prog_clk_0_S_out(prog_clk_0_wires[455]),
    .Reset_W_in(ResetWires[133]),
    .pReset_N_in(pResetWires[304]),
    .Test_en_W_in(Test_enWires[133]),
    .SC_OUT_TOP(scff_Wires[302]),
    .SC_IN_BOT(scff_Wires[301]),
    .top_width_0_height_0__pin_0_(cbx_1__1__125_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__125_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__125_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__125_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__125_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__125_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__125_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__125_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__125_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__125_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__125_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__125_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__125_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__125_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__125_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__125_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[125]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[125]),
    .right_width_0_height_0__pin_16_(cby_12__1__4_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__4_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__4_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__4_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__4_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__4_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__4_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__4_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__4_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__4_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__4_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__4_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__4_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__4_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__4_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__4_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__124_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_136_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_136_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_136_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_136_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_136_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_136_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_136_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_136_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_136_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_136_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_136_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_136_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_136_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_136_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_136_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_136_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_136_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_136_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_136_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_136_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_136_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_136_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_136_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_136_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_136_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_136_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_136_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_136_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_136_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_136_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_136_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_136_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[124]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[124]),
    .ccff_tail(grid_clb_136_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__6_
  (
    .clk_0_S_in(clk_1_wires[229]),
    .prog_clk_0_S_in(prog_clk_1_wires[229]),
    .prog_clk_0_E_out(prog_clk_0_wires[459]),
    .prog_clk_0_S_out(prog_clk_0_wires[458]),
    .Reset_W_in(ResetWires[155]),
    .pReset_N_in(pResetWires[353]),
    .Test_en_W_in(Test_enWires[155]),
    .SC_OUT_TOP(scff_Wires[304]),
    .SC_IN_BOT(scff_Wires[303]),
    .top_width_0_height_0__pin_0_(cbx_1__1__126_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__126_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__126_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__126_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__126_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__126_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__126_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__126_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__126_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__126_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__126_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__126_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__126_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__126_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__126_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__126_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[126]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[126]),
    .right_width_0_height_0__pin_16_(cby_12__1__5_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__5_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__5_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__5_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__5_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__5_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__5_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__5_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__5_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__5_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__5_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__5_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__5_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__5_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__5_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__5_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__125_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_137_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_137_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_137_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_137_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_137_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_137_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_137_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_137_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_137_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_137_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_137_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_137_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_137_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_137_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_137_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_137_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_137_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_137_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_137_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_137_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_137_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_137_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_137_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_137_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_137_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_137_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_137_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_137_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_137_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_137_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_137_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_137_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[125]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[125]),
    .ccff_tail(grid_clb_137_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__7_
  (
    .clk_0_N_in(clk_1_wires[237]),
    .prog_clk_0_N_in(prog_clk_1_wires[237]),
    .prog_clk_0_E_out(prog_clk_0_wires[462]),
    .prog_clk_0_S_out(prog_clk_0_wires[461]),
    .Reset_W_in(ResetWires[177]),
    .pReset_N_in(pResetWires[402]),
    .Test_en_W_in(Test_enWires[177]),
    .SC_OUT_TOP(scff_Wires[306]),
    .SC_IN_BOT(scff_Wires[305]),
    .top_width_0_height_0__pin_0_(cbx_1__1__127_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__127_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__127_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__127_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__127_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__127_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__127_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__127_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__127_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__127_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__127_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__127_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__127_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__127_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__127_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__127_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[127]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[127]),
    .right_width_0_height_0__pin_16_(cby_12__1__6_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__6_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__6_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__6_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__6_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__6_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__6_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__6_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__6_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__6_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__6_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__6_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__6_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__6_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__6_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__6_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__126_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_138_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_138_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_138_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_138_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_138_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_138_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_138_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_138_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_138_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_138_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_138_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_138_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_138_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_138_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_138_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_138_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_138_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_138_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_138_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_138_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_138_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_138_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_138_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_138_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_138_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_138_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_138_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_138_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_138_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_138_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_138_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_138_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[126]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[126]),
    .ccff_tail(grid_clb_138_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__8_
  (
    .clk_0_S_in(clk_1_wires[236]),
    .prog_clk_0_S_in(prog_clk_1_wires[236]),
    .prog_clk_0_E_out(prog_clk_0_wires[465]),
    .prog_clk_0_S_out(prog_clk_0_wires[464]),
    .Reset_W_in(ResetWires[199]),
    .pReset_N_in(pResetWires[451]),
    .Test_en_W_in(Test_enWires[199]),
    .SC_OUT_TOP(scff_Wires[308]),
    .SC_IN_BOT(scff_Wires[307]),
    .top_width_0_height_0__pin_0_(cbx_1__1__128_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__128_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__128_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__128_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__128_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__128_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__128_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__128_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__128_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__128_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__128_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__128_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__128_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__128_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__128_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__128_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[128]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[128]),
    .right_width_0_height_0__pin_16_(cby_12__1__7_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__7_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__7_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__7_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__7_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__7_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__7_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__7_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__7_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__7_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__7_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__7_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__7_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__7_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__7_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__7_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__127_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_139_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_139_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_139_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_139_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_139_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_139_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_139_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_139_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_139_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_139_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_139_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_139_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_139_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_139_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_139_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_139_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_139_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_139_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_139_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_139_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_139_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_139_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_139_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_139_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_139_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_139_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_139_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_139_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_139_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_139_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_139_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_139_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[127]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[127]),
    .ccff_tail(grid_clb_139_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__9_
  (
    .clk_0_N_in(clk_1_wires[244]),
    .prog_clk_0_N_in(prog_clk_1_wires[244]),
    .prog_clk_0_E_out(prog_clk_0_wires[468]),
    .prog_clk_0_S_out(prog_clk_0_wires[467]),
    .Reset_W_in(ResetWires[221]),
    .pReset_N_in(pResetWires[500]),
    .Test_en_W_in(Test_enWires[221]),
    .SC_OUT_TOP(scff_Wires[310]),
    .SC_IN_BOT(scff_Wires[309]),
    .top_width_0_height_0__pin_0_(cbx_1__1__129_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__129_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__129_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__129_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__129_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__129_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__129_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__129_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__129_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__129_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__129_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__129_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__129_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__129_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__129_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__129_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[129]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[129]),
    .right_width_0_height_0__pin_16_(cby_12__1__8_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__8_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__8_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__8_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__8_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__8_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__8_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__8_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__8_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__8_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__8_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__8_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__8_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__8_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__8_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__8_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__128_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_140_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_140_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_140_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_140_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_140_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_140_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_140_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_140_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_140_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_140_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_140_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_140_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_140_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_140_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_140_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_140_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_140_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_140_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_140_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_140_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_140_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_140_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_140_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_140_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_140_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_140_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_140_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_140_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_140_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_140_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_140_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_140_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[128]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[128]),
    .ccff_tail(grid_clb_140_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__10_
  (
    .clk_0_S_in(clk_1_wires[243]),
    .prog_clk_0_S_in(prog_clk_1_wires[243]),
    .prog_clk_0_E_out(prog_clk_0_wires[471]),
    .prog_clk_0_S_out(prog_clk_0_wires[470]),
    .Reset_W_in(ResetWires[243]),
    .pReset_N_in(pResetWires[549]),
    .Test_en_W_in(Test_enWires[243]),
    .SC_OUT_TOP(scff_Wires[312]),
    .SC_IN_BOT(scff_Wires[311]),
    .top_width_0_height_0__pin_0_(cbx_1__1__130_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__130_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__130_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__130_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__130_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__130_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__130_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__130_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__130_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__130_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__130_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__130_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__130_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__130_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__130_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__130_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[130]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[130]),
    .right_width_0_height_0__pin_16_(cby_12__1__9_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__9_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__9_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__9_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__9_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__9_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__9_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__9_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__9_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__9_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__9_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__9_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__9_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__9_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__9_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__9_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__129_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_141_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_141_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_141_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_141_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_141_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_141_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_141_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_141_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_141_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_141_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_141_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_141_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_141_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_141_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_141_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_141_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_141_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_141_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_141_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_141_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_141_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_141_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_141_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_141_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_141_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_141_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_141_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_141_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_141_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_141_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_141_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_141_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[129]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[129]),
    .ccff_tail(grid_clb_141_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__11_
  (
    .clk_0_N_in(clk_1_wires[251]),
    .prog_clk_0_N_in(prog_clk_1_wires[251]),
    .prog_clk_0_E_out(prog_clk_0_wires[474]),
    .prog_clk_0_S_out(prog_clk_0_wires[473]),
    .Reset_W_in(ResetWires[265]),
    .pReset_N_in(pResetWires[598]),
    .Test_en_W_in(Test_enWires[265]),
    .SC_OUT_TOP(scff_Wires[314]),
    .SC_IN_BOT(scff_Wires[313]),
    .top_width_0_height_0__pin_0_(cbx_1__1__131_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__131_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__131_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__131_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__131_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__131_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__131_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__131_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__131_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__131_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__131_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__131_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__131_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__131_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__131_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__131_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[131]),
    .top_width_0_height_0__pin_34_(cout_feedthrough_wires[131]),
    .right_width_0_height_0__pin_16_(cby_12__1__10_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__10_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__10_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__10_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__10_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__10_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__10_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__10_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__10_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__10_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__10_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__10_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__10_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__10_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__10_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__10_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__130_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_142_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_142_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_142_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_142_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_142_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_142_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_142_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_142_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_142_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_142_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_142_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_142_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_142_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_142_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_142_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_142_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_142_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_142_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_142_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_142_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_142_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_142_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_142_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_142_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_142_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_142_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_142_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_142_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_142_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_142_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_142_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_142_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[130]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[130]),
    .ccff_tail(grid_clb_142_ccff_tail[0])
  );


  grid_clb
  grid_clb_12__12_
  (
    .clk_0_S_in(clk_1_wires[250]),
    .prog_clk_0_S_in(prog_clk_1_wires[250]),
    .prog_clk_0_N_out(prog_clk_0_wires[479]),
    .prog_clk_0_E_out(prog_clk_0_wires[477]),
    .prog_clk_0_S_out(prog_clk_0_wires[476]),
    .Reset_W_in(ResetWires[287]),
    .pReset_N_in(pResetWires[636]),
    .Test_en_W_in(Test_enWires[287]),
    .SC_OUT_TOP(scff_Wires[316]),
    .SC_IN_BOT(scff_Wires[315]),
    .top_width_0_height_0__pin_0_(cbx_1__12__11_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__12__11_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__12__11_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__12__11_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__12__11_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__12__11_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__12__11_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__12__11_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__12__11_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__12__11_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__12__11_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__12__11_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__12__11_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__12__11_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__12__11_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__12__11_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_12__12__undriven_top_width_0_height_0__pin_32_[0]),
    .top_width_0_height_0__pin_34_(grid_clb_12__12__undriven_top_width_0_height_0__pin_34_[0]),
    .right_width_0_height_0__pin_16_(cby_12__1__11_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_12__1__11_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_12__1__11_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_12__1__11_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_12__1__11_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_12__1__11_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_12__1__11_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_12__1__11_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_12__1__11_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_12__1__11_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_12__1__11_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_12__1__11_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_12__1__11_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_12__1__11_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_12__1__11_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_12__1__11_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__131_ccff_tail[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_143_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_143_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_143_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_143_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_143_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_143_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_143_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_143_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_143_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_143_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_143_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_143_top_width_0_height_0__pin_41_lower[0]),
    .top_width_0_height_0__pin_42_upper(grid_clb_143_top_width_0_height_0__pin_42_upper[0]),
    .top_width_0_height_0__pin_42_lower(grid_clb_143_top_width_0_height_0__pin_42_lower[0]),
    .top_width_0_height_0__pin_43_upper(grid_clb_143_top_width_0_height_0__pin_43_upper[0]),
    .top_width_0_height_0__pin_43_lower(grid_clb_143_top_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_143_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_143_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_143_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_143_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_143_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_143_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_143_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_143_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_143_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_143_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_143_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_143_right_width_0_height_0__pin_49_lower[0]),
    .right_width_0_height_0__pin_50_upper(grid_clb_143_right_width_0_height_0__pin_50_upper[0]),
    .right_width_0_height_0__pin_50_lower(grid_clb_143_right_width_0_height_0__pin_50_lower[0]),
    .right_width_0_height_0__pin_51_upper(grid_clb_143_right_width_0_height_0__pin_51_upper[0]),
    .right_width_0_height_0__pin_51_lower(grid_clb_143_right_width_0_height_0__pin_51_lower[0]),
    .bottom_width_0_height_0__pin_52_(regin_feedthrough_wires[131]),
    .bottom_width_0_height_0__pin_54_(cin_feedthrough_wires[131]),
    .ccff_tail(grid_clb_143_ccff_tail[0])
  );


  sb_0__0_
  sb_0__0_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[5]),
    .pReset_E_in(pResetWires[25]),
    .chany_top_in(cby_0__1__0_chany_bottom_out[0:29]),
    .top_left_grid_pin_1_(grid_io_left_0_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__0__0_chanx_left_out[0:29]),
    .right_bottom_grid_pin_1_(grid_io_bottom_11_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_11_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_11_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_11_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_11_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_11_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_11_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_11_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_11_top_width_0_height_0__pin_17_upper[0]),
    .ccff_head(grid_io_bottom_11_ccff_tail[0]),
    .chany_top_out(sb_0__0__0_chany_top_out[0:29]),
    .chanx_right_out(sb_0__0__0_chanx_right_out[0:29]),
    .ccff_tail(ccff_tail[0])
  );


  sb_0__1_
  sb_0__1_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[4]),
    .pReset_S_out(pResetWires[64]),
    .pReset_E_in(pResetWires[61]),
    .chany_top_in(cby_0__1__1_chany_bottom_out[0:29]),
    .top_left_grid_pin_1_(grid_io_left_1_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__0_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_0_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_0_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_0_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_0_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_0_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_0_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_0_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_0_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_0__1__0_chany_top_out[0:29]),
    .bottom_left_grid_pin_1_(grid_io_left_0_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__0_ccff_tail[0]),
    .chany_top_out(sb_0__1__0_chany_top_out[0:29]),
    .chanx_right_out(sb_0__1__0_chanx_right_out[0:29]),
    .chany_bottom_out(sb_0__1__0_chany_bottom_out[0:29]),
    .ccff_tail(sb_0__1__0_ccff_tail[0])
  );


  sb_0__1_
  sb_0__2_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[10]),
    .pReset_S_out(pResetWires[113]),
    .pReset_E_in(pResetWires[110]),
    .chany_top_in(cby_0__1__2_chany_bottom_out[0:29]),
    .top_left_grid_pin_1_(grid_io_left_2_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__1_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_1_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_1_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_1_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_1_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_1_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_1_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_1_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_1_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_0__1__1_chany_top_out[0:29]),
    .bottom_left_grid_pin_1_(grid_io_left_1_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__1_ccff_tail[0]),
    .chany_top_out(sb_0__1__1_chany_top_out[0:29]),
    .chanx_right_out(sb_0__1__1_chanx_right_out[0:29]),
    .chany_bottom_out(sb_0__1__1_chany_bottom_out[0:29]),
    .ccff_tail(sb_0__1__1_ccff_tail[0])
  );


  sb_0__1_
  sb_0__3_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[15]),
    .pReset_S_out(pResetWires[162]),
    .pReset_E_in(pResetWires[159]),
    .chany_top_in(cby_0__1__3_chany_bottom_out[0:29]),
    .top_left_grid_pin_1_(grid_io_left_3_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__2_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_2_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_2_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_2_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_2_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_2_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_2_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_2_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_2_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_0__1__2_chany_top_out[0:29]),
    .bottom_left_grid_pin_1_(grid_io_left_2_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__2_ccff_tail[0]),
    .chany_top_out(sb_0__1__2_chany_top_out[0:29]),
    .chanx_right_out(sb_0__1__2_chanx_right_out[0:29]),
    .chany_bottom_out(sb_0__1__2_chany_bottom_out[0:29]),
    .ccff_tail(sb_0__1__2_ccff_tail[0])
  );


  sb_0__1_
  sb_0__4_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[20]),
    .pReset_S_out(pResetWires[211]),
    .pReset_E_in(pResetWires[208]),
    .chany_top_in(cby_0__1__4_chany_bottom_out[0:29]),
    .top_left_grid_pin_1_(grid_io_left_4_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__3_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_3_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_3_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_3_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_3_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_3_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_3_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_3_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_3_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_0__1__3_chany_top_out[0:29]),
    .bottom_left_grid_pin_1_(grid_io_left_3_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__3_ccff_tail[0]),
    .chany_top_out(sb_0__1__3_chany_top_out[0:29]),
    .chanx_right_out(sb_0__1__3_chanx_right_out[0:29]),
    .chany_bottom_out(sb_0__1__3_chany_bottom_out[0:29]),
    .ccff_tail(sb_0__1__3_ccff_tail[0])
  );


  sb_0__1_
  sb_0__5_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[25]),
    .pReset_S_out(pResetWires[260]),
    .pReset_E_in(pResetWires[257]),
    .chany_top_in(cby_0__1__5_chany_bottom_out[0:29]),
    .top_left_grid_pin_1_(grid_io_left_5_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__4_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_4_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_4_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_4_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_4_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_4_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_4_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_4_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_4_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_0__1__4_chany_top_out[0:29]),
    .bottom_left_grid_pin_1_(grid_io_left_4_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__4_ccff_tail[0]),
    .chany_top_out(sb_0__1__4_chany_top_out[0:29]),
    .chanx_right_out(sb_0__1__4_chanx_right_out[0:29]),
    .chany_bottom_out(sb_0__1__4_chany_bottom_out[0:29]),
    .ccff_tail(sb_0__1__4_ccff_tail[0])
  );


  sb_0__1_
  sb_0__6_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[30]),
    .pReset_S_out(pResetWires[309]),
    .pReset_E_in(pResetWires[306]),
    .chany_top_in(cby_0__1__6_chany_bottom_out[0:29]),
    .top_left_grid_pin_1_(grid_io_left_6_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__5_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_5_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_5_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_5_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_5_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_5_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_5_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_5_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_5_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_0__1__5_chany_top_out[0:29]),
    .bottom_left_grid_pin_1_(grid_io_left_5_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__5_ccff_tail[0]),
    .chany_top_out(sb_0__1__5_chany_top_out[0:29]),
    .chanx_right_out(sb_0__1__5_chanx_right_out[0:29]),
    .chany_bottom_out(sb_0__1__5_chany_bottom_out[0:29]),
    .ccff_tail(sb_0__1__5_ccff_tail[0])
  );


  sb_0__1_
  sb_0__7_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[35]),
    .pReset_S_out(pResetWires[358]),
    .pReset_E_in(pResetWires[355]),
    .chany_top_in(cby_0__1__7_chany_bottom_out[0:29]),
    .top_left_grid_pin_1_(grid_io_left_7_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__6_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_6_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_6_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_6_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_6_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_6_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_6_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_6_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_6_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_0__1__6_chany_top_out[0:29]),
    .bottom_left_grid_pin_1_(grid_io_left_6_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__6_ccff_tail[0]),
    .chany_top_out(sb_0__1__6_chany_top_out[0:29]),
    .chanx_right_out(sb_0__1__6_chanx_right_out[0:29]),
    .chany_bottom_out(sb_0__1__6_chany_bottom_out[0:29]),
    .ccff_tail(sb_0__1__6_ccff_tail[0])
  );


  sb_0__1_
  sb_0__8_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[40]),
    .pReset_S_out(pResetWires[407]),
    .pReset_E_in(pResetWires[404]),
    .chany_top_in(cby_0__1__8_chany_bottom_out[0:29]),
    .top_left_grid_pin_1_(grid_io_left_8_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__7_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_7_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_7_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_7_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_7_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_7_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_7_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_7_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_7_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_0__1__7_chany_top_out[0:29]),
    .bottom_left_grid_pin_1_(grid_io_left_7_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__7_ccff_tail[0]),
    .chany_top_out(sb_0__1__7_chany_top_out[0:29]),
    .chanx_right_out(sb_0__1__7_chanx_right_out[0:29]),
    .chany_bottom_out(sb_0__1__7_chany_bottom_out[0:29]),
    .ccff_tail(sb_0__1__7_ccff_tail[0])
  );


  sb_0__1_
  sb_0__9_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[45]),
    .pReset_S_out(pResetWires[456]),
    .pReset_E_in(pResetWires[453]),
    .chany_top_in(cby_0__1__9_chany_bottom_out[0:29]),
    .top_left_grid_pin_1_(grid_io_left_9_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__8_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_8_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_8_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_8_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_8_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_8_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_8_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_8_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_8_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_0__1__8_chany_top_out[0:29]),
    .bottom_left_grid_pin_1_(grid_io_left_8_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__8_ccff_tail[0]),
    .chany_top_out(sb_0__1__8_chany_top_out[0:29]),
    .chanx_right_out(sb_0__1__8_chanx_right_out[0:29]),
    .chany_bottom_out(sb_0__1__8_chany_bottom_out[0:29]),
    .ccff_tail(sb_0__1__8_ccff_tail[0])
  );


  sb_0__1_
  sb_0__10_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[50]),
    .pReset_S_out(pResetWires[505]),
    .pReset_E_in(pResetWires[502]),
    .chany_top_in(cby_0__1__10_chany_bottom_out[0:29]),
    .top_left_grid_pin_1_(grid_io_left_10_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__9_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_9_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_9_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_9_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_9_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_9_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_9_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_9_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_9_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_0__1__9_chany_top_out[0:29]),
    .bottom_left_grid_pin_1_(grid_io_left_9_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__9_ccff_tail[0]),
    .chany_top_out(sb_0__1__9_chany_top_out[0:29]),
    .chanx_right_out(sb_0__1__9_chanx_right_out[0:29]),
    .chany_bottom_out(sb_0__1__9_chany_bottom_out[0:29]),
    .ccff_tail(sb_0__1__9_ccff_tail[0])
  );


  sb_0__1_
  sb_0__11_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[55]),
    .pReset_S_out(pResetWires[554]),
    .pReset_E_in(pResetWires[551]),
    .chany_top_in(cby_0__1__11_chany_bottom_out[0:29]),
    .top_left_grid_pin_1_(grid_io_left_11_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__10_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_10_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_10_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_10_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_10_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_10_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_10_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_10_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_10_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_0__1__10_chany_top_out[0:29]),
    .bottom_left_grid_pin_1_(grid_io_left_10_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__10_ccff_tail[0]),
    .chany_top_out(sb_0__1__10_chany_top_out[0:29]),
    .chanx_right_out(sb_0__1__10_chanx_right_out[0:29]),
    .chany_bottom_out(sb_0__1__10_chany_bottom_out[0:29]),
    .ccff_tail(sb_0__1__10_ccff_tail[0])
  );


  sb_0__2_
  sb_0__12_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[62]),
    .pReset_S_out(pResetWires[603]),
    .pReset_E_in(pResetWires[600]),
    .SC_OUT_BOT(scff_Wires[0]),
    .SC_IN_TOP(sc_head),
    .chanx_right_in(cbx_1__12__0_chanx_left_out[0:29]),
    .right_top_grid_pin_1_(grid_io_top_0_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_11_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_11_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_11_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_11_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_11_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_11_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_11_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_11_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_0__1__11_chany_top_out[0:29]),
    .bottom_left_grid_pin_1_(grid_io_left_11_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(grid_io_top_0_ccff_tail[0]),
    .chanx_right_out(sb_0__12__0_chanx_right_out[0:29]),
    .chany_bottom_out(sb_0__12__0_chany_bottom_out[0:29]),
    .ccff_tail(sb_0__12__0_ccff_tail[0])
  );


  sb_1__0_
  sb_1__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[2]),
    .pReset_E_in(pResetWires[28]),
    .pReset_N_out(pResetWires[27]),
    .pReset_W_out(pResetWires[26]),
    .SC_OUT_TOP(scff_Wires[27]),
    .SC_IN_TOP(scff_Wires[26]),
    .chany_top_in(cby_1__1__0_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_0_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_0_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_0_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_0_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_0_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_0_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_0_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_0_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__0__1_chanx_left_out[0:29]),
    .right_bottom_grid_pin_1_(grid_io_bottom_10_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_10_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_10_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_10_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_10_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_10_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_10_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_10_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_10_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__0_chanx_right_out[0:29]),
    .left_bottom_grid_pin_1_(grid_io_bottom_11_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_11_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_11_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_11_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_11_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_11_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_11_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_11_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_11_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_10_ccff_tail[0]),
    .chany_top_out(sb_1__0__0_chany_top_out[0:29]),
    .chanx_right_out(sb_1__0__0_chanx_right_out[0:29]),
    .chanx_left_out(sb_1__0__0_chanx_left_out[0:29]),
    .ccff_tail(sb_1__0__0_ccff_tail[0])
  );


  sb_1__0_
  sb_2__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[65]),
    .pReset_E_in(pResetWires[31]),
    .pReset_N_out(pResetWires[30]),
    .pReset_W_out(pResetWires[29]),
    .chany_top_in(cby_1__1__12_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_12_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_12_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_12_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_12_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_12_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_12_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_12_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_12_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__0__2_chanx_left_out[0:29]),
    .right_bottom_grid_pin_1_(grid_io_bottom_9_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_9_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_9_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_9_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_9_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_9_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_9_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_9_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_9_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__1_chanx_right_out[0:29]),
    .left_bottom_grid_pin_1_(grid_io_bottom_10_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_10_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_10_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_10_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_10_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_10_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_10_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_10_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_10_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_9_ccff_tail[0]),
    .chany_top_out(sb_1__0__1_chany_top_out[0:29]),
    .chanx_right_out(sb_1__0__1_chanx_right_out[0:29]),
    .chanx_left_out(sb_1__0__1_chanx_left_out[0:29]),
    .ccff_tail(sb_1__0__1_ccff_tail[0])
  );


  sb_1__0_
  sb_3__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[103]),
    .pReset_E_in(pResetWires[34]),
    .pReset_N_out(pResetWires[33]),
    .pReset_W_out(pResetWires[32]),
    .SC_OUT_TOP(scff_Wires[80]),
    .SC_IN_TOP(scff_Wires[79]),
    .chany_top_in(cby_1__1__24_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_24_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_24_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_24_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_24_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_24_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_24_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_24_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_24_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__0__3_chanx_left_out[0:29]),
    .right_bottom_grid_pin_1_(grid_io_bottom_8_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_8_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_8_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_8_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_8_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_8_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_8_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_8_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_8_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__2_chanx_right_out[0:29]),
    .left_bottom_grid_pin_1_(grid_io_bottom_9_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_9_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_9_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_9_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_9_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_9_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_9_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_9_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_9_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_8_ccff_tail[0]),
    .chany_top_out(sb_1__0__2_chany_top_out[0:29]),
    .chanx_right_out(sb_1__0__2_chanx_right_out[0:29]),
    .chanx_left_out(sb_1__0__2_chanx_left_out[0:29]),
    .ccff_tail(sb_1__0__2_ccff_tail[0])
  );


  sb_1__0_
  sb_4__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[141]),
    .pReset_E_in(pResetWires[37]),
    .pReset_N_out(pResetWires[36]),
    .pReset_W_out(pResetWires[35]),
    .chany_top_in(cby_1__1__36_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_36_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_36_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_36_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_36_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_36_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_36_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_36_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_36_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__0__4_chanx_left_out[0:29]),
    .right_bottom_grid_pin_1_(grid_io_bottom_7_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_7_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_7_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_7_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_7_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_7_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_7_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_7_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_7_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__3_chanx_right_out[0:29]),
    .left_bottom_grid_pin_1_(grid_io_bottom_8_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_8_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_8_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_8_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_8_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_8_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_8_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_8_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_8_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_7_ccff_tail[0]),
    .chany_top_out(sb_1__0__3_chany_top_out[0:29]),
    .chanx_right_out(sb_1__0__3_chanx_right_out[0:29]),
    .chanx_left_out(sb_1__0__3_chanx_left_out[0:29]),
    .ccff_tail(sb_1__0__3_ccff_tail[0])
  );


  sb_1__0_
  sb_5__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[179]),
    .pReset_E_in(pResetWires[40]),
    .pReset_N_out(pResetWires[39]),
    .pReset_W_out(pResetWires[38]),
    .SC_OUT_TOP(scff_Wires[133]),
    .SC_IN_TOP(scff_Wires[132]),
    .chany_top_in(cby_1__1__48_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_48_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_48_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_48_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_48_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_48_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_48_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_48_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_48_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__0__5_chanx_left_out[0:29]),
    .right_bottom_grid_pin_1_(grid_io_bottom_6_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_6_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_6_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_6_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_6_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_6_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_6_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_6_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_6_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__4_chanx_right_out[0:29]),
    .left_bottom_grid_pin_1_(grid_io_bottom_7_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_7_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_7_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_7_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_7_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_7_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_7_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_7_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_7_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_6_ccff_tail[0]),
    .chany_top_out(sb_1__0__4_chany_top_out[0:29]),
    .chanx_right_out(sb_1__0__4_chanx_right_out[0:29]),
    .chanx_left_out(sb_1__0__4_chanx_left_out[0:29]),
    .ccff_tail(sb_1__0__4_ccff_tail[0])
  );


  sb_1__0_
  sb_6__0_
  (
    .clk_3_N_out(clk_3_wires[90]),
    .clk_3_S_in(clk),
    .prog_clk_3_N_out(prog_clk_3_wires[90]),
    .prog_clk_3_S_in(prog_clk),
    .prog_clk_0_N_in(prog_clk_0_wires[217]),
    .Reset_N_out(ResetWires[1]),
    .Reset_S_in(Reset),
    .pReset_E_out(pResetWires[43]),
    .pReset_W_out(pResetWires[41]),
    .pReset_N_out(pResetWires[42]),
    .pReset_S_in(pReset),
    .Test_en_N_out(Test_enWires[1]),
    .Test_en_S_in(Test_en),
    .chany_top_in(cby_1__1__60_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_60_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_60_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_60_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_60_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_60_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_60_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_60_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_60_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__0__6_chanx_left_out[0:29]),
    .right_bottom_grid_pin_1_(grid_io_bottom_5_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_5_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_5_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_5_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_5_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_5_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_5_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_5_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_5_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__5_chanx_right_out[0:29]),
    .left_bottom_grid_pin_1_(grid_io_bottom_6_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_6_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_6_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_6_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_6_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_6_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_6_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_6_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_6_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_5_ccff_tail[0]),
    .chany_top_out(sb_1__0__5_chany_top_out[0:29]),
    .chanx_right_out(sb_1__0__5_chanx_right_out[0:29]),
    .chanx_left_out(sb_1__0__5_chanx_left_out[0:29]),
    .ccff_tail(sb_1__0__5_ccff_tail[0])
  );


  sb_1__0_
  sb_7__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[255]),
    .pReset_E_out(pResetWires[46]),
    .pReset_N_out(pResetWires[45]),
    .pReset_W_in(pResetWires[44]),
    .SC_OUT_TOP(scff_Wires[186]),
    .SC_IN_TOP(scff_Wires[185]),
    .chany_top_in(cby_1__1__72_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_72_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_72_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_72_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_72_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_72_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_72_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_72_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_72_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__0__7_chanx_left_out[0:29]),
    .right_bottom_grid_pin_1_(grid_io_bottom_4_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_4_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_4_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_4_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_4_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_4_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_4_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_4_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_4_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__6_chanx_right_out[0:29]),
    .left_bottom_grid_pin_1_(grid_io_bottom_5_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_5_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_5_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_5_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_5_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_5_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_5_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_5_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_5_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_4_ccff_tail[0]),
    .chany_top_out(sb_1__0__6_chany_top_out[0:29]),
    .chanx_right_out(sb_1__0__6_chanx_right_out[0:29]),
    .chanx_left_out(sb_1__0__6_chanx_left_out[0:29]),
    .ccff_tail(sb_1__0__6_ccff_tail[0])
  );


  sb_1__0_
  sb_8__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[293]),
    .pReset_E_out(pResetWires[49]),
    .pReset_N_out(pResetWires[48]),
    .pReset_W_in(pResetWires[47]),
    .chany_top_in(cby_1__1__84_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_84_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_84_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_84_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_84_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_84_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_84_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_84_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_84_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__0__8_chanx_left_out[0:29]),
    .right_bottom_grid_pin_1_(grid_io_bottom_3_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_3_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_3_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_3_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_3_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_3_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_3_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_3_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_3_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__7_chanx_right_out[0:29]),
    .left_bottom_grid_pin_1_(grid_io_bottom_4_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_4_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_4_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_4_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_4_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_4_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_4_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_4_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_4_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_3_ccff_tail[0]),
    .chany_top_out(sb_1__0__7_chany_top_out[0:29]),
    .chanx_right_out(sb_1__0__7_chanx_right_out[0:29]),
    .chanx_left_out(sb_1__0__7_chanx_left_out[0:29]),
    .ccff_tail(sb_1__0__7_ccff_tail[0])
  );


  sb_1__0_
  sb_9__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[331]),
    .pReset_E_out(pResetWires[52]),
    .pReset_N_out(pResetWires[51]),
    .pReset_W_in(pResetWires[50]),
    .SC_OUT_TOP(scff_Wires[239]),
    .SC_IN_TOP(scff_Wires[238]),
    .chany_top_in(cby_1__1__96_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_96_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_96_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_96_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_96_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_96_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_96_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_96_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_96_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__0__9_chanx_left_out[0:29]),
    .right_bottom_grid_pin_1_(grid_io_bottom_2_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_2_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_2_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_2_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_2_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_2_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_2_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_2_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_2_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__8_chanx_right_out[0:29]),
    .left_bottom_grid_pin_1_(grid_io_bottom_3_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_3_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_3_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_3_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_3_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_3_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_3_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_3_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_3_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_2_ccff_tail[0]),
    .chany_top_out(sb_1__0__8_chany_top_out[0:29]),
    .chanx_right_out(sb_1__0__8_chanx_right_out[0:29]),
    .chanx_left_out(sb_1__0__8_chanx_left_out[0:29]),
    .ccff_tail(sb_1__0__8_ccff_tail[0])
  );


  sb_1__0_
  sb_10__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[369]),
    .pReset_E_out(pResetWires[55]),
    .pReset_N_out(pResetWires[54]),
    .pReset_W_in(pResetWires[53]),
    .chany_top_in(cby_1__1__108_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_108_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_108_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_108_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_108_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_108_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_108_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_108_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_108_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__0__10_chanx_left_out[0:29]),
    .right_bottom_grid_pin_1_(grid_io_bottom_1_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_1_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_1_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_1_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_1_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_1_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_1_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_1_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_1_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__9_chanx_right_out[0:29]),
    .left_bottom_grid_pin_1_(grid_io_bottom_2_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_2_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_2_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_2_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_2_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_2_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_2_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_2_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_2_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_1_ccff_tail[0]),
    .chany_top_out(sb_1__0__9_chany_top_out[0:29]),
    .chanx_right_out(sb_1__0__9_chanx_right_out[0:29]),
    .chanx_left_out(sb_1__0__9_chanx_left_out[0:29]),
    .ccff_tail(sb_1__0__9_ccff_tail[0])
  );


  sb_1__0_
  sb_11__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[407]),
    .pReset_E_out(pResetWires[58]),
    .pReset_N_out(pResetWires[57]),
    .pReset_W_in(pResetWires[56]),
    .SC_OUT_TOP(scff_Wires[292]),
    .SC_IN_TOP(scff_Wires[291]),
    .chany_top_in(cby_1__1__120_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_120_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_120_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_120_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_120_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_120_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_120_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_120_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_120_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__0__11_chanx_left_out[0:29]),
    .right_bottom_grid_pin_1_(grid_io_bottom_0_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_0_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_0_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_0_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_0_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_0_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_0_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_0_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_0_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__10_chanx_right_out[0:29]),
    .left_bottom_grid_pin_1_(grid_io_bottom_1_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_1_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_1_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_1_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_1_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_1_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_1_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_1_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_1_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_0_ccff_tail[0]),
    .chany_top_out(sb_1__0__10_chany_top_out[0:29]),
    .chanx_right_out(sb_1__0__10_chanx_right_out[0:29]),
    .chanx_left_out(sb_1__0__10_chanx_left_out[0:29]),
    .ccff_tail(sb_1__0__10_ccff_tail[0])
  );


  sb_1__1_
  sb_1__1_
  (
    .clk_1_N_in(clk_2_wires[4]),
    .clk_1_W_out(clk_1_wires[2]),
    .clk_1_E_out(clk_1_wires[1]),
    .prog_clk_1_N_in(prog_clk_2_wires[4]),
    .prog_clk_1_W_out(prog_clk_1_wires[2]),
    .prog_clk_1_E_out(prog_clk_1_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[8]),
    .pReset_E_in(pResetWires[66]),
    .pReset_N_out(pResetWires[65]),
    .pReset_W_out(pResetWires[62]),
    .chany_top_in(cby_1__1__1_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_1_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_1_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_1_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_1_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_1_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_1_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_1_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_1_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__11_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_12_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_12_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_12_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_12_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_12_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_12_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_12_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_12_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__0_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_0_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_0_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_0_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_0_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_0_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_0_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_0_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_0_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__0_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_0_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_0_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_0_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_0_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_0_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_0_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_0_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_0_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__11_ccff_tail[0]),
    .chany_top_out(sb_1__1__0_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__0_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__0_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__0_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__0_ccff_tail[0])
  );


  sb_1__1_
  sb_1__2_
  (
    .clk_2_S_out(clk_2_wires[3]),
    .clk_2_E_in(clk_2_wires[1]),
    .prog_clk_2_S_out(prog_clk_2_wires[3]),
    .prog_clk_2_E_in(prog_clk_2_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[13]),
    .pReset_E_in(pResetWires[115]),
    .pReset_N_out(pResetWires[114]),
    .pReset_W_out(pResetWires[111]),
    .chany_top_in(cby_1__1__2_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_2_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_2_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_2_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_2_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_2_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_2_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_2_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_2_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__12_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_13_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_13_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_13_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_13_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_13_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_13_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_13_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_13_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__1_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_1_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_1_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_1_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_1_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_1_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_1_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_1_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_1_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__1_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_1_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_1_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_1_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_1_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_1_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_1_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_1_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_1_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__12_ccff_tail[0]),
    .chany_top_out(sb_1__1__1_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__1_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__1_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__1_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__1_ccff_tail[0])
  );


  sb_1__1_
  sb_1__3_
  (
    .clk_1_N_in(clk_2_wires[11]),
    .clk_1_W_out(clk_1_wires[9]),
    .clk_1_E_out(clk_1_wires[8]),
    .prog_clk_1_N_in(prog_clk_2_wires[11]),
    .prog_clk_1_W_out(prog_clk_1_wires[9]),
    .prog_clk_1_E_out(prog_clk_1_wires[8]),
    .prog_clk_0_N_in(prog_clk_0_wires[18]),
    .pReset_E_in(pResetWires[164]),
    .pReset_N_out(pResetWires[163]),
    .pReset_W_out(pResetWires[160]),
    .chany_top_in(cby_1__1__3_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_3_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_3_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_3_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_3_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_3_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_3_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_3_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_3_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__13_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_14_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_14_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_14_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_14_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_14_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_14_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_14_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_14_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__2_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_2_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_2_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_2_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_2_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_2_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_2_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_2_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_2_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__2_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_2_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_2_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_2_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_2_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_2_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_2_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_2_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_2_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__13_ccff_tail[0]),
    .chany_top_out(sb_1__1__2_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__2_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__2_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__2_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__2_ccff_tail[0])
  );


  sb_1__1_
  sb_1__4_
  (
    .clk_2_S_out(clk_2_wires[10]),
    .clk_2_N_out(clk_2_wires[8]),
    .clk_2_E_in(clk_2_wires[6]),
    .prog_clk_2_S_out(prog_clk_2_wires[10]),
    .prog_clk_2_N_out(prog_clk_2_wires[8]),
    .prog_clk_2_E_in(prog_clk_2_wires[6]),
    .prog_clk_0_N_in(prog_clk_0_wires[23]),
    .pReset_E_in(pResetWires[213]),
    .pReset_N_out(pResetWires[212]),
    .pReset_W_out(pResetWires[209]),
    .chany_top_in(cby_1__1__4_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_4_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_4_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_4_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_4_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_4_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_4_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_4_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_4_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__14_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_15_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_15_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_15_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_15_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_15_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_15_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_15_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_15_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__3_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_3_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_3_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_3_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_3_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_3_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_3_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_3_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_3_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__3_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_3_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_3_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_3_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_3_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_3_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_3_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_3_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_3_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__14_ccff_tail[0]),
    .chany_top_out(sb_1__1__3_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__3_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__3_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__3_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__3_ccff_tail[0])
  );


  sb_1__1_
  sb_1__5_
  (
    .clk_1_S_in(clk_2_wires[9]),
    .clk_1_W_out(clk_1_wires[16]),
    .clk_1_E_out(clk_1_wires[15]),
    .prog_clk_1_S_in(prog_clk_2_wires[9]),
    .prog_clk_1_W_out(prog_clk_1_wires[16]),
    .prog_clk_1_E_out(prog_clk_1_wires[15]),
    .prog_clk_0_N_in(prog_clk_0_wires[28]),
    .pReset_E_in(pResetWires[262]),
    .pReset_N_out(pResetWires[261]),
    .pReset_W_out(pResetWires[258]),
    .chany_top_in(cby_1__1__5_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_5_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_5_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_5_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_5_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_5_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_5_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_5_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_5_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__15_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_16_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_16_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_16_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_16_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_16_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_16_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_16_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_16_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__4_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_4_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_4_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_4_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_4_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_4_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_4_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_4_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_4_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__4_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_4_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_4_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_4_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_4_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_4_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_4_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_4_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_4_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__15_ccff_tail[0]),
    .chany_top_out(sb_1__1__4_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__4_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__4_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__4_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__4_ccff_tail[0])
  );


  sb_1__1_
  sb_1__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[33]),
    .pReset_E_in(pResetWires[311]),
    .pReset_N_out(pResetWires[310]),
    .pReset_W_out(pResetWires[307]),
    .chany_top_in(cby_1__1__6_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_6_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_6_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_6_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_6_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_6_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_6_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_6_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_6_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__16_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_17_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_17_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_17_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_17_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_17_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_17_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_17_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_17_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__5_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_5_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_5_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_5_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_5_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_5_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_5_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_5_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_5_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__5_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_5_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_5_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_5_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_5_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_5_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_5_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_5_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_5_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__16_ccff_tail[0]),
    .chany_top_out(sb_1__1__5_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__5_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__5_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__5_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__5_ccff_tail[0])
  );


  sb_1__1_
  sb_1__7_
  (
    .clk_1_N_in(clk_2_wires[18]),
    .clk_1_W_out(clk_1_wires[23]),
    .clk_1_E_out(clk_1_wires[22]),
    .prog_clk_1_N_in(prog_clk_2_wires[18]),
    .prog_clk_1_W_out(prog_clk_1_wires[23]),
    .prog_clk_1_E_out(prog_clk_1_wires[22]),
    .prog_clk_0_N_in(prog_clk_0_wires[38]),
    .pReset_E_in(pResetWires[360]),
    .pReset_N_out(pResetWires[359]),
    .pReset_W_out(pResetWires[356]),
    .chany_top_in(cby_1__1__7_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_7_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_7_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_7_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_7_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_7_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_7_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_7_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_7_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__17_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_18_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_18_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_18_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_18_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_18_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_18_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_18_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_18_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__6_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_6_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_6_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_6_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_6_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_6_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_6_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_6_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_6_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__6_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_6_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_6_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_6_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_6_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_6_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_6_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_6_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_6_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__17_ccff_tail[0]),
    .chany_top_out(sb_1__1__6_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__6_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__6_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__6_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__6_ccff_tail[0])
  );


  sb_1__1_
  sb_1__8_
  (
    .clk_2_S_out(clk_2_wires[17]),
    .clk_2_N_out(clk_2_wires[15]),
    .clk_2_E_in(clk_2_wires[13]),
    .prog_clk_2_S_out(prog_clk_2_wires[17]),
    .prog_clk_2_N_out(prog_clk_2_wires[15]),
    .prog_clk_2_E_in(prog_clk_2_wires[13]),
    .prog_clk_0_N_in(prog_clk_0_wires[43]),
    .pReset_E_in(pResetWires[409]),
    .pReset_N_out(pResetWires[408]),
    .pReset_W_out(pResetWires[405]),
    .chany_top_in(cby_1__1__8_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_8_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_8_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_8_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_8_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_8_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_8_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_8_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_8_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__18_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_19_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_19_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_19_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_19_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_19_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_19_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_19_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_19_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__7_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_7_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_7_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_7_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_7_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_7_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_7_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_7_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_7_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__7_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_7_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_7_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_7_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_7_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_7_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_7_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_7_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_7_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__18_ccff_tail[0]),
    .chany_top_out(sb_1__1__7_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__7_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__7_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__7_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__7_ccff_tail[0])
  );


  sb_1__1_
  sb_1__9_
  (
    .clk_1_S_in(clk_2_wires[16]),
    .clk_1_W_out(clk_1_wires[30]),
    .clk_1_E_out(clk_1_wires[29]),
    .prog_clk_1_S_in(prog_clk_2_wires[16]),
    .prog_clk_1_W_out(prog_clk_1_wires[30]),
    .prog_clk_1_E_out(prog_clk_1_wires[29]),
    .prog_clk_0_N_in(prog_clk_0_wires[48]),
    .pReset_E_in(pResetWires[458]),
    .pReset_N_out(pResetWires[457]),
    .pReset_W_out(pResetWires[454]),
    .chany_top_in(cby_1__1__9_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_9_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_9_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_9_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_9_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_9_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_9_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_9_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_9_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__19_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_20_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_20_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_20_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_20_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_20_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_20_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_20_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_20_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__8_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_8_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_8_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_8_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_8_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_8_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_8_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_8_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_8_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__8_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_8_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_8_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_8_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_8_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_8_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_8_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_8_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_8_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__19_ccff_tail[0]),
    .chany_top_out(sb_1__1__8_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__8_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__8_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__8_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__8_ccff_tail[0])
  );


  sb_1__1_
  sb_1__10_
  (
    .clk_2_N_out(clk_2_wires[22]),
    .clk_2_E_in(clk_2_wires[20]),
    .prog_clk_2_N_out(prog_clk_2_wires[22]),
    .prog_clk_2_E_in(prog_clk_2_wires[20]),
    .prog_clk_0_N_in(prog_clk_0_wires[53]),
    .pReset_E_in(pResetWires[507]),
    .pReset_N_out(pResetWires[506]),
    .pReset_W_out(pResetWires[503]),
    .chany_top_in(cby_1__1__10_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_10_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_10_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_10_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_10_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_10_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_10_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_10_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_10_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__20_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_21_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_21_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_21_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_21_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_21_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_21_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_21_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_21_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__9_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_9_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_9_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_9_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_9_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_9_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_9_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_9_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_9_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__9_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_9_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_9_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_9_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_9_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_9_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_9_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_9_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_9_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__20_ccff_tail[0]),
    .chany_top_out(sb_1__1__9_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__9_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__9_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__9_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__9_ccff_tail[0])
  );


  sb_1__1_
  sb_1__11_
  (
    .clk_1_S_in(clk_2_wires[23]),
    .clk_1_W_out(clk_1_wires[37]),
    .clk_1_E_out(clk_1_wires[36]),
    .prog_clk_1_S_in(prog_clk_2_wires[23]),
    .prog_clk_1_W_out(prog_clk_1_wires[37]),
    .prog_clk_1_E_out(prog_clk_1_wires[36]),
    .prog_clk_0_N_in(prog_clk_0_wires[58]),
    .pReset_E_in(pResetWires[556]),
    .pReset_N_out(pResetWires[555]),
    .pReset_W_out(pResetWires[552]),
    .chany_top_in(cby_1__1__11_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_11_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_11_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_11_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_11_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_11_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_11_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_11_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_11_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__21_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_22_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_22_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_22_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_22_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_22_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_22_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_22_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_22_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__10_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_10_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_10_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_10_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_10_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_10_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_10_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_10_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_10_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__10_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_10_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_10_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_10_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_10_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_10_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_10_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_10_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_10_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__21_ccff_tail[0]),
    .chany_top_out(sb_1__1__10_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__10_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__10_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__10_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__10_ccff_tail[0])
  );


  sb_1__1_
  sb_2__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[68]),
    .pReset_E_in(pResetWires[70]),
    .pReset_N_out(pResetWires[69]),
    .pReset_W_out(pResetWires[67]),
    .chany_top_in(cby_1__1__13_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_13_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_13_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_13_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_13_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_13_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_13_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_13_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_13_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__22_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_24_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_24_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_24_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_24_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_24_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_24_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_24_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_24_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__12_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_12_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_12_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_12_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_12_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_12_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_12_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_12_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_12_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__11_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_12_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_12_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_12_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_12_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_12_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_12_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_12_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_12_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__22_ccff_tail[0]),
    .chany_top_out(sb_1__1__11_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__11_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__11_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__11_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__11_ccff_tail[0])
  );


  sb_1__1_
  sb_2__2_
  (
    .clk_2_N_in(clk_3_wires[69]),
    .clk_2_W_out(clk_2_wires[2]),
    .prog_clk_2_N_in(prog_clk_3_wires[69]),
    .prog_clk_2_W_out(prog_clk_2_wires[2]),
    .prog_clk_0_N_in(prog_clk_0_wires[71]),
    .pReset_E_in(pResetWires[119]),
    .pReset_N_out(pResetWires[118]),
    .pReset_W_out(pResetWires[116]),
    .chany_top_in(cby_1__1__14_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_14_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_14_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_14_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_14_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_14_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_14_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_14_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_14_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__23_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_25_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_25_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_25_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_25_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_25_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_25_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_25_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_25_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__13_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_13_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_13_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_13_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_13_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_13_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_13_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_13_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_13_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__12_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_13_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_13_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_13_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_13_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_13_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_13_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_13_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_13_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__23_ccff_tail[0]),
    .chany_top_out(sb_1__1__12_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__12_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__12_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__12_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__12_ccff_tail[0])
  );


  sb_1__1_
  sb_2__3_
  (
    .clk_3_S_out(clk_3_wires[68]),
    .clk_3_N_in(clk_3_wires[65]),
    .prog_clk_3_S_out(prog_clk_3_wires[68]),
    .prog_clk_3_N_in(prog_clk_3_wires[65]),
    .prog_clk_0_N_in(prog_clk_0_wires[74]),
    .pReset_E_in(pResetWires[168]),
    .pReset_N_out(pResetWires[167]),
    .pReset_W_out(pResetWires[165]),
    .chany_top_in(cby_1__1__15_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_15_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_15_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_15_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_15_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_15_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_15_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_15_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_15_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__24_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_26_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_26_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_26_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_26_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_26_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_26_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_26_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_26_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__14_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_14_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_14_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_14_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_14_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_14_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_14_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_14_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_14_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__13_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_14_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_14_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_14_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_14_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_14_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_14_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_14_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_14_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__24_ccff_tail[0]),
    .chany_top_out(sb_1__1__13_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__13_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__13_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__13_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__13_ccff_tail[0])
  );


  sb_1__1_
  sb_2__4_
  (
    .clk_3_S_out(clk_3_wires[64]),
    .clk_2_N_in(clk_3_wires[59]),
    .clk_3_N_in(clk_3_wires[59]),
    .clk_2_W_out(clk_2_wires[7]),
    .prog_clk_3_S_out(prog_clk_3_wires[64]),
    .prog_clk_2_N_in(prog_clk_3_wires[59]),
    .prog_clk_3_N_in(prog_clk_3_wires[59]),
    .prog_clk_2_W_out(prog_clk_2_wires[7]),
    .prog_clk_0_N_in(prog_clk_0_wires[77]),
    .pReset_E_in(pResetWires[217]),
    .pReset_N_out(pResetWires[216]),
    .pReset_W_out(pResetWires[214]),
    .chany_top_in(cby_1__1__16_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_16_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_16_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_16_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_16_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_16_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_16_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_16_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_16_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__25_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_27_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_27_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_27_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_27_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_27_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_27_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_27_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_27_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__15_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_15_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_15_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_15_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_15_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_15_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_15_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_15_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_15_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__14_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_15_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_15_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_15_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_15_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_15_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_15_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_15_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_15_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__25_ccff_tail[0]),
    .chany_top_out(sb_1__1__14_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__14_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__14_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__14_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__14_ccff_tail[0])
  );


  sb_1__1_
  sb_2__5_
  (
    .clk_3_S_out(clk_3_wires[58]),
    .clk_3_N_in(clk_3_wires[55]),
    .prog_clk_3_S_out(prog_clk_3_wires[58]),
    .prog_clk_3_N_in(prog_clk_3_wires[55]),
    .prog_clk_0_N_in(prog_clk_0_wires[80]),
    .pReset_E_in(pResetWires[266]),
    .pReset_N_out(pResetWires[265]),
    .pReset_W_out(pResetWires[263]),
    .chany_top_in(cby_1__1__17_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_17_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_17_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_17_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_17_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_17_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_17_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_17_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_17_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__26_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_28_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_28_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_28_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_28_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_28_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_28_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_28_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_28_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__16_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_16_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_16_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_16_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_16_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_16_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_16_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_16_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_16_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__15_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_16_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_16_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_16_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_16_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_16_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_16_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_16_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_16_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__26_ccff_tail[0]),
    .chany_top_out(sb_1__1__15_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__15_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__15_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__15_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__15_ccff_tail[0])
  );


  sb_1__1_
  sb_2__6_
  (
    .clk_3_S_out(clk_3_wires[54]),
    .clk_3_N_out(clk_3_wires[52]),
    .clk_3_E_in(clk_3_wires[51]),
    .prog_clk_3_S_out(prog_clk_3_wires[54]),
    .prog_clk_3_N_out(prog_clk_3_wires[52]),
    .prog_clk_3_E_in(prog_clk_3_wires[51]),
    .prog_clk_0_N_in(prog_clk_0_wires[83]),
    .pReset_E_in(pResetWires[315]),
    .pReset_N_out(pResetWires[314]),
    .pReset_W_out(pResetWires[312]),
    .chany_top_in(cby_1__1__18_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_18_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_18_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_18_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_18_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_18_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_18_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_18_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_18_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__27_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_29_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_29_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_29_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_29_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_29_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_29_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_29_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_29_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__17_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_17_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_17_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_17_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_17_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_17_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_17_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_17_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_17_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__16_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_17_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_17_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_17_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_17_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_17_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_17_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_17_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_17_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__27_ccff_tail[0]),
    .chany_top_out(sb_1__1__16_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__16_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__16_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__16_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__16_ccff_tail[0])
  );


  sb_1__1_
  sb_2__7_
  (
    .clk_3_N_out(clk_3_wires[56]),
    .clk_3_S_in(clk_3_wires[53]),
    .prog_clk_3_N_out(prog_clk_3_wires[56]),
    .prog_clk_3_S_in(prog_clk_3_wires[53]),
    .prog_clk_0_N_in(prog_clk_0_wires[86]),
    .pReset_E_in(pResetWires[364]),
    .pReset_N_out(pResetWires[363]),
    .pReset_W_out(pResetWires[361]),
    .chany_top_in(cby_1__1__19_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_19_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_19_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_19_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_19_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_19_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_19_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_19_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_19_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__28_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_30_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_30_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_30_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_30_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_30_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_30_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_30_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_30_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__18_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_18_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_18_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_18_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_18_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_18_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_18_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_18_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_18_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__17_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_18_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_18_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_18_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_18_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_18_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_18_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_18_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_18_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__28_ccff_tail[0]),
    .chany_top_out(sb_1__1__17_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__17_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__17_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__17_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__17_ccff_tail[0])
  );


  sb_1__1_
  sb_2__8_
  (
    .clk_3_N_out(clk_3_wires[62]),
    .clk_2_S_in(clk_3_wires[57]),
    .clk_3_S_in(clk_3_wires[57]),
    .clk_2_W_out(clk_2_wires[14]),
    .prog_clk_3_N_out(prog_clk_3_wires[62]),
    .prog_clk_2_S_in(prog_clk_3_wires[57]),
    .prog_clk_3_S_in(prog_clk_3_wires[57]),
    .prog_clk_2_W_out(prog_clk_2_wires[14]),
    .prog_clk_0_N_in(prog_clk_0_wires[89]),
    .pReset_E_in(pResetWires[413]),
    .pReset_N_out(pResetWires[412]),
    .pReset_W_out(pResetWires[410]),
    .chany_top_in(cby_1__1__20_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_20_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_20_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_20_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_20_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_20_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_20_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_20_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_20_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__29_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_31_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_31_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_31_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_31_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_31_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_31_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_31_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_31_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__19_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_19_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_19_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_19_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_19_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_19_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_19_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_19_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_19_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__18_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_19_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_19_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_19_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_19_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_19_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_19_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_19_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_19_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__29_ccff_tail[0]),
    .chany_top_out(sb_1__1__18_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__18_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__18_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__18_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__18_ccff_tail[0])
  );


  sb_1__1_
  sb_2__9_
  (
    .clk_3_N_out(clk_3_wires[66]),
    .clk_3_S_in(clk_3_wires[63]),
    .prog_clk_3_N_out(prog_clk_3_wires[66]),
    .prog_clk_3_S_in(prog_clk_3_wires[63]),
    .prog_clk_0_N_in(prog_clk_0_wires[92]),
    .pReset_E_in(pResetWires[462]),
    .pReset_N_out(pResetWires[461]),
    .pReset_W_out(pResetWires[459]),
    .chany_top_in(cby_1__1__21_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_21_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_21_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_21_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_21_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_21_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_21_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_21_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_21_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__30_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_32_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_32_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_32_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_32_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_32_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_32_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_32_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_32_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__20_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_20_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_20_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_20_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_20_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_20_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_20_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_20_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_20_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__19_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_20_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_20_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_20_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_20_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_20_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_20_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_20_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_20_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__30_ccff_tail[0]),
    .chany_top_out(sb_1__1__19_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__19_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__19_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__19_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__19_ccff_tail[0])
  );


  sb_1__1_
  sb_2__10_
  (
    .clk_2_S_in(clk_3_wires[67]),
    .clk_2_W_out(clk_2_wires[21]),
    .prog_clk_2_S_in(prog_clk_3_wires[67]),
    .prog_clk_2_W_out(prog_clk_2_wires[21]),
    .prog_clk_0_N_in(prog_clk_0_wires[95]),
    .pReset_E_in(pResetWires[511]),
    .pReset_N_out(pResetWires[510]),
    .pReset_W_out(pResetWires[508]),
    .chany_top_in(cby_1__1__22_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_22_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_22_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_22_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_22_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_22_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_22_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_22_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_22_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__31_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_33_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_33_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_33_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_33_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_33_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_33_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_33_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_33_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__21_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_21_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_21_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_21_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_21_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_21_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_21_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_21_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_21_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__20_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_21_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_21_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_21_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_21_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_21_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_21_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_21_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_21_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__31_ccff_tail[0]),
    .chany_top_out(sb_1__1__20_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__20_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__20_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__20_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__20_ccff_tail[0])
  );


  sb_1__1_
  sb_2__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[98]),
    .pReset_E_in(pResetWires[560]),
    .pReset_N_out(pResetWires[559]),
    .pReset_W_out(pResetWires[557]),
    .chany_top_in(cby_1__1__23_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_23_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_23_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_23_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_23_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_23_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_23_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_23_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_23_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__32_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_34_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_34_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_34_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_34_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_34_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_34_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_34_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_34_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__22_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_22_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_22_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_22_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_22_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_22_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_22_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_22_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_22_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__21_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_22_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_22_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_22_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_22_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_22_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_22_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_22_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_22_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__32_ccff_tail[0]),
    .chany_top_out(sb_1__1__21_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__21_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__21_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__21_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__21_ccff_tail[0])
  );


  sb_1__1_
  sb_3__1_
  (
    .clk_1_N_in(clk_2_wires[30]),
    .clk_1_W_out(clk_1_wires[44]),
    .clk_1_E_out(clk_1_wires[43]),
    .prog_clk_1_N_in(prog_clk_2_wires[30]),
    .prog_clk_1_W_out(prog_clk_1_wires[44]),
    .prog_clk_1_E_out(prog_clk_1_wires[43]),
    .prog_clk_0_N_in(prog_clk_0_wires[106]),
    .pReset_E_in(pResetWires[74]),
    .pReset_N_out(pResetWires[73]),
    .pReset_W_out(pResetWires[71]),
    .chany_top_in(cby_1__1__25_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_25_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_25_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_25_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_25_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_25_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_25_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_25_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_25_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__33_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_36_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_36_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_36_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_36_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_36_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_36_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_36_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_36_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__24_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_24_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_24_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_24_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_24_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_24_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_24_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_24_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_24_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__22_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_24_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_24_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_24_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_24_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_24_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_24_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_24_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_24_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__33_ccff_tail[0]),
    .chany_top_out(sb_1__1__22_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__22_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__22_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__22_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__22_ccff_tail[0])
  );


  sb_1__1_
  sb_3__2_
  (
    .clk_2_S_out(clk_2_wires[29]),
    .clk_2_E_in(clk_2_wires[28]),
    .prog_clk_2_S_out(prog_clk_2_wires[29]),
    .prog_clk_2_E_in(prog_clk_2_wires[28]),
    .prog_clk_0_N_in(prog_clk_0_wires[109]),
    .pReset_E_in(pResetWires[123]),
    .pReset_N_out(pResetWires[122]),
    .pReset_W_out(pResetWires[120]),
    .chany_top_in(cby_1__1__26_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_26_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_26_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_26_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_26_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_26_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_26_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_26_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_26_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__34_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_37_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_37_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_37_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_37_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_37_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_37_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_37_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_37_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__25_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_25_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_25_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_25_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_25_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_25_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_25_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_25_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_25_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__23_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_25_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_25_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_25_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_25_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_25_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_25_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_25_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_25_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__34_ccff_tail[0]),
    .chany_top_out(sb_1__1__23_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__23_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__23_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__23_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__23_ccff_tail[0])
  );


  sb_1__1_
  sb_3__3_
  (
    .clk_1_N_in(clk_2_wires[41]),
    .clk_1_W_out(clk_1_wires[51]),
    .clk_1_E_out(clk_1_wires[50]),
    .prog_clk_1_N_in(prog_clk_2_wires[41]),
    .prog_clk_1_W_out(prog_clk_1_wires[51]),
    .prog_clk_1_E_out(prog_clk_1_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[112]),
    .pReset_E_in(pResetWires[172]),
    .pReset_N_out(pResetWires[171]),
    .pReset_W_out(pResetWires[169]),
    .chany_top_in(cby_1__1__27_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_27_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_27_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_27_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_27_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_27_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_27_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_27_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_27_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__35_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_38_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_38_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_38_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_38_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_38_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_38_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_38_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_38_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__26_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_26_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_26_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_26_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_26_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_26_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_26_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_26_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_26_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__24_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_26_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_26_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_26_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_26_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_26_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_26_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_26_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_26_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__35_ccff_tail[0]),
    .chany_top_out(sb_1__1__24_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__24_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__24_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__24_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__24_ccff_tail[0])
  );


  sb_1__1_
  sb_3__4_
  (
    .clk_2_S_out(clk_2_wires[40]),
    .clk_2_N_out(clk_2_wires[38]),
    .clk_2_E_in(clk_2_wires[37]),
    .prog_clk_2_S_out(prog_clk_2_wires[40]),
    .prog_clk_2_N_out(prog_clk_2_wires[38]),
    .prog_clk_2_E_in(prog_clk_2_wires[37]),
    .prog_clk_0_N_in(prog_clk_0_wires[115]),
    .pReset_E_in(pResetWires[221]),
    .pReset_N_out(pResetWires[220]),
    .pReset_W_out(pResetWires[218]),
    .chany_top_in(cby_1__1__28_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_28_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_28_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_28_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_28_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_28_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_28_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_28_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_28_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__36_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_39_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_39_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_39_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_39_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_39_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_39_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_39_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_39_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__27_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_27_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_27_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_27_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_27_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_27_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_27_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_27_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_27_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__25_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_27_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_27_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_27_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_27_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_27_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_27_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_27_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_27_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__36_ccff_tail[0]),
    .chany_top_out(sb_1__1__25_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__25_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__25_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__25_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__25_ccff_tail[0])
  );


  sb_1__1_
  sb_3__5_
  (
    .clk_1_S_in(clk_2_wires[39]),
    .clk_1_W_out(clk_1_wires[58]),
    .clk_1_E_out(clk_1_wires[57]),
    .prog_clk_1_S_in(prog_clk_2_wires[39]),
    .prog_clk_1_W_out(prog_clk_1_wires[58]),
    .prog_clk_1_E_out(prog_clk_1_wires[57]),
    .prog_clk_0_N_in(prog_clk_0_wires[118]),
    .pReset_E_in(pResetWires[270]),
    .pReset_N_out(pResetWires[269]),
    .pReset_W_out(pResetWires[267]),
    .chany_top_in(cby_1__1__29_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_29_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_29_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_29_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_29_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_29_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_29_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_29_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_29_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__37_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_40_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_40_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_40_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_40_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_40_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_40_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_40_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_40_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__28_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_28_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_28_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_28_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_28_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_28_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_28_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_28_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_28_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__26_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_28_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_28_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_28_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_28_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_28_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_28_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_28_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_28_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__37_ccff_tail[0]),
    .chany_top_out(sb_1__1__26_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__26_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__26_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__26_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__26_ccff_tail[0])
  );


  sb_1__1_
  sb_3__6_
  (
    .clk_3_W_out(clk_3_wires[50]),
    .clk_3_E_in(clk_3_wires[47]),
    .prog_clk_3_W_out(prog_clk_3_wires[50]),
    .prog_clk_3_E_in(prog_clk_3_wires[47]),
    .prog_clk_0_N_in(prog_clk_0_wires[121]),
    .pReset_E_in(pResetWires[319]),
    .pReset_N_out(pResetWires[318]),
    .pReset_W_out(pResetWires[316]),
    .chany_top_in(cby_1__1__30_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_30_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_30_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_30_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_30_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_30_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_30_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_30_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_30_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__38_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_41_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_41_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_41_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_41_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_41_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_41_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_41_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_41_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__29_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_29_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_29_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_29_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_29_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_29_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_29_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_29_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_29_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__27_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_29_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_29_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_29_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_29_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_29_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_29_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_29_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_29_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__38_ccff_tail[0]),
    .chany_top_out(sb_1__1__27_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__27_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__27_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__27_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__27_ccff_tail[0])
  );


  sb_1__1_
  sb_3__7_
  (
    .clk_1_N_in(clk_2_wires[54]),
    .clk_1_W_out(clk_1_wires[65]),
    .clk_1_E_out(clk_1_wires[64]),
    .prog_clk_1_N_in(prog_clk_2_wires[54]),
    .prog_clk_1_W_out(prog_clk_1_wires[65]),
    .prog_clk_1_E_out(prog_clk_1_wires[64]),
    .prog_clk_0_N_in(prog_clk_0_wires[124]),
    .pReset_E_in(pResetWires[368]),
    .pReset_N_out(pResetWires[367]),
    .pReset_W_out(pResetWires[365]),
    .chany_top_in(cby_1__1__31_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_31_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_31_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_31_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_31_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_31_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_31_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_31_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_31_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__39_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_42_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_42_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_42_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_42_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_42_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_42_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_42_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_42_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__30_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_30_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_30_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_30_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_30_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_30_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_30_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_30_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_30_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__28_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_30_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_30_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_30_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_30_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_30_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_30_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_30_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_30_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__39_ccff_tail[0]),
    .chany_top_out(sb_1__1__28_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__28_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__28_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__28_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__28_ccff_tail[0])
  );


  sb_1__1_
  sb_3__8_
  (
    .clk_2_S_out(clk_2_wires[53]),
    .clk_2_N_out(clk_2_wires[51]),
    .clk_2_E_in(clk_2_wires[50]),
    .prog_clk_2_S_out(prog_clk_2_wires[53]),
    .prog_clk_2_N_out(prog_clk_2_wires[51]),
    .prog_clk_2_E_in(prog_clk_2_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[127]),
    .pReset_E_in(pResetWires[417]),
    .pReset_N_out(pResetWires[416]),
    .pReset_W_out(pResetWires[414]),
    .chany_top_in(cby_1__1__32_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_32_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_32_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_32_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_32_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_32_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_32_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_32_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_32_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__40_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_43_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_43_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_43_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_43_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_43_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_43_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_43_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_43_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__31_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_31_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_31_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_31_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_31_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_31_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_31_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_31_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_31_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__29_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_31_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_31_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_31_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_31_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_31_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_31_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_31_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_31_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__40_ccff_tail[0]),
    .chany_top_out(sb_1__1__29_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__29_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__29_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__29_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__29_ccff_tail[0])
  );


  sb_1__1_
  sb_3__9_
  (
    .clk_1_S_in(clk_2_wires[52]),
    .clk_1_W_out(clk_1_wires[72]),
    .clk_1_E_out(clk_1_wires[71]),
    .prog_clk_1_S_in(prog_clk_2_wires[52]),
    .prog_clk_1_W_out(prog_clk_1_wires[72]),
    .prog_clk_1_E_out(prog_clk_1_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[130]),
    .pReset_E_in(pResetWires[466]),
    .pReset_N_out(pResetWires[465]),
    .pReset_W_out(pResetWires[463]),
    .chany_top_in(cby_1__1__33_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_33_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_33_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_33_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_33_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_33_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_33_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_33_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_33_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__41_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_44_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_44_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_44_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_44_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_44_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_44_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_44_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_44_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__32_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_32_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_32_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_32_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_32_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_32_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_32_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_32_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_32_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__30_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_32_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_32_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_32_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_32_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_32_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_32_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_32_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_32_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__41_ccff_tail[0]),
    .chany_top_out(sb_1__1__30_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__30_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__30_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__30_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__30_ccff_tail[0])
  );


  sb_1__1_
  sb_3__10_
  (
    .clk_2_N_out(clk_2_wires[64]),
    .clk_2_E_in(clk_2_wires[63]),
    .prog_clk_2_N_out(prog_clk_2_wires[64]),
    .prog_clk_2_E_in(prog_clk_2_wires[63]),
    .prog_clk_0_N_in(prog_clk_0_wires[133]),
    .pReset_E_in(pResetWires[515]),
    .pReset_N_out(pResetWires[514]),
    .pReset_W_out(pResetWires[512]),
    .chany_top_in(cby_1__1__34_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_34_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_34_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_34_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_34_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_34_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_34_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_34_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_34_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__42_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_45_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_45_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_45_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_45_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_45_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_45_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_45_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_45_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__33_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_33_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_33_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_33_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_33_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_33_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_33_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_33_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_33_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__31_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_33_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_33_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_33_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_33_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_33_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_33_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_33_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_33_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__42_ccff_tail[0]),
    .chany_top_out(sb_1__1__31_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__31_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__31_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__31_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__31_ccff_tail[0])
  );


  sb_1__1_
  sb_3__11_
  (
    .clk_1_S_in(clk_2_wires[65]),
    .clk_1_W_out(clk_1_wires[79]),
    .clk_1_E_out(clk_1_wires[78]),
    .prog_clk_1_S_in(prog_clk_2_wires[65]),
    .prog_clk_1_W_out(prog_clk_1_wires[79]),
    .prog_clk_1_E_out(prog_clk_1_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[136]),
    .pReset_E_in(pResetWires[564]),
    .pReset_N_out(pResetWires[563]),
    .pReset_W_out(pResetWires[561]),
    .chany_top_in(cby_1__1__35_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_35_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_35_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_35_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_35_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_35_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_35_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_35_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_35_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__43_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_46_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_46_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_46_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_46_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_46_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_46_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_46_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_46_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__34_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_34_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_34_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_34_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_34_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_34_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_34_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_34_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_34_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__32_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_34_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_34_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_34_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_34_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_34_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_34_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_34_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_34_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__43_ccff_tail[0]),
    .chany_top_out(sb_1__1__32_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__32_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__32_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__32_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__32_ccff_tail[0])
  );


  sb_1__1_
  sb_4__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[144]),
    .pReset_E_in(pResetWires[78]),
    .pReset_N_out(pResetWires[77]),
    .pReset_W_out(pResetWires[75]),
    .chany_top_in(cby_1__1__37_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_37_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_37_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_37_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_37_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_37_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_37_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_37_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_37_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__44_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_48_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_48_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_48_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_48_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_48_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_48_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_48_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_48_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__36_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_36_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_36_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_36_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_36_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_36_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_36_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_36_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_36_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__33_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_36_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_36_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_36_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_36_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_36_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_36_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_36_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_36_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__44_ccff_tail[0]),
    .chany_top_out(sb_1__1__33_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__33_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__33_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__33_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__33_ccff_tail[0])
  );


  sb_1__1_
  sb_4__2_
  (
    .clk_2_N_in(clk_3_wires[25]),
    .clk_2_W_out(clk_2_wires[27]),
    .clk_2_E_out(clk_2_wires[25]),
    .prog_clk_2_N_in(prog_clk_3_wires[25]),
    .prog_clk_2_W_out(prog_clk_2_wires[27]),
    .prog_clk_2_E_out(prog_clk_2_wires[25]),
    .prog_clk_0_N_in(prog_clk_0_wires[147]),
    .pReset_E_in(pResetWires[127]),
    .pReset_N_out(pResetWires[126]),
    .pReset_W_out(pResetWires[124]),
    .chany_top_in(cby_1__1__38_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_38_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_38_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_38_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_38_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_38_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_38_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_38_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_38_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__45_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_49_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_49_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_49_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_49_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_49_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_49_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_49_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_49_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__37_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_37_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_37_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_37_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_37_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_37_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_37_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_37_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_37_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__34_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_37_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_37_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_37_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_37_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_37_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_37_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_37_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_37_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__45_ccff_tail[0]),
    .chany_top_out(sb_1__1__34_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__34_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__34_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__34_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__34_ccff_tail[0])
  );


  sb_1__1_
  sb_4__3_
  (
    .clk_3_S_out(clk_3_wires[24]),
    .clk_3_N_in(clk_3_wires[21]),
    .prog_clk_3_S_out(prog_clk_3_wires[24]),
    .prog_clk_3_N_in(prog_clk_3_wires[21]),
    .prog_clk_0_N_in(prog_clk_0_wires[150]),
    .pReset_E_in(pResetWires[176]),
    .pReset_N_out(pResetWires[175]),
    .pReset_W_out(pResetWires[173]),
    .chany_top_in(cby_1__1__39_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_39_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_39_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_39_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_39_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_39_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_39_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_39_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_39_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__46_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_50_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_50_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_50_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_50_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_50_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_50_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_50_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_50_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__38_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_38_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_38_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_38_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_38_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_38_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_38_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_38_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_38_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__35_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_38_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_38_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_38_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_38_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_38_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_38_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_38_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_38_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__46_ccff_tail[0]),
    .chany_top_out(sb_1__1__35_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__35_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__35_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__35_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__35_ccff_tail[0])
  );


  sb_1__1_
  sb_4__4_
  (
    .clk_3_S_out(clk_3_wires[20]),
    .clk_2_N_in(clk_3_wires[15]),
    .clk_3_N_in(clk_3_wires[15]),
    .clk_2_W_out(clk_2_wires[36]),
    .clk_2_E_out(clk_2_wires[34]),
    .prog_clk_3_S_out(prog_clk_3_wires[20]),
    .prog_clk_2_N_in(prog_clk_3_wires[15]),
    .prog_clk_3_N_in(prog_clk_3_wires[15]),
    .prog_clk_2_W_out(prog_clk_2_wires[36]),
    .prog_clk_2_E_out(prog_clk_2_wires[34]),
    .prog_clk_0_N_in(prog_clk_0_wires[153]),
    .pReset_E_in(pResetWires[225]),
    .pReset_N_out(pResetWires[224]),
    .pReset_W_out(pResetWires[222]),
    .chany_top_in(cby_1__1__40_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_40_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_40_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_40_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_40_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_40_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_40_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_40_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_40_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__47_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_51_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_51_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_51_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_51_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_51_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_51_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_51_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_51_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__39_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_39_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_39_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_39_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_39_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_39_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_39_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_39_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_39_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__36_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_39_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_39_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_39_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_39_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_39_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_39_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_39_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_39_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__47_ccff_tail[0]),
    .chany_top_out(sb_1__1__36_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__36_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__36_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__36_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__36_ccff_tail[0])
  );


  sb_1__1_
  sb_4__5_
  (
    .clk_3_S_out(clk_3_wires[14]),
    .clk_3_N_in(clk_3_wires[11]),
    .prog_clk_3_S_out(prog_clk_3_wires[14]),
    .prog_clk_3_N_in(prog_clk_3_wires[11]),
    .prog_clk_0_N_in(prog_clk_0_wires[156]),
    .pReset_E_in(pResetWires[274]),
    .pReset_N_out(pResetWires[273]),
    .pReset_W_out(pResetWires[271]),
    .chany_top_in(cby_1__1__41_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_41_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_41_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_41_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_41_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_41_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_41_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_41_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_41_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__48_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_52_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_52_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_52_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_52_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_52_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_52_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_52_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_52_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__40_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_40_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_40_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_40_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_40_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_40_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_40_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_40_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_40_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__37_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_40_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_40_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_40_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_40_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_40_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_40_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_40_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_40_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__48_ccff_tail[0]),
    .chany_top_out(sb_1__1__37_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__37_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__37_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__37_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__37_ccff_tail[0])
  );


  sb_1__1_
  sb_4__6_
  (
    .clk_3_W_out(clk_3_wires[46]),
    .clk_3_S_out(clk_3_wires[10]),
    .clk_3_N_out(clk_3_wires[8]),
    .clk_3_E_in(clk_3_wires[7]),
    .prog_clk_3_W_out(prog_clk_3_wires[46]),
    .prog_clk_3_S_out(prog_clk_3_wires[10]),
    .prog_clk_3_N_out(prog_clk_3_wires[8]),
    .prog_clk_3_E_in(prog_clk_3_wires[7]),
    .prog_clk_0_N_in(prog_clk_0_wires[159]),
    .pReset_E_in(pResetWires[323]),
    .pReset_N_out(pResetWires[322]),
    .pReset_W_out(pResetWires[320]),
    .chany_top_in(cby_1__1__42_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_42_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_42_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_42_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_42_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_42_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_42_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_42_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_42_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__49_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_53_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_53_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_53_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_53_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_53_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_53_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_53_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_53_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__41_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_41_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_41_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_41_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_41_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_41_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_41_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_41_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_41_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__38_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_41_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_41_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_41_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_41_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_41_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_41_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_41_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_41_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__49_ccff_tail[0]),
    .chany_top_out(sb_1__1__38_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__38_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__38_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__38_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__38_ccff_tail[0])
  );


  sb_1__1_
  sb_4__7_
  (
    .clk_3_N_out(clk_3_wires[12]),
    .clk_3_S_in(clk_3_wires[9]),
    .prog_clk_3_N_out(prog_clk_3_wires[12]),
    .prog_clk_3_S_in(prog_clk_3_wires[9]),
    .prog_clk_0_N_in(prog_clk_0_wires[162]),
    .pReset_E_in(pResetWires[372]),
    .pReset_N_out(pResetWires[371]),
    .pReset_W_out(pResetWires[369]),
    .chany_top_in(cby_1__1__43_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_43_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_43_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_43_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_43_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_43_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_43_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_43_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_43_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__50_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_54_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_54_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_54_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_54_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_54_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_54_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_54_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_54_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__42_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_42_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_42_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_42_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_42_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_42_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_42_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_42_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_42_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__39_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_42_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_42_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_42_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_42_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_42_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_42_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_42_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_42_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__50_ccff_tail[0]),
    .chany_top_out(sb_1__1__39_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__39_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__39_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__39_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__39_ccff_tail[0])
  );


  sb_1__1_
  sb_4__8_
  (
    .clk_3_N_out(clk_3_wires[18]),
    .clk_2_S_in(clk_3_wires[13]),
    .clk_3_S_in(clk_3_wires[13]),
    .clk_2_W_out(clk_2_wires[49]),
    .clk_2_E_out(clk_2_wires[47]),
    .prog_clk_3_N_out(prog_clk_3_wires[18]),
    .prog_clk_2_S_in(prog_clk_3_wires[13]),
    .prog_clk_3_S_in(prog_clk_3_wires[13]),
    .prog_clk_2_W_out(prog_clk_2_wires[49]),
    .prog_clk_2_E_out(prog_clk_2_wires[47]),
    .prog_clk_0_N_in(prog_clk_0_wires[165]),
    .pReset_E_in(pResetWires[421]),
    .pReset_N_out(pResetWires[420]),
    .pReset_W_out(pResetWires[418]),
    .chany_top_in(cby_1__1__44_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_44_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_44_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_44_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_44_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_44_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_44_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_44_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_44_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__51_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_55_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_55_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_55_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_55_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_55_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_55_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_55_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_55_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__43_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_43_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_43_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_43_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_43_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_43_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_43_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_43_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_43_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__40_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_43_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_43_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_43_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_43_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_43_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_43_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_43_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_43_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__51_ccff_tail[0]),
    .chany_top_out(sb_1__1__40_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__40_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__40_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__40_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__40_ccff_tail[0])
  );


  sb_1__1_
  sb_4__9_
  (
    .clk_3_N_out(clk_3_wires[22]),
    .clk_3_S_in(clk_3_wires[19]),
    .prog_clk_3_N_out(prog_clk_3_wires[22]),
    .prog_clk_3_S_in(prog_clk_3_wires[19]),
    .prog_clk_0_N_in(prog_clk_0_wires[168]),
    .pReset_E_in(pResetWires[470]),
    .pReset_N_out(pResetWires[469]),
    .pReset_W_out(pResetWires[467]),
    .chany_top_in(cby_1__1__45_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_45_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_45_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_45_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_45_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_45_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_45_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_45_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_45_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__52_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_56_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_56_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_56_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_56_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_56_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_56_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_56_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_56_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__44_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_44_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_44_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_44_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_44_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_44_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_44_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_44_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_44_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__41_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_44_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_44_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_44_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_44_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_44_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_44_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_44_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_44_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__52_ccff_tail[0]),
    .chany_top_out(sb_1__1__41_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__41_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__41_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__41_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__41_ccff_tail[0])
  );


  sb_1__1_
  sb_4__10_
  (
    .clk_2_S_in(clk_3_wires[23]),
    .clk_2_W_out(clk_2_wires[62]),
    .clk_2_E_out(clk_2_wires[60]),
    .prog_clk_2_S_in(prog_clk_3_wires[23]),
    .prog_clk_2_W_out(prog_clk_2_wires[62]),
    .prog_clk_2_E_out(prog_clk_2_wires[60]),
    .prog_clk_0_N_in(prog_clk_0_wires[171]),
    .pReset_E_in(pResetWires[519]),
    .pReset_N_out(pResetWires[518]),
    .pReset_W_out(pResetWires[516]),
    .chany_top_in(cby_1__1__46_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_46_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_46_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_46_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_46_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_46_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_46_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_46_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_46_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__53_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_57_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_57_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_57_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_57_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_57_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_57_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_57_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_57_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__45_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_45_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_45_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_45_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_45_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_45_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_45_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_45_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_45_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__42_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_45_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_45_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_45_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_45_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_45_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_45_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_45_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_45_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__53_ccff_tail[0]),
    .chany_top_out(sb_1__1__42_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__42_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__42_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__42_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__42_ccff_tail[0])
  );


  sb_1__1_
  sb_4__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[174]),
    .pReset_E_in(pResetWires[568]),
    .pReset_N_out(pResetWires[567]),
    .pReset_W_out(pResetWires[565]),
    .chany_top_in(cby_1__1__47_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_47_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_47_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_47_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_47_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_47_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_47_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_47_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_47_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__54_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_58_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_58_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_58_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_58_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_58_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_58_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_58_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_58_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__46_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_46_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_46_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_46_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_46_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_46_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_46_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_46_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_46_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__43_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_46_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_46_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_46_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_46_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_46_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_46_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_46_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_46_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__54_ccff_tail[0]),
    .chany_top_out(sb_1__1__43_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__43_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__43_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__43_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__43_ccff_tail[0])
  );


  sb_1__1_
  sb_5__1_
  (
    .clk_1_N_in(clk_2_wires[32]),
    .clk_1_W_out(clk_1_wires[86]),
    .clk_1_E_out(clk_1_wires[85]),
    .prog_clk_1_N_in(prog_clk_2_wires[32]),
    .prog_clk_1_W_out(prog_clk_1_wires[86]),
    .prog_clk_1_E_out(prog_clk_1_wires[85]),
    .prog_clk_0_N_in(prog_clk_0_wires[182]),
    .pReset_E_in(pResetWires[82]),
    .pReset_N_out(pResetWires[81]),
    .pReset_W_out(pResetWires[79]),
    .chany_top_in(cby_1__1__49_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_49_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_49_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_49_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_49_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_49_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_49_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_49_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_49_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__55_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_60_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_60_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_60_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_60_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_60_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_60_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_60_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_60_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__48_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_48_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_48_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_48_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_48_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_48_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_48_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_48_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_48_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__44_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_48_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_48_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_48_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_48_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_48_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_48_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_48_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_48_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__55_ccff_tail[0]),
    .chany_top_out(sb_1__1__44_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__44_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__44_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__44_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__44_ccff_tail[0])
  );


  sb_1__1_
  sb_5__2_
  (
    .clk_2_S_out(clk_2_wires[31]),
    .clk_2_W_in(clk_2_wires[26]),
    .prog_clk_2_S_out(prog_clk_2_wires[31]),
    .prog_clk_2_W_in(prog_clk_2_wires[26]),
    .prog_clk_0_N_in(prog_clk_0_wires[185]),
    .pReset_E_in(pResetWires[131]),
    .pReset_N_out(pResetWires[130]),
    .pReset_W_out(pResetWires[128]),
    .chany_top_in(cby_1__1__50_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_50_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_50_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_50_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_50_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_50_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_50_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_50_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_50_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__56_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_61_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_61_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_61_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_61_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_61_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_61_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_61_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_61_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__49_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_49_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_49_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_49_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_49_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_49_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_49_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_49_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_49_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__45_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_49_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_49_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_49_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_49_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_49_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_49_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_49_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_49_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__56_ccff_tail[0]),
    .chany_top_out(sb_1__1__45_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__45_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__45_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__45_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__45_ccff_tail[0])
  );


  sb_1__1_
  sb_5__3_
  (
    .clk_1_N_in(clk_2_wires[45]),
    .clk_1_W_out(clk_1_wires[93]),
    .clk_1_E_out(clk_1_wires[92]),
    .prog_clk_1_N_in(prog_clk_2_wires[45]),
    .prog_clk_1_W_out(prog_clk_1_wires[93]),
    .prog_clk_1_E_out(prog_clk_1_wires[92]),
    .prog_clk_0_N_in(prog_clk_0_wires[188]),
    .pReset_E_in(pResetWires[180]),
    .pReset_N_out(pResetWires[179]),
    .pReset_W_out(pResetWires[177]),
    .chany_top_in(cby_1__1__51_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_51_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_51_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_51_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_51_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_51_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_51_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_51_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_51_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__57_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_62_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_62_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_62_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_62_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_62_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_62_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_62_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_62_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__50_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_50_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_50_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_50_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_50_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_50_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_50_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_50_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_50_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__46_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_50_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_50_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_50_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_50_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_50_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_50_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_50_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_50_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__57_ccff_tail[0]),
    .chany_top_out(sb_1__1__46_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__46_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__46_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__46_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__46_ccff_tail[0])
  );


  sb_1__1_
  sb_5__4_
  (
    .clk_2_S_out(clk_2_wires[44]),
    .clk_2_N_out(clk_2_wires[42]),
    .clk_2_W_in(clk_2_wires[35]),
    .prog_clk_2_S_out(prog_clk_2_wires[44]),
    .prog_clk_2_N_out(prog_clk_2_wires[42]),
    .prog_clk_2_W_in(prog_clk_2_wires[35]),
    .prog_clk_0_N_in(prog_clk_0_wires[191]),
    .pReset_E_in(pResetWires[229]),
    .pReset_N_out(pResetWires[228]),
    .pReset_W_out(pResetWires[226]),
    .chany_top_in(cby_1__1__52_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_52_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_52_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_52_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_52_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_52_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_52_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_52_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_52_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__58_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_63_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_63_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_63_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_63_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_63_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_63_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_63_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_63_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__51_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_51_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_51_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_51_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_51_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_51_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_51_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_51_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_51_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__47_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_51_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_51_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_51_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_51_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_51_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_51_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_51_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_51_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__58_ccff_tail[0]),
    .chany_top_out(sb_1__1__47_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__47_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__47_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__47_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__47_ccff_tail[0])
  );


  sb_1__1_
  sb_5__5_
  (
    .clk_1_S_in(clk_2_wires[43]),
    .clk_1_W_out(clk_1_wires[100]),
    .clk_1_E_out(clk_1_wires[99]),
    .prog_clk_1_S_in(prog_clk_2_wires[43]),
    .prog_clk_1_W_out(prog_clk_1_wires[100]),
    .prog_clk_1_E_out(prog_clk_1_wires[99]),
    .prog_clk_0_N_in(prog_clk_0_wires[194]),
    .pReset_E_in(pResetWires[278]),
    .pReset_N_out(pResetWires[277]),
    .pReset_W_out(pResetWires[275]),
    .chany_top_in(cby_1__1__53_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_53_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_53_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_53_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_53_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_53_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_53_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_53_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_53_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__59_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_64_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_64_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_64_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_64_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_64_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_64_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_64_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_64_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__52_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_52_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_52_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_52_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_52_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_52_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_52_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_52_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_52_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__48_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_52_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_52_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_52_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_52_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_52_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_52_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_52_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_52_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__59_ccff_tail[0]),
    .chany_top_out(sb_1__1__48_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__48_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__48_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__48_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__48_ccff_tail[0])
  );


  sb_1__1_
  sb_5__6_
  (
    .clk_3_W_out(clk_3_wires[6]),
    .clk_3_E_in(clk_3_wires[3]),
    .prog_clk_3_W_out(prog_clk_3_wires[6]),
    .prog_clk_3_E_in(prog_clk_3_wires[3]),
    .prog_clk_0_N_in(prog_clk_0_wires[197]),
    .pReset_E_in(pResetWires[327]),
    .pReset_N_out(pResetWires[326]),
    .pReset_W_out(pResetWires[324]),
    .chany_top_in(cby_1__1__54_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_54_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_54_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_54_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_54_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_54_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_54_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_54_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_54_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__60_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_65_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_65_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_65_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_65_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_65_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_65_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_65_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_65_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__53_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_53_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_53_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_53_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_53_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_53_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_53_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_53_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_53_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__49_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_53_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_53_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_53_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_53_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_53_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_53_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_53_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_53_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__60_ccff_tail[0]),
    .chany_top_out(sb_1__1__49_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__49_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__49_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__49_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__49_ccff_tail[0])
  );


  sb_1__1_
  sb_5__7_
  (
    .clk_1_N_in(clk_2_wires[58]),
    .clk_1_W_out(clk_1_wires[107]),
    .clk_1_E_out(clk_1_wires[106]),
    .prog_clk_1_N_in(prog_clk_2_wires[58]),
    .prog_clk_1_W_out(prog_clk_1_wires[107]),
    .prog_clk_1_E_out(prog_clk_1_wires[106]),
    .prog_clk_0_N_in(prog_clk_0_wires[200]),
    .pReset_E_in(pResetWires[376]),
    .pReset_N_out(pResetWires[375]),
    .pReset_W_out(pResetWires[373]),
    .chany_top_in(cby_1__1__55_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_55_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_55_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_55_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_55_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_55_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_55_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_55_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_55_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__61_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_66_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_66_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_66_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_66_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_66_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_66_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_66_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_66_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__54_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_54_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_54_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_54_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_54_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_54_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_54_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_54_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_54_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__50_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_54_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_54_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_54_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_54_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_54_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_54_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_54_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_54_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__61_ccff_tail[0]),
    .chany_top_out(sb_1__1__50_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__50_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__50_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__50_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__50_ccff_tail[0])
  );


  sb_1__1_
  sb_5__8_
  (
    .clk_2_S_out(clk_2_wires[57]),
    .clk_2_N_out(clk_2_wires[55]),
    .clk_2_W_in(clk_2_wires[48]),
    .prog_clk_2_S_out(prog_clk_2_wires[57]),
    .prog_clk_2_N_out(prog_clk_2_wires[55]),
    .prog_clk_2_W_in(prog_clk_2_wires[48]),
    .prog_clk_0_N_in(prog_clk_0_wires[203]),
    .pReset_E_in(pResetWires[425]),
    .pReset_N_out(pResetWires[424]),
    .pReset_W_out(pResetWires[422]),
    .chany_top_in(cby_1__1__56_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_56_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_56_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_56_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_56_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_56_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_56_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_56_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_56_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__62_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_67_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_67_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_67_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_67_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_67_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_67_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_67_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_67_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__55_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_55_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_55_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_55_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_55_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_55_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_55_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_55_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_55_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__51_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_55_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_55_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_55_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_55_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_55_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_55_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_55_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_55_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__62_ccff_tail[0]),
    .chany_top_out(sb_1__1__51_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__51_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__51_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__51_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__51_ccff_tail[0])
  );


  sb_1__1_
  sb_5__9_
  (
    .clk_1_S_in(clk_2_wires[56]),
    .clk_1_W_out(clk_1_wires[114]),
    .clk_1_E_out(clk_1_wires[113]),
    .prog_clk_1_S_in(prog_clk_2_wires[56]),
    .prog_clk_1_W_out(prog_clk_1_wires[114]),
    .prog_clk_1_E_out(prog_clk_1_wires[113]),
    .prog_clk_0_N_in(prog_clk_0_wires[206]),
    .pReset_E_in(pResetWires[474]),
    .pReset_N_out(pResetWires[473]),
    .pReset_W_out(pResetWires[471]),
    .chany_top_in(cby_1__1__57_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_57_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_57_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_57_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_57_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_57_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_57_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_57_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_57_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__63_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_68_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_68_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_68_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_68_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_68_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_68_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_68_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_68_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__56_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_56_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_56_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_56_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_56_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_56_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_56_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_56_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_56_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__52_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_56_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_56_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_56_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_56_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_56_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_56_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_56_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_56_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__63_ccff_tail[0]),
    .chany_top_out(sb_1__1__52_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__52_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__52_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__52_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__52_ccff_tail[0])
  );


  sb_1__1_
  sb_5__10_
  (
    .clk_2_N_out(clk_2_wires[66]),
    .clk_2_W_in(clk_2_wires[61]),
    .prog_clk_2_N_out(prog_clk_2_wires[66]),
    .prog_clk_2_W_in(prog_clk_2_wires[61]),
    .prog_clk_0_N_in(prog_clk_0_wires[209]),
    .pReset_E_in(pResetWires[523]),
    .pReset_N_out(pResetWires[522]),
    .pReset_W_out(pResetWires[520]),
    .chany_top_in(cby_1__1__58_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_58_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_58_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_58_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_58_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_58_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_58_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_58_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_58_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__64_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_69_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_69_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_69_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_69_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_69_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_69_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_69_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_69_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__57_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_57_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_57_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_57_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_57_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_57_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_57_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_57_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_57_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__53_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_57_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_57_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_57_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_57_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_57_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_57_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_57_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_57_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__64_ccff_tail[0]),
    .chany_top_out(sb_1__1__53_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__53_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__53_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__53_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__53_ccff_tail[0])
  );


  sb_1__1_
  sb_5__11_
  (
    .clk_1_S_in(clk_2_wires[67]),
    .clk_1_W_out(clk_1_wires[121]),
    .clk_1_E_out(clk_1_wires[120]),
    .prog_clk_1_S_in(prog_clk_2_wires[67]),
    .prog_clk_1_W_out(prog_clk_1_wires[121]),
    .prog_clk_1_E_out(prog_clk_1_wires[120]),
    .prog_clk_0_N_in(prog_clk_0_wires[212]),
    .pReset_E_in(pResetWires[572]),
    .pReset_N_out(pResetWires[571]),
    .pReset_W_out(pResetWires[569]),
    .chany_top_in(cby_1__1__59_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_59_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_59_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_59_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_59_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_59_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_59_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_59_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_59_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__65_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_70_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_70_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_70_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_70_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_70_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_70_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_70_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_70_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__58_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_58_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_58_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_58_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_58_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_58_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_58_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_58_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_58_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__54_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_58_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_58_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_58_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_58_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_58_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_58_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_58_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_58_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__65_ccff_tail[0]),
    .chany_top_out(sb_1__1__54_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__54_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__54_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__54_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__54_ccff_tail[0])
  );


  sb_1__1_
  sb_6__1_
  (
    .clk_3_N_out(clk_3_wires[92]),
    .clk_3_S_in(clk_3_wires[89]),
    .prog_clk_3_N_out(prog_clk_3_wires[92]),
    .prog_clk_3_S_in(prog_clk_3_wires[89]),
    .prog_clk_0_N_in(prog_clk_0_wires[220]),
    .Reset_N_out(ResetWires[3]),
    .Reset_S_in(ResetWires[2]),
    .pReset_E_out(pResetWires[86]),
    .pReset_W_out(pResetWires[83]),
    .pReset_N_out(pResetWires[85]),
    .pReset_S_in(pResetWires[2]),
    .Test_en_N_out(Test_enWires[3]),
    .Test_en_S_in(Test_enWires[2]),
    .chany_top_in(cby_1__1__61_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_61_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_61_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_61_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_61_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_61_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_61_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_61_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_61_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__66_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_72_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_72_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_72_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_72_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_72_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_72_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_72_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_72_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__60_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_60_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_60_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_60_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_60_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_60_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_60_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_60_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_60_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__55_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_60_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_60_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_60_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_60_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_60_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_60_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_60_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_60_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__66_ccff_tail[0]),
    .chany_top_out(sb_1__1__55_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__55_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__55_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__55_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__55_ccff_tail[0])
  );


  sb_1__1_
  sb_6__2_
  (
    .clk_3_N_out(clk_3_wires[94]),
    .clk_3_S_in(clk_3_wires[91]),
    .prog_clk_3_N_out(prog_clk_3_wires[94]),
    .prog_clk_3_S_in(prog_clk_3_wires[91]),
    .prog_clk_0_N_in(prog_clk_0_wires[223]),
    .Reset_N_out(ResetWires[5]),
    .Reset_S_in(ResetWires[4]),
    .pReset_E_out(pResetWires[135]),
    .pReset_W_out(pResetWires[132]),
    .pReset_N_out(pResetWires[134]),
    .pReset_S_in(pResetWires[4]),
    .Test_en_N_out(Test_enWires[5]),
    .Test_en_S_in(Test_enWires[4]),
    .chany_top_in(cby_1__1__62_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_62_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_62_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_62_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_62_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_62_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_62_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_62_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_62_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__67_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_73_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_73_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_73_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_73_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_73_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_73_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_73_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_73_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__61_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_61_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_61_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_61_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_61_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_61_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_61_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_61_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_61_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__56_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_61_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_61_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_61_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_61_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_61_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_61_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_61_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_61_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__67_ccff_tail[0]),
    .chany_top_out(sb_1__1__56_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__56_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__56_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__56_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__56_ccff_tail[0])
  );


  sb_1__1_
  sb_6__3_
  (
    .clk_3_N_out(clk_3_wires[96]),
    .clk_3_S_in(clk_3_wires[93]),
    .prog_clk_3_N_out(prog_clk_3_wires[96]),
    .prog_clk_3_S_in(prog_clk_3_wires[93]),
    .prog_clk_0_N_in(prog_clk_0_wires[226]),
    .Reset_N_out(ResetWires[7]),
    .Reset_S_in(ResetWires[6]),
    .pReset_E_out(pResetWires[184]),
    .pReset_W_out(pResetWires[181]),
    .pReset_N_out(pResetWires[183]),
    .pReset_S_in(pResetWires[6]),
    .Test_en_N_out(Test_enWires[7]),
    .Test_en_S_in(Test_enWires[6]),
    .chany_top_in(cby_1__1__63_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_63_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_63_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_63_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_63_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_63_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_63_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_63_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_63_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__68_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_74_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_74_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_74_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_74_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_74_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_74_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_74_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_74_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__62_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_62_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_62_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_62_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_62_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_62_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_62_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_62_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_62_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__57_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_62_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_62_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_62_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_62_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_62_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_62_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_62_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_62_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__68_ccff_tail[0]),
    .chany_top_out(sb_1__1__57_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__57_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__57_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__57_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__57_ccff_tail[0])
  );


  sb_1__1_
  sb_6__4_
  (
    .clk_3_N_out(clk_3_wires[98]),
    .clk_3_S_in(clk_3_wires[95]),
    .prog_clk_3_N_out(prog_clk_3_wires[98]),
    .prog_clk_3_S_in(prog_clk_3_wires[95]),
    .prog_clk_0_N_in(prog_clk_0_wires[229]),
    .Reset_N_out(ResetWires[9]),
    .Reset_S_in(ResetWires[8]),
    .pReset_E_out(pResetWires[233]),
    .pReset_W_out(pResetWires[230]),
    .pReset_N_out(pResetWires[232]),
    .pReset_S_in(pResetWires[8]),
    .Test_en_N_out(Test_enWires[9]),
    .Test_en_S_in(Test_enWires[8]),
    .chany_top_in(cby_1__1__64_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_64_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_64_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_64_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_64_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_64_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_64_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_64_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_64_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__69_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_75_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_75_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_75_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_75_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_75_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_75_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_75_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_75_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__63_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_63_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_63_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_63_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_63_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_63_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_63_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_63_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_63_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__58_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_63_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_63_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_63_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_63_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_63_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_63_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_63_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_63_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__69_ccff_tail[0]),
    .chany_top_out(sb_1__1__58_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__58_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__58_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__58_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__58_ccff_tail[0])
  );


  sb_1__1_
  sb_6__5_
  (
    .clk_3_N_out(clk_3_wires[100]),
    .clk_3_S_in(clk_3_wires[97]),
    .prog_clk_3_N_out(prog_clk_3_wires[100]),
    .prog_clk_3_S_in(prog_clk_3_wires[97]),
    .prog_clk_0_N_in(prog_clk_0_wires[232]),
    .Reset_N_out(ResetWires[11]),
    .Reset_S_in(ResetWires[10]),
    .pReset_E_out(pResetWires[282]),
    .pReset_W_out(pResetWires[279]),
    .pReset_N_out(pResetWires[281]),
    .pReset_S_in(pResetWires[10]),
    .Test_en_N_out(Test_enWires[11]),
    .Test_en_S_in(Test_enWires[10]),
    .chany_top_in(cby_1__1__65_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_65_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_65_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_65_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_65_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_65_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_65_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_65_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_65_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__70_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_76_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_76_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_76_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_76_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_76_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_76_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_76_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_76_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__64_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_64_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_64_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_64_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_64_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_64_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_64_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_64_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_64_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__59_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_64_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_64_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_64_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_64_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_64_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_64_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_64_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_64_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__70_ccff_tail[0]),
    .chany_top_out(sb_1__1__59_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__59_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__59_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__59_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__59_ccff_tail[0])
  );


  sb_1__1_
  sb_6__6_
  (
    .clk_3_S_in(clk_3_wires[99]),
    .clk_3_W_out(clk_3_wires[2]),
    .clk_3_E_out(clk_3_wires[0]),
    .prog_clk_3_S_in(prog_clk_3_wires[99]),
    .prog_clk_3_W_out(prog_clk_3_wires[2]),
    .prog_clk_3_E_out(prog_clk_3_wires[0]),
    .prog_clk_0_N_in(prog_clk_0_wires[235]),
    .Reset_N_out(ResetWires[13]),
    .Reset_S_in(ResetWires[12]),
    .pReset_E_out(pResetWires[331]),
    .pReset_W_out(pResetWires[328]),
    .pReset_N_out(pResetWires[330]),
    .pReset_S_in(pResetWires[12]),
    .Test_en_N_out(Test_enWires[13]),
    .Test_en_S_in(Test_enWires[12]),
    .chany_top_in(cby_1__1__66_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_66_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_66_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_66_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_66_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_66_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_66_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_66_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_66_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__71_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_77_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_77_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_77_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_77_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_77_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_77_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_77_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_77_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__65_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_65_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_65_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_65_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_65_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_65_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_65_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_65_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_65_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__60_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_65_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_65_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_65_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_65_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_65_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_65_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_65_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_65_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__71_ccff_tail[0]),
    .chany_top_out(sb_1__1__60_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__60_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__60_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__60_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__60_ccff_tail[0])
  );


  sb_1__1_
  sb_6__7_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[238]),
    .Reset_N_out(ResetWires[15]),
    .Reset_S_in(ResetWires[14]),
    .pReset_E_out(pResetWires[380]),
    .pReset_W_out(pResetWires[377]),
    .pReset_N_out(pResetWires[379]),
    .pReset_S_in(pResetWires[14]),
    .Test_en_N_out(Test_enWires[15]),
    .Test_en_S_in(Test_enWires[14]),
    .chany_top_in(cby_1__1__67_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_67_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_67_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_67_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_67_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_67_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_67_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_67_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_67_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__72_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_78_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_78_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_78_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_78_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_78_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_78_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_78_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_78_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__66_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_66_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_66_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_66_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_66_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_66_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_66_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_66_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_66_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__61_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_66_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_66_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_66_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_66_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_66_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_66_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_66_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_66_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__72_ccff_tail[0]),
    .chany_top_out(sb_1__1__61_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__61_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__61_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__61_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__61_ccff_tail[0])
  );


  sb_1__1_
  sb_6__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[241]),
    .Reset_N_out(ResetWires[17]),
    .Reset_S_in(ResetWires[16]),
    .pReset_E_out(pResetWires[429]),
    .pReset_W_out(pResetWires[426]),
    .pReset_N_out(pResetWires[428]),
    .pReset_S_in(pResetWires[16]),
    .Test_en_N_out(Test_enWires[17]),
    .Test_en_S_in(Test_enWires[16]),
    .chany_top_in(cby_1__1__68_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_68_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_68_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_68_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_68_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_68_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_68_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_68_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_68_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__73_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_79_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_79_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_79_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_79_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_79_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_79_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_79_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_79_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__67_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_67_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_67_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_67_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_67_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_67_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_67_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_67_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_67_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__62_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_67_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_67_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_67_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_67_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_67_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_67_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_67_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_67_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__73_ccff_tail[0]),
    .chany_top_out(sb_1__1__62_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__62_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__62_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__62_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__62_ccff_tail[0])
  );


  sb_1__1_
  sb_6__9_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[244]),
    .Reset_N_out(ResetWires[19]),
    .Reset_S_in(ResetWires[18]),
    .pReset_E_out(pResetWires[478]),
    .pReset_W_out(pResetWires[475]),
    .pReset_N_out(pResetWires[477]),
    .pReset_S_in(pResetWires[18]),
    .Test_en_N_out(Test_enWires[19]),
    .Test_en_S_in(Test_enWires[18]),
    .chany_top_in(cby_1__1__69_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_69_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_69_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_69_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_69_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_69_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_69_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_69_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_69_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__74_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_80_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_80_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_80_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_80_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_80_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_80_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_80_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_80_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__68_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_68_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_68_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_68_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_68_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_68_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_68_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_68_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_68_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__63_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_68_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_68_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_68_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_68_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_68_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_68_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_68_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_68_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__74_ccff_tail[0]),
    .chany_top_out(sb_1__1__63_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__63_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__63_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__63_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__63_ccff_tail[0])
  );


  sb_1__1_
  sb_6__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[247]),
    .Reset_N_out(ResetWires[21]),
    .Reset_S_in(ResetWires[20]),
    .pReset_E_out(pResetWires[527]),
    .pReset_W_out(pResetWires[524]),
    .pReset_N_out(pResetWires[526]),
    .pReset_S_in(pResetWires[20]),
    .Test_en_N_out(Test_enWires[21]),
    .Test_en_S_in(Test_enWires[20]),
    .chany_top_in(cby_1__1__70_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_70_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_70_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_70_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_70_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_70_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_70_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_70_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_70_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__75_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_81_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_81_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_81_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_81_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_81_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_81_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_81_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_81_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__69_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_69_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_69_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_69_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_69_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_69_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_69_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_69_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_69_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__64_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_69_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_69_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_69_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_69_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_69_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_69_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_69_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_69_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__75_ccff_tail[0]),
    .chany_top_out(sb_1__1__64_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__64_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__64_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__64_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__64_ccff_tail[0])
  );


  sb_1__1_
  sb_6__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[250]),
    .Reset_N_out(ResetWires[23]),
    .Reset_S_in(ResetWires[22]),
    .pReset_E_out(pResetWires[576]),
    .pReset_W_out(pResetWires[573]),
    .pReset_N_out(pResetWires[575]),
    .pReset_S_in(pResetWires[22]),
    .Test_en_N_out(Test_enWires[23]),
    .Test_en_S_in(Test_enWires[22]),
    .chany_top_in(cby_1__1__71_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_71_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_71_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_71_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_71_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_71_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_71_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_71_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_71_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__76_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_82_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_82_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_82_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_82_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_82_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_82_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_82_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_82_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__70_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_70_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_70_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_70_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_70_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_70_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_70_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_70_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_70_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__65_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_70_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_70_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_70_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_70_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_70_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_70_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_70_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_70_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__76_ccff_tail[0]),
    .chany_top_out(sb_1__1__65_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__65_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__65_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__65_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__65_ccff_tail[0])
  );


  sb_1__1_
  sb_7__1_
  (
    .clk_1_N_in(clk_2_wires[74]),
    .clk_1_W_out(clk_1_wires[128]),
    .clk_1_E_out(clk_1_wires[127]),
    .prog_clk_1_N_in(prog_clk_2_wires[74]),
    .prog_clk_1_W_out(prog_clk_1_wires[128]),
    .prog_clk_1_E_out(prog_clk_1_wires[127]),
    .prog_clk_0_N_in(prog_clk_0_wires[258]),
    .pReset_E_out(pResetWires[90]),
    .pReset_N_out(pResetWires[89]),
    .pReset_W_in(pResetWires[87]),
    .chany_top_in(cby_1__1__73_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_73_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_73_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_73_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_73_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_73_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_73_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_73_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_73_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__77_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_84_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_84_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_84_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_84_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_84_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_84_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_84_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_84_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__72_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_72_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_72_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_72_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_72_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_72_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_72_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_72_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_72_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__66_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_72_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_72_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_72_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_72_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_72_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_72_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_72_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_72_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__77_ccff_tail[0]),
    .chany_top_out(sb_1__1__66_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__66_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__66_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__66_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__66_ccff_tail[0])
  );


  sb_1__1_
  sb_7__2_
  (
    .clk_2_S_out(clk_2_wires[73]),
    .clk_2_E_in(clk_2_wires[72]),
    .prog_clk_2_S_out(prog_clk_2_wires[73]),
    .prog_clk_2_E_in(prog_clk_2_wires[72]),
    .prog_clk_0_N_in(prog_clk_0_wires[261]),
    .pReset_E_out(pResetWires[139]),
    .pReset_N_out(pResetWires[138]),
    .pReset_W_in(pResetWires[136]),
    .chany_top_in(cby_1__1__74_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_74_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_74_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_74_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_74_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_74_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_74_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_74_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_74_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__78_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_85_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_85_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_85_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_85_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_85_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_85_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_85_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_85_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__73_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_73_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_73_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_73_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_73_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_73_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_73_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_73_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_73_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__67_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_73_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_73_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_73_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_73_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_73_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_73_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_73_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_73_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__78_ccff_tail[0]),
    .chany_top_out(sb_1__1__67_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__67_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__67_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__67_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__67_ccff_tail[0])
  );


  sb_1__1_
  sb_7__3_
  (
    .clk_1_N_in(clk_2_wires[85]),
    .clk_1_W_out(clk_1_wires[135]),
    .clk_1_E_out(clk_1_wires[134]),
    .prog_clk_1_N_in(prog_clk_2_wires[85]),
    .prog_clk_1_W_out(prog_clk_1_wires[135]),
    .prog_clk_1_E_out(prog_clk_1_wires[134]),
    .prog_clk_0_N_in(prog_clk_0_wires[264]),
    .pReset_E_out(pResetWires[188]),
    .pReset_N_out(pResetWires[187]),
    .pReset_W_in(pResetWires[185]),
    .chany_top_in(cby_1__1__75_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_75_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_75_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_75_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_75_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_75_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_75_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_75_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_75_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__79_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_86_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_86_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_86_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_86_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_86_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_86_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_86_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_86_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__74_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_74_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_74_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_74_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_74_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_74_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_74_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_74_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_74_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__68_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_74_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_74_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_74_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_74_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_74_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_74_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_74_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_74_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__79_ccff_tail[0]),
    .chany_top_out(sb_1__1__68_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__68_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__68_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__68_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__68_ccff_tail[0])
  );


  sb_1__1_
  sb_7__4_
  (
    .clk_2_S_out(clk_2_wires[84]),
    .clk_2_N_out(clk_2_wires[82]),
    .clk_2_E_in(clk_2_wires[81]),
    .prog_clk_2_S_out(prog_clk_2_wires[84]),
    .prog_clk_2_N_out(prog_clk_2_wires[82]),
    .prog_clk_2_E_in(prog_clk_2_wires[81]),
    .prog_clk_0_N_in(prog_clk_0_wires[267]),
    .pReset_E_out(pResetWires[237]),
    .pReset_N_out(pResetWires[236]),
    .pReset_W_in(pResetWires[234]),
    .chany_top_in(cby_1__1__76_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_76_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_76_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_76_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_76_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_76_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_76_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_76_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_76_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__80_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_87_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_87_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_87_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_87_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_87_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_87_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_87_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_87_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__75_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_75_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_75_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_75_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_75_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_75_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_75_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_75_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_75_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__69_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_75_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_75_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_75_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_75_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_75_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_75_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_75_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_75_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__80_ccff_tail[0]),
    .chany_top_out(sb_1__1__69_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__69_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__69_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__69_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__69_ccff_tail[0])
  );


  sb_1__1_
  sb_7__5_
  (
    .clk_1_S_in(clk_2_wires[83]),
    .clk_1_W_out(clk_1_wires[142]),
    .clk_1_E_out(clk_1_wires[141]),
    .prog_clk_1_S_in(prog_clk_2_wires[83]),
    .prog_clk_1_W_out(prog_clk_1_wires[142]),
    .prog_clk_1_E_out(prog_clk_1_wires[141]),
    .prog_clk_0_N_in(prog_clk_0_wires[270]),
    .pReset_E_out(pResetWires[286]),
    .pReset_N_out(pResetWires[285]),
    .pReset_W_in(pResetWires[283]),
    .chany_top_in(cby_1__1__77_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_77_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_77_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_77_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_77_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_77_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_77_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_77_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_77_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__81_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_88_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_88_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_88_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_88_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_88_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_88_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_88_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_88_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__76_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_76_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_76_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_76_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_76_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_76_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_76_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_76_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_76_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__70_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_76_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_76_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_76_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_76_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_76_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_76_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_76_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_76_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__81_ccff_tail[0]),
    .chany_top_out(sb_1__1__70_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__70_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__70_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__70_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__70_ccff_tail[0])
  );


  sb_1__1_
  sb_7__6_
  (
    .clk_3_E_out(clk_3_wires[4]),
    .clk_3_W_in(clk_3_wires[1]),
    .prog_clk_3_E_out(prog_clk_3_wires[4]),
    .prog_clk_3_W_in(prog_clk_3_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[273]),
    .pReset_E_out(pResetWires[335]),
    .pReset_N_out(pResetWires[334]),
    .pReset_W_in(pResetWires[332]),
    .chany_top_in(cby_1__1__78_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_78_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_78_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_78_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_78_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_78_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_78_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_78_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_78_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__82_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_89_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_89_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_89_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_89_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_89_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_89_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_89_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_89_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__77_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_77_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_77_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_77_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_77_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_77_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_77_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_77_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_77_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__71_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_77_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_77_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_77_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_77_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_77_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_77_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_77_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_77_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__82_ccff_tail[0]),
    .chany_top_out(sb_1__1__71_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__71_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__71_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__71_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__71_ccff_tail[0])
  );


  sb_1__1_
  sb_7__7_
  (
    .clk_1_N_in(clk_2_wires[98]),
    .clk_1_W_out(clk_1_wires[149]),
    .clk_1_E_out(clk_1_wires[148]),
    .prog_clk_1_N_in(prog_clk_2_wires[98]),
    .prog_clk_1_W_out(prog_clk_1_wires[149]),
    .prog_clk_1_E_out(prog_clk_1_wires[148]),
    .prog_clk_0_N_in(prog_clk_0_wires[276]),
    .pReset_E_out(pResetWires[384]),
    .pReset_N_out(pResetWires[383]),
    .pReset_W_in(pResetWires[381]),
    .chany_top_in(cby_1__1__79_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_79_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_79_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_79_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_79_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_79_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_79_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_79_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_79_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__83_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_90_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_90_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_90_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_90_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_90_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_90_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_90_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_90_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__78_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_78_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_78_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_78_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_78_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_78_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_78_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_78_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_78_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__72_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_78_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_78_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_78_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_78_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_78_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_78_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_78_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_78_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__83_ccff_tail[0]),
    .chany_top_out(sb_1__1__72_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__72_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__72_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__72_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__72_ccff_tail[0])
  );


  sb_1__1_
  sb_7__8_
  (
    .clk_2_S_out(clk_2_wires[97]),
    .clk_2_N_out(clk_2_wires[95]),
    .clk_2_E_in(clk_2_wires[94]),
    .prog_clk_2_S_out(prog_clk_2_wires[97]),
    .prog_clk_2_N_out(prog_clk_2_wires[95]),
    .prog_clk_2_E_in(prog_clk_2_wires[94]),
    .prog_clk_0_N_in(prog_clk_0_wires[279]),
    .pReset_E_out(pResetWires[433]),
    .pReset_N_out(pResetWires[432]),
    .pReset_W_in(pResetWires[430]),
    .chany_top_in(cby_1__1__80_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_80_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_80_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_80_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_80_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_80_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_80_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_80_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_80_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__84_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_91_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_91_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_91_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_91_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_91_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_91_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_91_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_91_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__79_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_79_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_79_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_79_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_79_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_79_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_79_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_79_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_79_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__73_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_79_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_79_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_79_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_79_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_79_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_79_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_79_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_79_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__84_ccff_tail[0]),
    .chany_top_out(sb_1__1__73_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__73_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__73_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__73_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__73_ccff_tail[0])
  );


  sb_1__1_
  sb_7__9_
  (
    .clk_1_S_in(clk_2_wires[96]),
    .clk_1_W_out(clk_1_wires[156]),
    .clk_1_E_out(clk_1_wires[155]),
    .prog_clk_1_S_in(prog_clk_2_wires[96]),
    .prog_clk_1_W_out(prog_clk_1_wires[156]),
    .prog_clk_1_E_out(prog_clk_1_wires[155]),
    .prog_clk_0_N_in(prog_clk_0_wires[282]),
    .pReset_E_out(pResetWires[482]),
    .pReset_N_out(pResetWires[481]),
    .pReset_W_in(pResetWires[479]),
    .chany_top_in(cby_1__1__81_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_81_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_81_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_81_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_81_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_81_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_81_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_81_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_81_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__85_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_92_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_92_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_92_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_92_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_92_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_92_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_92_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_92_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__80_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_80_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_80_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_80_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_80_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_80_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_80_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_80_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_80_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__74_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_80_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_80_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_80_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_80_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_80_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_80_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_80_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_80_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__85_ccff_tail[0]),
    .chany_top_out(sb_1__1__74_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__74_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__74_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__74_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__74_ccff_tail[0])
  );


  sb_1__1_
  sb_7__10_
  (
    .clk_2_N_out(clk_2_wires[108]),
    .clk_2_E_in(clk_2_wires[107]),
    .prog_clk_2_N_out(prog_clk_2_wires[108]),
    .prog_clk_2_E_in(prog_clk_2_wires[107]),
    .prog_clk_0_N_in(prog_clk_0_wires[285]),
    .pReset_E_out(pResetWires[531]),
    .pReset_N_out(pResetWires[530]),
    .pReset_W_in(pResetWires[528]),
    .chany_top_in(cby_1__1__82_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_82_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_82_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_82_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_82_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_82_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_82_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_82_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_82_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__86_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_93_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_93_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_93_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_93_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_93_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_93_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_93_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_93_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__81_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_81_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_81_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_81_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_81_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_81_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_81_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_81_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_81_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__75_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_81_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_81_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_81_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_81_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_81_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_81_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_81_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_81_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__86_ccff_tail[0]),
    .chany_top_out(sb_1__1__75_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__75_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__75_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__75_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__75_ccff_tail[0])
  );


  sb_1__1_
  sb_7__11_
  (
    .clk_1_S_in(clk_2_wires[109]),
    .clk_1_W_out(clk_1_wires[163]),
    .clk_1_E_out(clk_1_wires[162]),
    .prog_clk_1_S_in(prog_clk_2_wires[109]),
    .prog_clk_1_W_out(prog_clk_1_wires[163]),
    .prog_clk_1_E_out(prog_clk_1_wires[162]),
    .prog_clk_0_N_in(prog_clk_0_wires[288]),
    .pReset_E_out(pResetWires[580]),
    .pReset_N_out(pResetWires[579]),
    .pReset_W_in(pResetWires[577]),
    .chany_top_in(cby_1__1__83_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_83_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_83_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_83_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_83_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_83_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_83_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_83_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_83_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__87_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_94_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_94_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_94_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_94_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_94_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_94_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_94_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_94_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__82_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_82_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_82_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_82_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_82_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_82_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_82_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_82_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_82_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__76_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_82_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_82_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_82_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_82_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_82_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_82_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_82_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_82_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__87_ccff_tail[0]),
    .chany_top_out(sb_1__1__76_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__76_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__76_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__76_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__76_ccff_tail[0])
  );


  sb_1__1_
  sb_8__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[296]),
    .pReset_E_out(pResetWires[94]),
    .pReset_N_out(pResetWires[93]),
    .pReset_W_in(pResetWires[91]),
    .chany_top_in(cby_1__1__85_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_85_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_85_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_85_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_85_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_85_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_85_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_85_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_85_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__88_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_96_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_96_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_96_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_96_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_96_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_96_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_96_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_96_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__84_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_84_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_84_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_84_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_84_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_84_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_84_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_84_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_84_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__77_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_84_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_84_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_84_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_84_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_84_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_84_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_84_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_84_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__88_ccff_tail[0]),
    .chany_top_out(sb_1__1__77_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__77_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__77_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__77_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__77_ccff_tail[0])
  );


  sb_1__1_
  sb_8__2_
  (
    .clk_2_N_in(clk_3_wires[43]),
    .clk_2_W_out(clk_2_wires[71]),
    .clk_2_E_out(clk_2_wires[69]),
    .prog_clk_2_N_in(prog_clk_3_wires[43]),
    .prog_clk_2_W_out(prog_clk_2_wires[71]),
    .prog_clk_2_E_out(prog_clk_2_wires[69]),
    .prog_clk_0_N_in(prog_clk_0_wires[299]),
    .pReset_E_out(pResetWires[143]),
    .pReset_N_out(pResetWires[142]),
    .pReset_W_in(pResetWires[140]),
    .chany_top_in(cby_1__1__86_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_86_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_86_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_86_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_86_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_86_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_86_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_86_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_86_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__89_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_97_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_97_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_97_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_97_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_97_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_97_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_97_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_97_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__85_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_85_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_85_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_85_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_85_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_85_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_85_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_85_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_85_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__78_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_85_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_85_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_85_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_85_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_85_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_85_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_85_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_85_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__89_ccff_tail[0]),
    .chany_top_out(sb_1__1__78_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__78_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__78_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__78_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__78_ccff_tail[0])
  );


  sb_1__1_
  sb_8__3_
  (
    .clk_3_S_out(clk_3_wires[42]),
    .clk_3_N_in(clk_3_wires[39]),
    .prog_clk_3_S_out(prog_clk_3_wires[42]),
    .prog_clk_3_N_in(prog_clk_3_wires[39]),
    .prog_clk_0_N_in(prog_clk_0_wires[302]),
    .pReset_E_out(pResetWires[192]),
    .pReset_N_out(pResetWires[191]),
    .pReset_W_in(pResetWires[189]),
    .chany_top_in(cby_1__1__87_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_87_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_87_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_87_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_87_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_87_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_87_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_87_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_87_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__90_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_98_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_98_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_98_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_98_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_98_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_98_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_98_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_98_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__86_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_86_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_86_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_86_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_86_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_86_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_86_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_86_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_86_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__79_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_86_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_86_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_86_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_86_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_86_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_86_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_86_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_86_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__90_ccff_tail[0]),
    .chany_top_out(sb_1__1__79_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__79_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__79_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__79_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__79_ccff_tail[0])
  );


  sb_1__1_
  sb_8__4_
  (
    .clk_3_S_out(clk_3_wires[38]),
    .clk_2_N_in(clk_3_wires[33]),
    .clk_3_N_in(clk_3_wires[33]),
    .clk_2_W_out(clk_2_wires[80]),
    .clk_2_E_out(clk_2_wires[78]),
    .prog_clk_3_S_out(prog_clk_3_wires[38]),
    .prog_clk_2_N_in(prog_clk_3_wires[33]),
    .prog_clk_3_N_in(prog_clk_3_wires[33]),
    .prog_clk_2_W_out(prog_clk_2_wires[80]),
    .prog_clk_2_E_out(prog_clk_2_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[305]),
    .pReset_E_out(pResetWires[241]),
    .pReset_N_out(pResetWires[240]),
    .pReset_W_in(pResetWires[238]),
    .chany_top_in(cby_1__1__88_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_88_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_88_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_88_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_88_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_88_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_88_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_88_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_88_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__91_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_99_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_99_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_99_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_99_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_99_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_99_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_99_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_99_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__87_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_87_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_87_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_87_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_87_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_87_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_87_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_87_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_87_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__80_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_87_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_87_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_87_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_87_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_87_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_87_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_87_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_87_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__91_ccff_tail[0]),
    .chany_top_out(sb_1__1__80_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__80_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__80_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__80_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__80_ccff_tail[0])
  );


  sb_1__1_
  sb_8__5_
  (
    .clk_3_S_out(clk_3_wires[32]),
    .clk_3_N_in(clk_3_wires[29]),
    .prog_clk_3_S_out(prog_clk_3_wires[32]),
    .prog_clk_3_N_in(prog_clk_3_wires[29]),
    .prog_clk_0_N_in(prog_clk_0_wires[308]),
    .pReset_E_out(pResetWires[290]),
    .pReset_N_out(pResetWires[289]),
    .pReset_W_in(pResetWires[287]),
    .chany_top_in(cby_1__1__89_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_89_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_89_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_89_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_89_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_89_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_89_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_89_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_89_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__92_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_100_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_100_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_100_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_100_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_100_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_100_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_100_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_100_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__88_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_88_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_88_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_88_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_88_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_88_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_88_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_88_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_88_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__81_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_88_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_88_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_88_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_88_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_88_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_88_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_88_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_88_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__92_ccff_tail[0]),
    .chany_top_out(sb_1__1__81_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__81_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__81_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__81_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__81_ccff_tail[0])
  );


  sb_1__1_
  sb_8__6_
  (
    .clk_3_E_out(clk_3_wires[44]),
    .clk_3_S_out(clk_3_wires[28]),
    .clk_3_N_out(clk_3_wires[26]),
    .clk_3_W_in(clk_3_wires[5]),
    .prog_clk_3_E_out(prog_clk_3_wires[44]),
    .prog_clk_3_S_out(prog_clk_3_wires[28]),
    .prog_clk_3_N_out(prog_clk_3_wires[26]),
    .prog_clk_3_W_in(prog_clk_3_wires[5]),
    .prog_clk_0_N_in(prog_clk_0_wires[311]),
    .pReset_E_out(pResetWires[339]),
    .pReset_N_out(pResetWires[338]),
    .pReset_W_in(pResetWires[336]),
    .chany_top_in(cby_1__1__90_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_90_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_90_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_90_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_90_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_90_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_90_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_90_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_90_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__93_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_101_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_101_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_101_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_101_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_101_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_101_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_101_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_101_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__89_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_89_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_89_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_89_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_89_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_89_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_89_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_89_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_89_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__82_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_89_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_89_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_89_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_89_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_89_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_89_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_89_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_89_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__93_ccff_tail[0]),
    .chany_top_out(sb_1__1__82_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__82_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__82_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__82_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__82_ccff_tail[0])
  );


  sb_1__1_
  sb_8__7_
  (
    .clk_3_N_out(clk_3_wires[30]),
    .clk_3_S_in(clk_3_wires[27]),
    .prog_clk_3_N_out(prog_clk_3_wires[30]),
    .prog_clk_3_S_in(prog_clk_3_wires[27]),
    .prog_clk_0_N_in(prog_clk_0_wires[314]),
    .pReset_E_out(pResetWires[388]),
    .pReset_N_out(pResetWires[387]),
    .pReset_W_in(pResetWires[385]),
    .chany_top_in(cby_1__1__91_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_91_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_91_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_91_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_91_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_91_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_91_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_91_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_91_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__94_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_102_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_102_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_102_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_102_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_102_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_102_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_102_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_102_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__90_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_90_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_90_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_90_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_90_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_90_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_90_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_90_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_90_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__83_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_90_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_90_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_90_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_90_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_90_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_90_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_90_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_90_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__94_ccff_tail[0]),
    .chany_top_out(sb_1__1__83_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__83_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__83_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__83_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__83_ccff_tail[0])
  );


  sb_1__1_
  sb_8__8_
  (
    .clk_3_N_out(clk_3_wires[36]),
    .clk_2_S_in(clk_3_wires[31]),
    .clk_3_S_in(clk_3_wires[31]),
    .clk_2_W_out(clk_2_wires[93]),
    .clk_2_E_out(clk_2_wires[91]),
    .prog_clk_3_N_out(prog_clk_3_wires[36]),
    .prog_clk_2_S_in(prog_clk_3_wires[31]),
    .prog_clk_3_S_in(prog_clk_3_wires[31]),
    .prog_clk_2_W_out(prog_clk_2_wires[93]),
    .prog_clk_2_E_out(prog_clk_2_wires[91]),
    .prog_clk_0_N_in(prog_clk_0_wires[317]),
    .pReset_E_out(pResetWires[437]),
    .pReset_N_out(pResetWires[436]),
    .pReset_W_in(pResetWires[434]),
    .chany_top_in(cby_1__1__92_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_92_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_92_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_92_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_92_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_92_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_92_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_92_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_92_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__95_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_103_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_103_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_103_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_103_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_103_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_103_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_103_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_103_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__91_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_91_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_91_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_91_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_91_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_91_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_91_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_91_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_91_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__84_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_91_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_91_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_91_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_91_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_91_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_91_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_91_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_91_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__95_ccff_tail[0]),
    .chany_top_out(sb_1__1__84_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__84_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__84_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__84_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__84_ccff_tail[0])
  );


  sb_1__1_
  sb_8__9_
  (
    .clk_3_N_out(clk_3_wires[40]),
    .clk_3_S_in(clk_3_wires[37]),
    .prog_clk_3_N_out(prog_clk_3_wires[40]),
    .prog_clk_3_S_in(prog_clk_3_wires[37]),
    .prog_clk_0_N_in(prog_clk_0_wires[320]),
    .pReset_E_out(pResetWires[486]),
    .pReset_N_out(pResetWires[485]),
    .pReset_W_in(pResetWires[483]),
    .chany_top_in(cby_1__1__93_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_93_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_93_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_93_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_93_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_93_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_93_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_93_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_93_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__96_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_104_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_104_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_104_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_104_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_104_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_104_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_104_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_104_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__92_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_92_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_92_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_92_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_92_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_92_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_92_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_92_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_92_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__85_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_92_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_92_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_92_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_92_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_92_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_92_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_92_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_92_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__96_ccff_tail[0]),
    .chany_top_out(sb_1__1__85_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__85_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__85_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__85_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__85_ccff_tail[0])
  );


  sb_1__1_
  sb_8__10_
  (
    .clk_2_S_in(clk_3_wires[41]),
    .clk_2_W_out(clk_2_wires[106]),
    .clk_2_E_out(clk_2_wires[104]),
    .prog_clk_2_S_in(prog_clk_3_wires[41]),
    .prog_clk_2_W_out(prog_clk_2_wires[106]),
    .prog_clk_2_E_out(prog_clk_2_wires[104]),
    .prog_clk_0_N_in(prog_clk_0_wires[323]),
    .pReset_E_out(pResetWires[535]),
    .pReset_N_out(pResetWires[534]),
    .pReset_W_in(pResetWires[532]),
    .chany_top_in(cby_1__1__94_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_94_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_94_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_94_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_94_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_94_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_94_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_94_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_94_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__97_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_105_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_105_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_105_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_105_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_105_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_105_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_105_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_105_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__93_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_93_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_93_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_93_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_93_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_93_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_93_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_93_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_93_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__86_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_93_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_93_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_93_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_93_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_93_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_93_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_93_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_93_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__97_ccff_tail[0]),
    .chany_top_out(sb_1__1__86_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__86_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__86_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__86_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__86_ccff_tail[0])
  );


  sb_1__1_
  sb_8__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[326]),
    .pReset_E_out(pResetWires[584]),
    .pReset_N_out(pResetWires[583]),
    .pReset_W_in(pResetWires[581]),
    .chany_top_in(cby_1__1__95_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_95_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_95_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_95_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_95_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_95_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_95_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_95_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_95_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__98_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_106_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_106_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_106_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_106_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_106_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_106_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_106_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_106_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__94_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_94_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_94_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_94_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_94_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_94_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_94_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_94_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_94_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__87_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_94_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_94_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_94_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_94_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_94_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_94_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_94_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_94_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__98_ccff_tail[0]),
    .chany_top_out(sb_1__1__87_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__87_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__87_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__87_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__87_ccff_tail[0])
  );


  sb_1__1_
  sb_9__1_
  (
    .clk_1_N_in(clk_2_wires[76]),
    .clk_1_W_out(clk_1_wires[170]),
    .clk_1_E_out(clk_1_wires[169]),
    .prog_clk_1_N_in(prog_clk_2_wires[76]),
    .prog_clk_1_W_out(prog_clk_1_wires[170]),
    .prog_clk_1_E_out(prog_clk_1_wires[169]),
    .prog_clk_0_N_in(prog_clk_0_wires[334]),
    .pReset_E_out(pResetWires[98]),
    .pReset_N_out(pResetWires[97]),
    .pReset_W_in(pResetWires[95]),
    .chany_top_in(cby_1__1__97_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_97_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_97_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_97_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_97_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_97_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_97_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_97_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_97_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__99_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_108_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_108_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_108_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_108_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_108_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_108_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_108_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_108_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__96_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_96_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_96_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_96_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_96_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_96_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_96_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_96_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_96_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__88_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_96_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_96_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_96_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_96_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_96_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_96_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_96_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_96_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__99_ccff_tail[0]),
    .chany_top_out(sb_1__1__88_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__88_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__88_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__88_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__88_ccff_tail[0])
  );


  sb_1__1_
  sb_9__2_
  (
    .clk_2_S_out(clk_2_wires[75]),
    .clk_2_W_in(clk_2_wires[70]),
    .prog_clk_2_S_out(prog_clk_2_wires[75]),
    .prog_clk_2_W_in(prog_clk_2_wires[70]),
    .prog_clk_0_N_in(prog_clk_0_wires[337]),
    .pReset_E_out(pResetWires[147]),
    .pReset_N_out(pResetWires[146]),
    .pReset_W_in(pResetWires[144]),
    .chany_top_in(cby_1__1__98_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_98_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_98_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_98_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_98_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_98_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_98_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_98_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_98_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__100_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_109_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_109_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_109_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_109_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_109_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_109_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_109_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_109_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__97_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_97_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_97_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_97_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_97_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_97_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_97_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_97_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_97_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__89_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_97_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_97_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_97_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_97_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_97_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_97_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_97_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_97_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__100_ccff_tail[0]),
    .chany_top_out(sb_1__1__89_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__89_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__89_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__89_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__89_ccff_tail[0])
  );


  sb_1__1_
  sb_9__3_
  (
    .clk_1_N_in(clk_2_wires[89]),
    .clk_1_W_out(clk_1_wires[177]),
    .clk_1_E_out(clk_1_wires[176]),
    .prog_clk_1_N_in(prog_clk_2_wires[89]),
    .prog_clk_1_W_out(prog_clk_1_wires[177]),
    .prog_clk_1_E_out(prog_clk_1_wires[176]),
    .prog_clk_0_N_in(prog_clk_0_wires[340]),
    .pReset_E_out(pResetWires[196]),
    .pReset_N_out(pResetWires[195]),
    .pReset_W_in(pResetWires[193]),
    .chany_top_in(cby_1__1__99_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_99_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_99_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_99_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_99_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_99_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_99_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_99_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_99_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__101_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_110_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_110_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_110_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_110_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_110_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_110_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_110_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_110_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__98_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_98_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_98_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_98_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_98_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_98_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_98_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_98_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_98_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__90_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_98_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_98_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_98_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_98_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_98_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_98_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_98_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_98_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__101_ccff_tail[0]),
    .chany_top_out(sb_1__1__90_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__90_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__90_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__90_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__90_ccff_tail[0])
  );


  sb_1__1_
  sb_9__4_
  (
    .clk_2_S_out(clk_2_wires[88]),
    .clk_2_N_out(clk_2_wires[86]),
    .clk_2_W_in(clk_2_wires[79]),
    .prog_clk_2_S_out(prog_clk_2_wires[88]),
    .prog_clk_2_N_out(prog_clk_2_wires[86]),
    .prog_clk_2_W_in(prog_clk_2_wires[79]),
    .prog_clk_0_N_in(prog_clk_0_wires[343]),
    .pReset_E_out(pResetWires[245]),
    .pReset_N_out(pResetWires[244]),
    .pReset_W_in(pResetWires[242]),
    .chany_top_in(cby_1__1__100_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_100_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_100_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_100_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_100_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_100_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_100_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_100_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_100_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__102_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_111_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_111_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_111_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_111_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_111_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_111_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_111_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_111_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__99_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_99_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_99_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_99_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_99_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_99_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_99_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_99_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_99_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__91_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_99_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_99_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_99_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_99_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_99_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_99_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_99_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_99_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__102_ccff_tail[0]),
    .chany_top_out(sb_1__1__91_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__91_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__91_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__91_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__91_ccff_tail[0])
  );


  sb_1__1_
  sb_9__5_
  (
    .clk_1_S_in(clk_2_wires[87]),
    .clk_1_W_out(clk_1_wires[184]),
    .clk_1_E_out(clk_1_wires[183]),
    .prog_clk_1_S_in(prog_clk_2_wires[87]),
    .prog_clk_1_W_out(prog_clk_1_wires[184]),
    .prog_clk_1_E_out(prog_clk_1_wires[183]),
    .prog_clk_0_N_in(prog_clk_0_wires[346]),
    .pReset_E_out(pResetWires[294]),
    .pReset_N_out(pResetWires[293]),
    .pReset_W_in(pResetWires[291]),
    .chany_top_in(cby_1__1__101_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_101_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_101_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_101_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_101_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_101_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_101_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_101_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_101_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__103_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_112_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_112_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_112_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_112_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_112_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_112_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_112_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_112_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__100_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_100_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_100_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_100_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_100_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_100_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_100_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_100_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_100_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__92_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_100_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_100_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_100_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_100_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_100_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_100_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_100_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_100_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__103_ccff_tail[0]),
    .chany_top_out(sb_1__1__92_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__92_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__92_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__92_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__92_ccff_tail[0])
  );


  sb_1__1_
  sb_9__6_
  (
    .clk_3_E_out(clk_3_wires[48]),
    .clk_3_W_in(clk_3_wires[45]),
    .prog_clk_3_E_out(prog_clk_3_wires[48]),
    .prog_clk_3_W_in(prog_clk_3_wires[45]),
    .prog_clk_0_N_in(prog_clk_0_wires[349]),
    .pReset_E_out(pResetWires[343]),
    .pReset_N_out(pResetWires[342]),
    .pReset_W_in(pResetWires[340]),
    .chany_top_in(cby_1__1__102_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_102_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_102_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_102_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_102_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_102_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_102_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_102_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_102_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__104_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_113_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_113_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_113_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_113_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_113_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_113_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_113_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_113_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__101_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_101_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_101_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_101_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_101_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_101_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_101_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_101_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_101_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__93_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_101_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_101_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_101_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_101_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_101_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_101_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_101_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_101_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__104_ccff_tail[0]),
    .chany_top_out(sb_1__1__93_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__93_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__93_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__93_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__93_ccff_tail[0])
  );


  sb_1__1_
  sb_9__7_
  (
    .clk_1_N_in(clk_2_wires[102]),
    .clk_1_W_out(clk_1_wires[191]),
    .clk_1_E_out(clk_1_wires[190]),
    .prog_clk_1_N_in(prog_clk_2_wires[102]),
    .prog_clk_1_W_out(prog_clk_1_wires[191]),
    .prog_clk_1_E_out(prog_clk_1_wires[190]),
    .prog_clk_0_N_in(prog_clk_0_wires[352]),
    .pReset_E_out(pResetWires[392]),
    .pReset_N_out(pResetWires[391]),
    .pReset_W_in(pResetWires[389]),
    .chany_top_in(cby_1__1__103_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_103_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_103_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_103_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_103_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_103_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_103_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_103_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_103_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__105_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_114_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_114_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_114_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_114_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_114_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_114_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_114_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_114_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__102_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_102_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_102_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_102_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_102_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_102_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_102_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_102_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_102_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__94_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_102_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_102_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_102_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_102_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_102_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_102_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_102_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_102_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__105_ccff_tail[0]),
    .chany_top_out(sb_1__1__94_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__94_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__94_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__94_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__94_ccff_tail[0])
  );


  sb_1__1_
  sb_9__8_
  (
    .clk_2_S_out(clk_2_wires[101]),
    .clk_2_N_out(clk_2_wires[99]),
    .clk_2_W_in(clk_2_wires[92]),
    .prog_clk_2_S_out(prog_clk_2_wires[101]),
    .prog_clk_2_N_out(prog_clk_2_wires[99]),
    .prog_clk_2_W_in(prog_clk_2_wires[92]),
    .prog_clk_0_N_in(prog_clk_0_wires[355]),
    .pReset_E_out(pResetWires[441]),
    .pReset_N_out(pResetWires[440]),
    .pReset_W_in(pResetWires[438]),
    .chany_top_in(cby_1__1__104_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_104_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_104_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_104_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_104_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_104_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_104_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_104_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_104_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__106_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_115_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_115_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_115_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_115_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_115_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_115_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_115_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_115_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__103_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_103_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_103_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_103_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_103_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_103_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_103_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_103_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_103_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__95_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_103_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_103_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_103_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_103_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_103_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_103_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_103_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_103_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__106_ccff_tail[0]),
    .chany_top_out(sb_1__1__95_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__95_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__95_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__95_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__95_ccff_tail[0])
  );


  sb_1__1_
  sb_9__9_
  (
    .clk_1_S_in(clk_2_wires[100]),
    .clk_1_W_out(clk_1_wires[198]),
    .clk_1_E_out(clk_1_wires[197]),
    .prog_clk_1_S_in(prog_clk_2_wires[100]),
    .prog_clk_1_W_out(prog_clk_1_wires[198]),
    .prog_clk_1_E_out(prog_clk_1_wires[197]),
    .prog_clk_0_N_in(prog_clk_0_wires[358]),
    .pReset_E_out(pResetWires[490]),
    .pReset_N_out(pResetWires[489]),
    .pReset_W_in(pResetWires[487]),
    .chany_top_in(cby_1__1__105_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_105_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_105_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_105_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_105_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_105_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_105_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_105_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_105_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__107_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_116_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_116_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_116_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_116_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_116_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_116_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_116_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_116_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__104_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_104_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_104_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_104_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_104_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_104_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_104_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_104_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_104_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__96_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_104_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_104_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_104_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_104_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_104_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_104_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_104_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_104_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__107_ccff_tail[0]),
    .chany_top_out(sb_1__1__96_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__96_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__96_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__96_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__96_ccff_tail[0])
  );


  sb_1__1_
  sb_9__10_
  (
    .clk_2_N_out(clk_2_wires[110]),
    .clk_2_W_in(clk_2_wires[105]),
    .prog_clk_2_N_out(prog_clk_2_wires[110]),
    .prog_clk_2_W_in(prog_clk_2_wires[105]),
    .prog_clk_0_N_in(prog_clk_0_wires[361]),
    .pReset_E_out(pResetWires[539]),
    .pReset_N_out(pResetWires[538]),
    .pReset_W_in(pResetWires[536]),
    .chany_top_in(cby_1__1__106_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_106_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_106_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_106_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_106_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_106_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_106_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_106_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_106_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__108_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_117_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_117_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_117_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_117_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_117_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_117_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_117_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_117_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__105_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_105_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_105_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_105_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_105_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_105_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_105_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_105_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_105_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__97_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_105_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_105_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_105_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_105_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_105_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_105_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_105_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_105_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__108_ccff_tail[0]),
    .chany_top_out(sb_1__1__97_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__97_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__97_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__97_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__97_ccff_tail[0])
  );


  sb_1__1_
  sb_9__11_
  (
    .clk_1_S_in(clk_2_wires[111]),
    .clk_1_W_out(clk_1_wires[205]),
    .clk_1_E_out(clk_1_wires[204]),
    .prog_clk_1_S_in(prog_clk_2_wires[111]),
    .prog_clk_1_W_out(prog_clk_1_wires[205]),
    .prog_clk_1_E_out(prog_clk_1_wires[204]),
    .prog_clk_0_N_in(prog_clk_0_wires[364]),
    .pReset_E_out(pResetWires[588]),
    .pReset_N_out(pResetWires[587]),
    .pReset_W_in(pResetWires[585]),
    .chany_top_in(cby_1__1__107_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_107_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_107_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_107_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_107_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_107_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_107_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_107_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_107_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__109_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_118_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_118_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_118_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_118_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_118_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_118_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_118_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_118_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__106_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_106_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_106_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_106_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_106_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_106_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_106_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_106_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_106_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__98_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_106_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_106_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_106_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_106_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_106_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_106_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_106_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_106_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__109_ccff_tail[0]),
    .chany_top_out(sb_1__1__98_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__98_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__98_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__98_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__98_ccff_tail[0])
  );


  sb_1__1_
  sb_10__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[372]),
    .pReset_E_out(pResetWires[102]),
    .pReset_N_out(pResetWires[101]),
    .pReset_W_in(pResetWires[99]),
    .chany_top_in(cby_1__1__109_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_109_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_109_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_109_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_109_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_109_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_109_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_109_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_109_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__110_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_120_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_120_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_120_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_120_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_120_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_120_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_120_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_120_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__108_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_108_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_108_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_108_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_108_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_108_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_108_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_108_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_108_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__99_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_108_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_108_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_108_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_108_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_108_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_108_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_108_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_108_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__110_ccff_tail[0]),
    .chany_top_out(sb_1__1__99_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__99_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__99_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__99_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__99_ccff_tail[0])
  );


  sb_1__1_
  sb_10__2_
  (
    .clk_2_N_in(clk_3_wires[87]),
    .clk_2_E_out(clk_2_wires[114]),
    .prog_clk_2_N_in(prog_clk_3_wires[87]),
    .prog_clk_2_E_out(prog_clk_2_wires[114]),
    .prog_clk_0_N_in(prog_clk_0_wires[375]),
    .pReset_E_out(pResetWires[151]),
    .pReset_N_out(pResetWires[150]),
    .pReset_W_in(pResetWires[148]),
    .chany_top_in(cby_1__1__110_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_110_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_110_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_110_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_110_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_110_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_110_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_110_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_110_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__111_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_121_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_121_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_121_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_121_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_121_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_121_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_121_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_121_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__109_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_109_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_109_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_109_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_109_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_109_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_109_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_109_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_109_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__100_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_109_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_109_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_109_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_109_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_109_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_109_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_109_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_109_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__111_ccff_tail[0]),
    .chany_top_out(sb_1__1__100_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__100_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__100_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__100_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__100_ccff_tail[0])
  );


  sb_1__1_
  sb_10__3_
  (
    .clk_3_S_out(clk_3_wires[86]),
    .clk_3_N_in(clk_3_wires[83]),
    .prog_clk_3_S_out(prog_clk_3_wires[86]),
    .prog_clk_3_N_in(prog_clk_3_wires[83]),
    .prog_clk_0_N_in(prog_clk_0_wires[378]),
    .pReset_E_out(pResetWires[200]),
    .pReset_N_out(pResetWires[199]),
    .pReset_W_in(pResetWires[197]),
    .chany_top_in(cby_1__1__111_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_111_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_111_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_111_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_111_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_111_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_111_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_111_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_111_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__112_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_122_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_122_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_122_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_122_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_122_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_122_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_122_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_122_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__110_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_110_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_110_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_110_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_110_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_110_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_110_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_110_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_110_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__101_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_110_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_110_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_110_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_110_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_110_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_110_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_110_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_110_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__112_ccff_tail[0]),
    .chany_top_out(sb_1__1__101_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__101_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__101_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__101_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__101_ccff_tail[0])
  );


  sb_1__1_
  sb_10__4_
  (
    .clk_3_S_out(clk_3_wires[82]),
    .clk_2_N_in(clk_3_wires[77]),
    .clk_3_N_in(clk_3_wires[77]),
    .clk_2_E_out(clk_2_wires[119]),
    .prog_clk_3_S_out(prog_clk_3_wires[82]),
    .prog_clk_2_N_in(prog_clk_3_wires[77]),
    .prog_clk_3_N_in(prog_clk_3_wires[77]),
    .prog_clk_2_E_out(prog_clk_2_wires[119]),
    .prog_clk_0_N_in(prog_clk_0_wires[381]),
    .pReset_E_out(pResetWires[249]),
    .pReset_N_out(pResetWires[248]),
    .pReset_W_in(pResetWires[246]),
    .chany_top_in(cby_1__1__112_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_112_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_112_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_112_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_112_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_112_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_112_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_112_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_112_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__113_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_123_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_123_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_123_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_123_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_123_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_123_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_123_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_123_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__111_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_111_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_111_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_111_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_111_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_111_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_111_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_111_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_111_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__102_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_111_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_111_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_111_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_111_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_111_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_111_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_111_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_111_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__113_ccff_tail[0]),
    .chany_top_out(sb_1__1__102_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__102_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__102_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__102_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__102_ccff_tail[0])
  );


  sb_1__1_
  sb_10__5_
  (
    .clk_3_S_out(clk_3_wires[76]),
    .clk_3_N_in(clk_3_wires[73]),
    .prog_clk_3_S_out(prog_clk_3_wires[76]),
    .prog_clk_3_N_in(prog_clk_3_wires[73]),
    .prog_clk_0_N_in(prog_clk_0_wires[384]),
    .pReset_E_out(pResetWires[298]),
    .pReset_N_out(pResetWires[297]),
    .pReset_W_in(pResetWires[295]),
    .chany_top_in(cby_1__1__113_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_113_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_113_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_113_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_113_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_113_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_113_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_113_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_113_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__114_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_124_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_124_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_124_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_124_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_124_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_124_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_124_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_124_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__112_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_112_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_112_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_112_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_112_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_112_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_112_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_112_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_112_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__103_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_112_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_112_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_112_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_112_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_112_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_112_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_112_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_112_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__114_ccff_tail[0]),
    .chany_top_out(sb_1__1__103_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__103_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__103_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__103_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__103_ccff_tail[0])
  );


  sb_1__1_
  sb_10__6_
  (
    .clk_3_S_out(clk_3_wires[72]),
    .clk_3_N_out(clk_3_wires[70]),
    .clk_3_W_in(clk_3_wires[49]),
    .prog_clk_3_S_out(prog_clk_3_wires[72]),
    .prog_clk_3_N_out(prog_clk_3_wires[70]),
    .prog_clk_3_W_in(prog_clk_3_wires[49]),
    .prog_clk_0_N_in(prog_clk_0_wires[387]),
    .pReset_E_out(pResetWires[347]),
    .pReset_N_out(pResetWires[346]),
    .pReset_W_in(pResetWires[344]),
    .chany_top_in(cby_1__1__114_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_114_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_114_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_114_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_114_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_114_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_114_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_114_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_114_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__115_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_125_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_125_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_125_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_125_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_125_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_125_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_125_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_125_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__113_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_113_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_113_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_113_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_113_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_113_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_113_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_113_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_113_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__104_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_113_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_113_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_113_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_113_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_113_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_113_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_113_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_113_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__115_ccff_tail[0]),
    .chany_top_out(sb_1__1__104_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__104_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__104_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__104_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__104_ccff_tail[0])
  );


  sb_1__1_
  sb_10__7_
  (
    .clk_3_N_out(clk_3_wires[74]),
    .clk_3_S_in(clk_3_wires[71]),
    .prog_clk_3_N_out(prog_clk_3_wires[74]),
    .prog_clk_3_S_in(prog_clk_3_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[390]),
    .pReset_E_out(pResetWires[396]),
    .pReset_N_out(pResetWires[395]),
    .pReset_W_in(pResetWires[393]),
    .chany_top_in(cby_1__1__115_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_115_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_115_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_115_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_115_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_115_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_115_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_115_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_115_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__116_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_126_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_126_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_126_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_126_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_126_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_126_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_126_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_126_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__114_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_114_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_114_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_114_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_114_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_114_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_114_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_114_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_114_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__105_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_114_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_114_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_114_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_114_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_114_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_114_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_114_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_114_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__116_ccff_tail[0]),
    .chany_top_out(sb_1__1__105_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__105_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__105_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__105_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__105_ccff_tail[0])
  );


  sb_1__1_
  sb_10__8_
  (
    .clk_3_N_out(clk_3_wires[80]),
    .clk_2_S_in(clk_3_wires[75]),
    .clk_3_S_in(clk_3_wires[75]),
    .clk_2_E_out(clk_2_wires[126]),
    .prog_clk_3_N_out(prog_clk_3_wires[80]),
    .prog_clk_2_S_in(prog_clk_3_wires[75]),
    .prog_clk_3_S_in(prog_clk_3_wires[75]),
    .prog_clk_2_E_out(prog_clk_2_wires[126]),
    .prog_clk_0_N_in(prog_clk_0_wires[393]),
    .pReset_E_out(pResetWires[445]),
    .pReset_N_out(pResetWires[444]),
    .pReset_W_in(pResetWires[442]),
    .chany_top_in(cby_1__1__116_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_116_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_116_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_116_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_116_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_116_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_116_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_116_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_116_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__117_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_127_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_127_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_127_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_127_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_127_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_127_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_127_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_127_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__115_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_115_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_115_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_115_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_115_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_115_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_115_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_115_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_115_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__106_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_115_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_115_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_115_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_115_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_115_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_115_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_115_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_115_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__117_ccff_tail[0]),
    .chany_top_out(sb_1__1__106_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__106_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__106_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__106_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__106_ccff_tail[0])
  );


  sb_1__1_
  sb_10__9_
  (
    .clk_3_N_out(clk_3_wires[84]),
    .clk_3_S_in(clk_3_wires[81]),
    .prog_clk_3_N_out(prog_clk_3_wires[84]),
    .prog_clk_3_S_in(prog_clk_3_wires[81]),
    .prog_clk_0_N_in(prog_clk_0_wires[396]),
    .pReset_E_out(pResetWires[494]),
    .pReset_N_out(pResetWires[493]),
    .pReset_W_in(pResetWires[491]),
    .chany_top_in(cby_1__1__117_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_117_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_117_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_117_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_117_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_117_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_117_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_117_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_117_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__118_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_128_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_128_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_128_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_128_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_128_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_128_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_128_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_128_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__116_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_116_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_116_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_116_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_116_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_116_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_116_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_116_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_116_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__107_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_116_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_116_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_116_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_116_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_116_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_116_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_116_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_116_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__118_ccff_tail[0]),
    .chany_top_out(sb_1__1__107_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__107_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__107_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__107_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__107_ccff_tail[0])
  );


  sb_1__1_
  sb_10__10_
  (
    .clk_2_S_in(clk_3_wires[85]),
    .clk_2_E_out(clk_2_wires[133]),
    .prog_clk_2_S_in(prog_clk_3_wires[85]),
    .prog_clk_2_E_out(prog_clk_2_wires[133]),
    .prog_clk_0_N_in(prog_clk_0_wires[399]),
    .pReset_E_out(pResetWires[543]),
    .pReset_N_out(pResetWires[542]),
    .pReset_W_in(pResetWires[540]),
    .chany_top_in(cby_1__1__118_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_118_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_118_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_118_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_118_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_118_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_118_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_118_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_118_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__119_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_129_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_129_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_129_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_129_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_129_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_129_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_129_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_129_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__117_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_117_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_117_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_117_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_117_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_117_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_117_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_117_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_117_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__108_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_117_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_117_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_117_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_117_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_117_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_117_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_117_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_117_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__119_ccff_tail[0]),
    .chany_top_out(sb_1__1__108_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__108_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__108_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__108_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__108_ccff_tail[0])
  );


  sb_1__1_
  sb_10__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[402]),
    .pReset_E_out(pResetWires[592]),
    .pReset_N_out(pResetWires[591]),
    .pReset_W_in(pResetWires[589]),
    .chany_top_in(cby_1__1__119_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_119_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_119_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_119_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_119_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_119_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_119_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_119_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_119_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__120_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_130_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_130_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_130_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_130_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_130_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_130_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_130_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_130_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__118_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_118_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_118_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_118_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_118_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_118_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_118_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_118_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_118_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__109_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_118_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_118_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_118_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_118_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_118_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_118_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_118_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_118_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__120_ccff_tail[0]),
    .chany_top_out(sb_1__1__109_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__109_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__109_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__109_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__109_ccff_tail[0])
  );


  sb_1__1_
  sb_11__1_
  (
    .clk_1_N_in(clk_2_wires[116]),
    .clk_1_W_out(clk_1_wires[212]),
    .clk_1_E_out(clk_1_wires[211]),
    .prog_clk_1_N_in(prog_clk_2_wires[116]),
    .prog_clk_1_W_out(prog_clk_1_wires[212]),
    .prog_clk_1_E_out(prog_clk_1_wires[211]),
    .prog_clk_0_N_in(prog_clk_0_wires[410]),
    .pReset_E_out(pResetWires[106]),
    .pReset_N_out(pResetWires[105]),
    .pReset_W_in(pResetWires[103]),
    .chany_top_in(cby_1__1__121_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_121_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_121_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_121_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_121_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_121_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_121_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_121_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_121_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__121_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_132_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_132_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_132_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_132_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_132_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_132_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_132_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_132_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__120_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_120_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_120_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_120_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_120_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_120_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_120_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_120_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_120_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__110_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_120_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_120_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_120_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_120_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_120_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_120_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_120_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_120_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__121_ccff_tail[0]),
    .chany_top_out(sb_1__1__110_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__110_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__110_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__110_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__110_ccff_tail[0])
  );


  sb_1__1_
  sb_11__2_
  (
    .clk_2_S_out(clk_2_wires[115]),
    .clk_2_W_in(clk_2_wires[113]),
    .prog_clk_2_S_out(prog_clk_2_wires[115]),
    .prog_clk_2_W_in(prog_clk_2_wires[113]),
    .prog_clk_0_N_in(prog_clk_0_wires[413]),
    .pReset_E_out(pResetWires[155]),
    .pReset_N_out(pResetWires[154]),
    .pReset_W_in(pResetWires[152]),
    .chany_top_in(cby_1__1__122_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_122_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_122_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_122_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_122_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_122_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_122_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_122_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_122_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__122_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_133_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_133_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_133_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_133_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_133_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_133_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_133_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_133_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__121_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_121_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_121_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_121_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_121_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_121_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_121_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_121_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_121_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__111_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_121_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_121_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_121_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_121_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_121_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_121_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_121_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_121_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__122_ccff_tail[0]),
    .chany_top_out(sb_1__1__111_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__111_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__111_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__111_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__111_ccff_tail[0])
  );


  sb_1__1_
  sb_11__3_
  (
    .clk_1_N_in(clk_2_wires[123]),
    .clk_1_W_out(clk_1_wires[219]),
    .clk_1_E_out(clk_1_wires[218]),
    .prog_clk_1_N_in(prog_clk_2_wires[123]),
    .prog_clk_1_W_out(prog_clk_1_wires[219]),
    .prog_clk_1_E_out(prog_clk_1_wires[218]),
    .prog_clk_0_N_in(prog_clk_0_wires[416]),
    .pReset_E_out(pResetWires[204]),
    .pReset_N_out(pResetWires[203]),
    .pReset_W_in(pResetWires[201]),
    .chany_top_in(cby_1__1__123_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_123_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_123_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_123_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_123_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_123_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_123_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_123_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_123_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__123_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_134_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_134_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_134_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_134_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_134_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_134_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_134_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_134_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__122_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_122_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_122_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_122_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_122_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_122_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_122_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_122_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_122_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__112_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_122_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_122_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_122_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_122_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_122_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_122_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_122_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_122_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__123_ccff_tail[0]),
    .chany_top_out(sb_1__1__112_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__112_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__112_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__112_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__112_ccff_tail[0])
  );


  sb_1__1_
  sb_11__4_
  (
    .clk_2_S_out(clk_2_wires[122]),
    .clk_2_N_out(clk_2_wires[120]),
    .clk_2_W_in(clk_2_wires[118]),
    .prog_clk_2_S_out(prog_clk_2_wires[122]),
    .prog_clk_2_N_out(prog_clk_2_wires[120]),
    .prog_clk_2_W_in(prog_clk_2_wires[118]),
    .prog_clk_0_N_in(prog_clk_0_wires[419]),
    .pReset_E_out(pResetWires[253]),
    .pReset_N_out(pResetWires[252]),
    .pReset_W_in(pResetWires[250]),
    .chany_top_in(cby_1__1__124_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_124_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_124_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_124_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_124_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_124_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_124_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_124_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_124_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__124_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_135_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_135_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_135_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_135_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_135_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_135_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_135_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_135_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__123_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_123_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_123_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_123_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_123_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_123_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_123_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_123_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_123_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__113_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_123_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_123_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_123_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_123_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_123_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_123_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_123_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_123_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__124_ccff_tail[0]),
    .chany_top_out(sb_1__1__113_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__113_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__113_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__113_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__113_ccff_tail[0])
  );


  sb_1__1_
  sb_11__5_
  (
    .clk_1_S_in(clk_2_wires[121]),
    .clk_1_W_out(clk_1_wires[226]),
    .clk_1_E_out(clk_1_wires[225]),
    .prog_clk_1_S_in(prog_clk_2_wires[121]),
    .prog_clk_1_W_out(prog_clk_1_wires[226]),
    .prog_clk_1_E_out(prog_clk_1_wires[225]),
    .prog_clk_0_N_in(prog_clk_0_wires[422]),
    .pReset_E_out(pResetWires[302]),
    .pReset_N_out(pResetWires[301]),
    .pReset_W_in(pResetWires[299]),
    .chany_top_in(cby_1__1__125_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_125_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_125_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_125_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_125_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_125_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_125_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_125_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_125_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__125_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_136_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_136_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_136_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_136_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_136_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_136_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_136_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_136_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__124_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_124_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_124_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_124_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_124_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_124_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_124_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_124_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_124_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__114_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_124_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_124_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_124_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_124_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_124_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_124_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_124_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_124_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__125_ccff_tail[0]),
    .chany_top_out(sb_1__1__114_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__114_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__114_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__114_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__114_ccff_tail[0])
  );


  sb_1__1_
  sb_11__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[425]),
    .pReset_E_out(pResetWires[351]),
    .pReset_N_out(pResetWires[350]),
    .pReset_W_in(pResetWires[348]),
    .chany_top_in(cby_1__1__126_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_126_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_126_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_126_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_126_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_126_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_126_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_126_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_126_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__126_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_137_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_137_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_137_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_137_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_137_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_137_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_137_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_137_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__125_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_125_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_125_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_125_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_125_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_125_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_125_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_125_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_125_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__115_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_125_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_125_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_125_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_125_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_125_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_125_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_125_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_125_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__126_ccff_tail[0]),
    .chany_top_out(sb_1__1__115_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__115_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__115_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__115_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__115_ccff_tail[0])
  );


  sb_1__1_
  sb_11__7_
  (
    .clk_1_N_in(clk_2_wires[130]),
    .clk_1_W_out(clk_1_wires[233]),
    .clk_1_E_out(clk_1_wires[232]),
    .prog_clk_1_N_in(prog_clk_2_wires[130]),
    .prog_clk_1_W_out(prog_clk_1_wires[233]),
    .prog_clk_1_E_out(prog_clk_1_wires[232]),
    .prog_clk_0_N_in(prog_clk_0_wires[428]),
    .pReset_E_out(pResetWires[400]),
    .pReset_N_out(pResetWires[399]),
    .pReset_W_in(pResetWires[397]),
    .chany_top_in(cby_1__1__127_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_127_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_127_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_127_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_127_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_127_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_127_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_127_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_127_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__127_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_138_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_138_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_138_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_138_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_138_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_138_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_138_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_138_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__126_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_126_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_126_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_126_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_126_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_126_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_126_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_126_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_126_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__116_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_126_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_126_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_126_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_126_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_126_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_126_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_126_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_126_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__127_ccff_tail[0]),
    .chany_top_out(sb_1__1__116_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__116_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__116_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__116_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__116_ccff_tail[0])
  );


  sb_1__1_
  sb_11__8_
  (
    .clk_2_S_out(clk_2_wires[129]),
    .clk_2_N_out(clk_2_wires[127]),
    .clk_2_W_in(clk_2_wires[125]),
    .prog_clk_2_S_out(prog_clk_2_wires[129]),
    .prog_clk_2_N_out(prog_clk_2_wires[127]),
    .prog_clk_2_W_in(prog_clk_2_wires[125]),
    .prog_clk_0_N_in(prog_clk_0_wires[431]),
    .pReset_E_out(pResetWires[449]),
    .pReset_N_out(pResetWires[448]),
    .pReset_W_in(pResetWires[446]),
    .chany_top_in(cby_1__1__128_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_128_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_128_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_128_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_128_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_128_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_128_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_128_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_128_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__128_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_139_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_139_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_139_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_139_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_139_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_139_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_139_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_139_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__127_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_127_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_127_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_127_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_127_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_127_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_127_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_127_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_127_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__117_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_127_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_127_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_127_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_127_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_127_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_127_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_127_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_127_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__128_ccff_tail[0]),
    .chany_top_out(sb_1__1__117_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__117_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__117_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__117_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__117_ccff_tail[0])
  );


  sb_1__1_
  sb_11__9_
  (
    .clk_1_S_in(clk_2_wires[128]),
    .clk_1_W_out(clk_1_wires[240]),
    .clk_1_E_out(clk_1_wires[239]),
    .prog_clk_1_S_in(prog_clk_2_wires[128]),
    .prog_clk_1_W_out(prog_clk_1_wires[240]),
    .prog_clk_1_E_out(prog_clk_1_wires[239]),
    .prog_clk_0_N_in(prog_clk_0_wires[434]),
    .pReset_E_out(pResetWires[498]),
    .pReset_N_out(pResetWires[497]),
    .pReset_W_in(pResetWires[495]),
    .chany_top_in(cby_1__1__129_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_129_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_129_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_129_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_129_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_129_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_129_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_129_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_129_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__129_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_140_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_140_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_140_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_140_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_140_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_140_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_140_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_140_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__128_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_128_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_128_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_128_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_128_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_128_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_128_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_128_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_128_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__118_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_128_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_128_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_128_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_128_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_128_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_128_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_128_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_128_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__129_ccff_tail[0]),
    .chany_top_out(sb_1__1__118_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__118_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__118_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__118_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__118_ccff_tail[0])
  );


  sb_1__1_
  sb_11__10_
  (
    .clk_2_N_out(clk_2_wires[134]),
    .clk_2_W_in(clk_2_wires[132]),
    .prog_clk_2_N_out(prog_clk_2_wires[134]),
    .prog_clk_2_W_in(prog_clk_2_wires[132]),
    .prog_clk_0_N_in(prog_clk_0_wires[437]),
    .pReset_E_out(pResetWires[547]),
    .pReset_N_out(pResetWires[546]),
    .pReset_W_in(pResetWires[544]),
    .chany_top_in(cby_1__1__130_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_130_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_130_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_130_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_130_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_130_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_130_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_130_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_130_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__130_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_141_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_141_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_141_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_141_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_141_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_141_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_141_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_141_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__129_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_129_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_129_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_129_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_129_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_129_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_129_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_129_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_129_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__119_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_129_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_129_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_129_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_129_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_129_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_129_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_129_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_129_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__130_ccff_tail[0]),
    .chany_top_out(sb_1__1__119_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__119_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__119_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__119_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__119_ccff_tail[0])
  );


  sb_1__1_
  sb_11__11_
  (
    .clk_1_S_in(clk_2_wires[135]),
    .clk_1_W_out(clk_1_wires[247]),
    .clk_1_E_out(clk_1_wires[246]),
    .prog_clk_1_S_in(prog_clk_2_wires[135]),
    .prog_clk_1_W_out(prog_clk_1_wires[247]),
    .prog_clk_1_E_out(prog_clk_1_wires[246]),
    .prog_clk_0_N_in(prog_clk_0_wires[440]),
    .pReset_E_out(pResetWires[596]),
    .pReset_N_out(pResetWires[595]),
    .pReset_W_in(pResetWires[593]),
    .chany_top_in(cby_1__1__131_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_131_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_131_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_131_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_131_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_131_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_131_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_131_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_131_right_width_0_height_0__pin_51_lower[0]),
    .chanx_right_in(cbx_1__1__131_chanx_left_out[0:29]),
    .right_bottom_grid_pin_36_(grid_clb_142_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_142_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_142_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_142_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_142_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_142_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_142_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_142_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__130_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_130_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_130_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_130_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_130_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_130_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_130_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_130_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_130_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__120_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_130_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_130_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_130_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_130_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_130_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_130_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_130_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_130_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(cbx_1__1__131_ccff_tail[0]),
    .chany_top_out(sb_1__1__120_chany_top_out[0:29]),
    .chanx_right_out(sb_1__1__120_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__1__120_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__1__120_chanx_left_out[0:29]),
    .ccff_tail(sb_1__1__120_ccff_tail[0])
  );


  sb_1__2_
  sb_1__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[60]),
    .pReset_E_in(pResetWires[604]),
    .pReset_W_out(pResetWires[601]),
    .chanx_right_in(cbx_1__12__1_chanx_left_out[0:29]),
    .right_top_grid_pin_1_(grid_io_top_1_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_23_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_23_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_23_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_23_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_23_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_23_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_23_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_23_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__11_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_11_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_11_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_11_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_11_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_11_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_11_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_11_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_11_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__12__0_chanx_right_out[0:29]),
    .left_top_grid_pin_1_(grid_io_top_0_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_11_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_11_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_11_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_11_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_11_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_11_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_11_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_11_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_top_1_ccff_tail[0]),
    .chanx_right_out(sb_1__12__0_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__12__0_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__12__0_chanx_left_out[0:29]),
    .ccff_tail(sb_1__12__0_ccff_tail[0])
  );


  sb_1__2_
  sb_2__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[100]),
    .pReset_E_in(pResetWires[607]),
    .pReset_W_out(pResetWires[605]),
    .SC_OUT_BOT(scff_Wires[53]),
    .SC_IN_BOT(scff_Wires[52]),
    .chanx_right_in(cbx_1__12__2_chanx_left_out[0:29]),
    .right_top_grid_pin_1_(grid_io_top_2_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_35_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_35_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_35_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_35_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_35_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_35_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_35_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_35_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__23_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_23_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_23_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_23_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_23_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_23_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_23_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_23_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_23_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__12__1_chanx_right_out[0:29]),
    .left_top_grid_pin_1_(grid_io_top_1_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_23_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_23_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_23_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_23_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_23_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_23_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_23_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_23_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_top_2_ccff_tail[0]),
    .chanx_right_out(sb_1__12__1_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__12__1_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__12__1_chanx_left_out[0:29]),
    .ccff_tail(sb_1__12__1_ccff_tail[0])
  );


  sb_1__2_
  sb_3__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[138]),
    .pReset_E_in(pResetWires[610]),
    .pReset_W_out(pResetWires[608]),
    .chanx_right_in(cbx_1__12__3_chanx_left_out[0:29]),
    .right_top_grid_pin_1_(grid_io_top_3_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_47_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_47_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_47_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_47_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_47_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_47_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_47_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_47_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__35_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_35_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_35_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_35_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_35_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_35_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_35_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_35_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_35_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__12__2_chanx_right_out[0:29]),
    .left_top_grid_pin_1_(grid_io_top_2_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_35_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_35_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_35_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_35_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_35_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_35_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_35_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_35_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_top_3_ccff_tail[0]),
    .chanx_right_out(sb_1__12__2_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__12__2_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__12__2_chanx_left_out[0:29]),
    .ccff_tail(sb_1__12__2_ccff_tail[0])
  );


  sb_1__2_
  sb_4__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[176]),
    .pReset_E_in(pResetWires[613]),
    .pReset_W_out(pResetWires[611]),
    .SC_OUT_BOT(scff_Wires[106]),
    .SC_IN_BOT(scff_Wires[105]),
    .chanx_right_in(cbx_1__12__4_chanx_left_out[0:29]),
    .right_top_grid_pin_1_(grid_io_top_4_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_59_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_59_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_59_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_59_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_59_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_59_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_59_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_59_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__47_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_47_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_47_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_47_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_47_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_47_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_47_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_47_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_47_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__12__3_chanx_right_out[0:29]),
    .left_top_grid_pin_1_(grid_io_top_3_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_47_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_47_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_47_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_47_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_47_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_47_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_47_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_47_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_top_4_ccff_tail[0]),
    .chanx_right_out(sb_1__12__3_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__12__3_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__12__3_chanx_left_out[0:29]),
    .ccff_tail(sb_1__12__3_ccff_tail[0])
  );


  sb_1__2_
  sb_5__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[214]),
    .pReset_E_in(pResetWires[616]),
    .pReset_W_out(pResetWires[614]),
    .chanx_right_in(cbx_1__12__5_chanx_left_out[0:29]),
    .right_top_grid_pin_1_(grid_io_top_5_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_71_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_71_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_71_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_71_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_71_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_71_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_71_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_71_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__59_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_59_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_59_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_59_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_59_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_59_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_59_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_59_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_59_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__12__4_chanx_right_out[0:29]),
    .left_top_grid_pin_1_(grid_io_top_4_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_59_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_59_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_59_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_59_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_59_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_59_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_59_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_59_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_top_5_ccff_tail[0]),
    .chanx_right_out(sb_1__12__4_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__12__4_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__12__4_chanx_left_out[0:29]),
    .ccff_tail(sb_1__12__4_ccff_tail[0])
  );


  sb_1__2_
  sb_6__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[252]),
    .pReset_E_out(pResetWires[619]),
    .pReset_W_out(pResetWires[617]),
    .pReset_S_in(pResetWires[24]),
    .SC_OUT_BOT(scff_Wires[159]),
    .SC_IN_BOT(scff_Wires[158]),
    .chanx_right_in(cbx_1__12__6_chanx_left_out[0:29]),
    .right_top_grid_pin_1_(grid_io_top_6_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_83_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_83_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_83_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_83_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_83_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_83_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_83_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_83_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__71_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_71_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_71_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_71_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_71_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_71_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_71_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_71_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_71_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__12__5_chanx_right_out[0:29]),
    .left_top_grid_pin_1_(grid_io_top_5_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_71_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_71_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_71_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_71_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_71_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_71_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_71_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_71_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_top_6_ccff_tail[0]),
    .chanx_right_out(sb_1__12__5_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__12__5_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__12__5_chanx_left_out[0:29]),
    .ccff_tail(sb_1__12__5_ccff_tail[0])
  );


  sb_1__2_
  sb_7__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[290]),
    .pReset_E_out(pResetWires[622]),
    .pReset_W_in(pResetWires[620]),
    .chanx_right_in(cbx_1__12__7_chanx_left_out[0:29]),
    .right_top_grid_pin_1_(grid_io_top_7_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_95_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_95_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_95_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_95_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_95_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_95_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_95_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_95_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__83_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_83_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_83_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_83_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_83_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_83_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_83_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_83_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_83_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__12__6_chanx_right_out[0:29]),
    .left_top_grid_pin_1_(grid_io_top_6_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_83_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_83_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_83_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_83_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_83_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_83_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_83_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_83_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_top_7_ccff_tail[0]),
    .chanx_right_out(sb_1__12__6_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__12__6_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__12__6_chanx_left_out[0:29]),
    .ccff_tail(sb_1__12__6_ccff_tail[0])
  );


  sb_1__2_
  sb_8__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[328]),
    .pReset_E_out(pResetWires[625]),
    .pReset_W_in(pResetWires[623]),
    .SC_OUT_BOT(scff_Wires[212]),
    .SC_IN_BOT(scff_Wires[211]),
    .chanx_right_in(cbx_1__12__8_chanx_left_out[0:29]),
    .right_top_grid_pin_1_(grid_io_top_8_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_107_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_107_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_107_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_107_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_107_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_107_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_107_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_107_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__95_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_95_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_95_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_95_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_95_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_95_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_95_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_95_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_95_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__12__7_chanx_right_out[0:29]),
    .left_top_grid_pin_1_(grid_io_top_7_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_95_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_95_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_95_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_95_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_95_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_95_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_95_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_95_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_top_8_ccff_tail[0]),
    .chanx_right_out(sb_1__12__7_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__12__7_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__12__7_chanx_left_out[0:29]),
    .ccff_tail(sb_1__12__7_ccff_tail[0])
  );


  sb_1__2_
  sb_9__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[366]),
    .pReset_E_out(pResetWires[628]),
    .pReset_W_in(pResetWires[626]),
    .chanx_right_in(cbx_1__12__9_chanx_left_out[0:29]),
    .right_top_grid_pin_1_(grid_io_top_9_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_119_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_119_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_119_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_119_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_119_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_119_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_119_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_119_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__107_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_107_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_107_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_107_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_107_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_107_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_107_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_107_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_107_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__12__8_chanx_right_out[0:29]),
    .left_top_grid_pin_1_(grid_io_top_8_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_107_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_107_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_107_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_107_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_107_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_107_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_107_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_107_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_top_9_ccff_tail[0]),
    .chanx_right_out(sb_1__12__8_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__12__8_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__12__8_chanx_left_out[0:29]),
    .ccff_tail(sb_1__12__8_ccff_tail[0])
  );


  sb_1__2_
  sb_10__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[404]),
    .pReset_E_out(pResetWires[631]),
    .pReset_W_in(pResetWires[629]),
    .SC_OUT_BOT(scff_Wires[265]),
    .SC_IN_BOT(scff_Wires[264]),
    .chanx_right_in(cbx_1__12__10_chanx_left_out[0:29]),
    .right_top_grid_pin_1_(grid_io_top_10_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_131_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_131_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_131_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_131_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_131_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_131_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_131_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_131_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__119_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_119_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_119_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_119_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_119_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_119_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_119_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_119_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_119_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__12__9_chanx_right_out[0:29]),
    .left_top_grid_pin_1_(grid_io_top_9_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_119_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_119_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_119_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_119_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_119_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_119_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_119_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_119_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_top_10_ccff_tail[0]),
    .chanx_right_out(sb_1__12__9_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__12__9_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__12__9_chanx_left_out[0:29]),
    .ccff_tail(sb_1__12__9_ccff_tail[0])
  );


  sb_1__2_
  sb_11__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[442]),
    .pReset_E_out(pResetWires[634]),
    .pReset_W_in(pResetWires[632]),
    .chanx_right_in(cbx_1__12__11_chanx_left_out[0:29]),
    .right_top_grid_pin_1_(grid_io_top_11_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_143_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_143_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_143_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_143_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_143_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_143_top_width_0_height_0__pin_41_upper[0]),
    .right_bottom_grid_pin_42_(grid_clb_143_top_width_0_height_0__pin_42_upper[0]),
    .right_bottom_grid_pin_43_(grid_clb_143_top_width_0_height_0__pin_43_upper[0]),
    .chany_bottom_in(cby_1__1__131_chany_top_out[0:29]),
    .bottom_left_grid_pin_44_(grid_clb_131_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_131_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_131_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_131_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_131_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_131_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_131_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_131_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__12__10_chanx_right_out[0:29]),
    .left_top_grid_pin_1_(grid_io_top_10_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_131_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_131_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_131_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_131_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_131_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_131_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_131_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_131_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_top_11_ccff_tail[0]),
    .chanx_right_out(sb_1__12__10_chanx_right_out[0:29]),
    .chany_bottom_out(sb_1__12__10_chany_bottom_out[0:29]),
    .chanx_left_out(sb_1__12__10_chanx_left_out[0:29]),
    .ccff_tail(sb_1__12__10_ccff_tail[0])
  );


  sb_2__0_
  sb_12__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[445]),
    .pReset_N_out(pResetWires[60]),
    .pReset_W_in(pResetWires[59]),
    .chany_top_in(cby_12__1__0_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_132_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_132_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_132_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_132_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_132_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_132_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_132_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_132_right_width_0_height_0__pin_51_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_11_left_width_0_height_0__pin_1_lower[0]),
    .chanx_left_in(cbx_1__0__11_chanx_right_out[0:29]),
    .left_bottom_grid_pin_1_(grid_io_bottom_0_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_0_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_0_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_0_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_0_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_0_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_0_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_0_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_0_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_right_11_ccff_tail[0]),
    .chany_top_out(sb_12__0__0_chany_top_out[0:29]),
    .chanx_left_out(sb_12__0__0_chanx_left_out[0:29]),
    .ccff_tail(sb_12__0__0_ccff_tail[0])
  );


  sb_2__1_
  sb_12__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[448]),
    .pReset_N_out(pResetWires[109]),
    .pReset_W_in(pResetWires[107]),
    .chany_top_in(cby_12__1__1_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_133_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_133_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_133_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_133_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_133_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_133_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_133_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_133_right_width_0_height_0__pin_51_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_10_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__0_chany_top_out[0:29]),
    .bottom_right_grid_pin_1_(grid_io_right_11_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_132_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_132_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_132_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_132_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_132_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_132_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_132_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_132_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__121_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_132_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_132_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_132_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_132_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_132_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_132_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_132_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_132_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_right_10_ccff_tail[0]),
    .chany_top_out(sb_12__1__0_chany_top_out[0:29]),
    .chany_bottom_out(sb_12__1__0_chany_bottom_out[0:29]),
    .chanx_left_out(sb_12__1__0_chanx_left_out[0:29]),
    .ccff_tail(sb_12__1__0_ccff_tail[0])
  );


  sb_2__1_
  sb_12__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[451]),
    .pReset_N_out(pResetWires[158]),
    .pReset_W_in(pResetWires[156]),
    .chany_top_in(cby_12__1__2_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_134_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_134_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_134_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_134_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_134_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_134_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_134_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_134_right_width_0_height_0__pin_51_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_9_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__1_chany_top_out[0:29]),
    .bottom_right_grid_pin_1_(grid_io_right_10_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_133_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_133_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_133_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_133_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_133_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_133_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_133_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_133_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__122_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_133_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_133_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_133_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_133_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_133_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_133_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_133_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_133_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_right_9_ccff_tail[0]),
    .chany_top_out(sb_12__1__1_chany_top_out[0:29]),
    .chany_bottom_out(sb_12__1__1_chany_bottom_out[0:29]),
    .chanx_left_out(sb_12__1__1_chanx_left_out[0:29]),
    .ccff_tail(sb_12__1__1_ccff_tail[0])
  );


  sb_2__1_
  sb_12__3_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[454]),
    .pReset_N_out(pResetWires[207]),
    .pReset_W_in(pResetWires[205]),
    .chany_top_in(cby_12__1__3_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_135_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_135_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_135_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_135_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_135_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_135_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_135_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_135_right_width_0_height_0__pin_51_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_8_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__2_chany_top_out[0:29]),
    .bottom_right_grid_pin_1_(grid_io_right_9_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_134_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_134_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_134_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_134_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_134_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_134_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_134_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_134_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__123_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_134_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_134_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_134_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_134_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_134_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_134_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_134_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_134_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_right_8_ccff_tail[0]),
    .chany_top_out(sb_12__1__2_chany_top_out[0:29]),
    .chany_bottom_out(sb_12__1__2_chany_bottom_out[0:29]),
    .chanx_left_out(sb_12__1__2_chanx_left_out[0:29]),
    .ccff_tail(sb_12__1__2_ccff_tail[0])
  );


  sb_2__1_
  sb_12__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[457]),
    .pReset_N_out(pResetWires[256]),
    .pReset_W_in(pResetWires[254]),
    .chany_top_in(cby_12__1__4_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_136_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_136_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_136_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_136_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_136_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_136_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_136_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_136_right_width_0_height_0__pin_51_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_7_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__3_chany_top_out[0:29]),
    .bottom_right_grid_pin_1_(grid_io_right_8_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_135_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_135_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_135_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_135_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_135_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_135_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_135_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_135_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__124_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_135_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_135_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_135_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_135_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_135_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_135_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_135_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_135_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_right_7_ccff_tail[0]),
    .chany_top_out(sb_12__1__3_chany_top_out[0:29]),
    .chany_bottom_out(sb_12__1__3_chany_bottom_out[0:29]),
    .chanx_left_out(sb_12__1__3_chanx_left_out[0:29]),
    .ccff_tail(sb_12__1__3_ccff_tail[0])
  );


  sb_2__1_
  sb_12__5_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[460]),
    .pReset_N_out(pResetWires[305]),
    .pReset_W_in(pResetWires[303]),
    .chany_top_in(cby_12__1__5_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_137_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_137_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_137_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_137_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_137_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_137_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_137_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_137_right_width_0_height_0__pin_51_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_6_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__4_chany_top_out[0:29]),
    .bottom_right_grid_pin_1_(grid_io_right_7_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_136_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_136_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_136_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_136_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_136_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_136_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_136_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_136_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__125_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_136_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_136_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_136_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_136_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_136_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_136_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_136_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_136_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_right_6_ccff_tail[0]),
    .chany_top_out(sb_12__1__4_chany_top_out[0:29]),
    .chany_bottom_out(sb_12__1__4_chany_bottom_out[0:29]),
    .chanx_left_out(sb_12__1__4_chanx_left_out[0:29]),
    .ccff_tail(sb_12__1__4_ccff_tail[0])
  );


  sb_2__1_
  sb_12__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[463]),
    .pReset_N_out(pResetWires[354]),
    .pReset_W_in(pResetWires[352]),
    .chany_top_in(cby_12__1__6_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_138_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_138_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_138_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_138_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_138_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_138_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_138_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_138_right_width_0_height_0__pin_51_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_5_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__5_chany_top_out[0:29]),
    .bottom_right_grid_pin_1_(grid_io_right_6_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_137_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_137_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_137_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_137_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_137_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_137_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_137_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_137_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__126_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_137_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_137_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_137_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_137_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_137_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_137_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_137_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_137_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_right_5_ccff_tail[0]),
    .chany_top_out(sb_12__1__5_chany_top_out[0:29]),
    .chany_bottom_out(sb_12__1__5_chany_bottom_out[0:29]),
    .chanx_left_out(sb_12__1__5_chanx_left_out[0:29]),
    .ccff_tail(sb_12__1__5_ccff_tail[0])
  );


  sb_2__1_
  sb_12__7_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[466]),
    .pReset_N_out(pResetWires[403]),
    .pReset_W_in(pResetWires[401]),
    .chany_top_in(cby_12__1__7_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_139_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_139_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_139_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_139_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_139_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_139_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_139_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_139_right_width_0_height_0__pin_51_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_4_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__6_chany_top_out[0:29]),
    .bottom_right_grid_pin_1_(grid_io_right_5_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_138_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_138_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_138_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_138_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_138_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_138_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_138_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_138_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__127_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_138_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_138_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_138_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_138_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_138_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_138_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_138_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_138_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_right_4_ccff_tail[0]),
    .chany_top_out(sb_12__1__6_chany_top_out[0:29]),
    .chany_bottom_out(sb_12__1__6_chany_bottom_out[0:29]),
    .chanx_left_out(sb_12__1__6_chanx_left_out[0:29]),
    .ccff_tail(sb_12__1__6_ccff_tail[0])
  );


  sb_2__1_
  sb_12__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[469]),
    .pReset_N_out(pResetWires[452]),
    .pReset_W_in(pResetWires[450]),
    .chany_top_in(cby_12__1__8_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_140_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_140_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_140_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_140_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_140_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_140_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_140_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_140_right_width_0_height_0__pin_51_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_3_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__7_chany_top_out[0:29]),
    .bottom_right_grid_pin_1_(grid_io_right_4_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_139_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_139_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_139_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_139_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_139_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_139_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_139_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_139_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__128_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_139_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_139_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_139_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_139_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_139_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_139_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_139_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_139_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_right_3_ccff_tail[0]),
    .chany_top_out(sb_12__1__7_chany_top_out[0:29]),
    .chany_bottom_out(sb_12__1__7_chany_bottom_out[0:29]),
    .chanx_left_out(sb_12__1__7_chanx_left_out[0:29]),
    .ccff_tail(sb_12__1__7_ccff_tail[0])
  );


  sb_2__1_
  sb_12__9_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[472]),
    .pReset_N_out(pResetWires[501]),
    .pReset_W_in(pResetWires[499]),
    .chany_top_in(cby_12__1__9_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_141_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_141_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_141_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_141_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_141_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_141_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_141_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_141_right_width_0_height_0__pin_51_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_2_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__8_chany_top_out[0:29]),
    .bottom_right_grid_pin_1_(grid_io_right_3_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_140_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_140_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_140_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_140_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_140_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_140_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_140_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_140_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__129_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_140_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_140_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_140_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_140_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_140_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_140_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_140_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_140_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_right_2_ccff_tail[0]),
    .chany_top_out(sb_12__1__8_chany_top_out[0:29]),
    .chany_bottom_out(sb_12__1__8_chany_bottom_out[0:29]),
    .chanx_left_out(sb_12__1__8_chanx_left_out[0:29]),
    .ccff_tail(sb_12__1__8_ccff_tail[0])
  );


  sb_2__1_
  sb_12__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[475]),
    .pReset_N_out(pResetWires[550]),
    .pReset_W_in(pResetWires[548]),
    .chany_top_in(cby_12__1__10_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_142_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_142_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_142_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_142_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_142_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_142_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_142_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_142_right_width_0_height_0__pin_51_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_1_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__9_chany_top_out[0:29]),
    .bottom_right_grid_pin_1_(grid_io_right_2_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_141_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_141_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_141_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_141_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_141_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_141_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_141_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_141_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__130_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_141_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_141_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_141_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_141_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_141_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_141_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_141_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_141_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_right_1_ccff_tail[0]),
    .chany_top_out(sb_12__1__9_chany_top_out[0:29]),
    .chany_bottom_out(sb_12__1__9_chany_bottom_out[0:29]),
    .chanx_left_out(sb_12__1__9_chanx_left_out[0:29]),
    .ccff_tail(sb_12__1__9_ccff_tail[0])
  );


  sb_2__1_
  sb_12__11_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[478]),
    .pReset_N_out(pResetWires[599]),
    .pReset_W_in(pResetWires[597]),
    .chany_top_in(cby_12__1__11_chany_bottom_out[0:29]),
    .top_left_grid_pin_44_(grid_clb_143_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_143_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_143_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_143_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_143_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_143_right_width_0_height_0__pin_49_lower[0]),
    .top_left_grid_pin_50_(grid_clb_143_right_width_0_height_0__pin_50_lower[0]),
    .top_left_grid_pin_51_(grid_clb_143_right_width_0_height_0__pin_51_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_0_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_12__1__10_chany_top_out[0:29]),
    .bottom_right_grid_pin_1_(grid_io_right_1_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_142_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_142_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_142_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_142_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_142_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_142_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_142_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_142_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__1__131_chanx_right_out[0:29]),
    .left_bottom_grid_pin_36_(grid_clb_142_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_142_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_142_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_142_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_142_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_142_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_142_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_142_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(grid_io_right_0_ccff_tail[0]),
    .chany_top_out(sb_12__1__10_chany_top_out[0:29]),
    .chany_bottom_out(sb_12__1__10_chany_bottom_out[0:29]),
    .chanx_left_out(sb_12__1__10_chanx_left_out[0:29]),
    .ccff_tail(sb_12__1__10_ccff_tail[0])
  );


  sb_2__2_
  sb_12__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[480]),
    .pReset_W_in(pResetWires[635]),
    .SC_OUT_BOT(sc_tail),
    .SC_IN_BOT(scff_Wires[317]),
    .chany_bottom_in(cby_12__1__11_chany_top_out[0:29]),
    .bottom_right_grid_pin_1_(grid_io_right_0_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_143_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_143_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_143_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_143_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_143_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_143_right_width_0_height_0__pin_49_upper[0]),
    .bottom_left_grid_pin_50_(grid_clb_143_right_width_0_height_0__pin_50_upper[0]),
    .bottom_left_grid_pin_51_(grid_clb_143_right_width_0_height_0__pin_51_upper[0]),
    .chanx_left_in(cbx_1__12__11_chanx_right_out[0:29]),
    .left_top_grid_pin_1_(grid_io_top_11_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_143_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_143_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_143_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_143_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_143_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_143_top_width_0_height_0__pin_41_lower[0]),
    .left_bottom_grid_pin_42_(grid_clb_143_top_width_0_height_0__pin_42_lower[0]),
    .left_bottom_grid_pin_43_(grid_clb_143_top_width_0_height_0__pin_43_lower[0]),
    .ccff_head(ccff_head[0]),
    .chany_bottom_out(sb_12__12__0_chany_bottom_out[0:29]),
    .chanx_left_out(sb_12__12__0_chanx_left_out[0:29]),
    .ccff_tail(sb_12__12__0_ccff_tail[0])
  );


  cbx_1__0_
  cbx_1__0_
  (
    .prog_clk_0_W_out(prog_clk_0_wires[5]),
    .prog_clk_0_N_in(prog_clk_0_wires[0]),
    .pReset_E_in(pResetWires[26]),
    .pReset_W_out(pResetWires[25]),
    .SC_OUT_BOT(scff_Wires[26]),
    .SC_IN_TOP(scff_Wires[25]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_11_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_11_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_11_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_11_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_11_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_11_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_11_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_11_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_11_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_11_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_11_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_11_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_11_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_11_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_11_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_11_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_11_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_11_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__0_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__0_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__0_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__0_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__0_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__0_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__0_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__0_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__0_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[123:131]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[123:131]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[123:131]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_0__0__0_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__0__0_chanx_left_out[0:29]),
    .ccff_head(sb_1__0__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__0_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__0__0_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__0__0_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__0_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__0_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__0_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__0_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__0_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__0_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__0_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__0_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_11_ccff_tail[0])
  );


  cbx_1__0_
  cbx_2__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[63]),
    .pReset_E_in(pResetWires[29]),
    .pReset_W_out(pResetWires[28]),
    .SC_OUT_TOP(scff_Wires[28]),
    .SC_IN_BOT(scff_Wires[27]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_10_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_10_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_10_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_10_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_10_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_10_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_10_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_10_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_10_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_10_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_10_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_10_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_10_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_10_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_10_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_10_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_10_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_10_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__1_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__1_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__1_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__1_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__1_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__1_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__1_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__1_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__1_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[114:122]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[114:122]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[114:122]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__0_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__0__1_chanx_left_out[0:29]),
    .ccff_head(sb_1__0__1_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__1_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__0__1_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__0__1_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__1_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__1_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__1_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__1_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__1_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__1_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__1_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__1_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_10_ccff_tail[0])
  );


  cbx_1__0_
  cbx_3__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[101]),
    .pReset_E_in(pResetWires[32]),
    .pReset_W_out(pResetWires[31]),
    .SC_OUT_BOT(scff_Wires[79]),
    .SC_IN_TOP(scff_Wires[78]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_9_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_9_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_9_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_9_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_9_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_9_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_9_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_9_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_9_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_9_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_9_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_9_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_9_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_9_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_9_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_9_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_9_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_9_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__2_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__2_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__2_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__2_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__2_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__2_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__2_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__2_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__2_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[105:113]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[105:113]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[105:113]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__1_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__0__2_chanx_left_out[0:29]),
    .ccff_head(sb_1__0__2_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__2_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__0__2_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__0__2_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__2_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__2_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__2_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__2_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__2_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__2_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__2_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__2_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_9_ccff_tail[0])
  );


  cbx_1__0_
  cbx_4__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[139]),
    .pReset_E_in(pResetWires[35]),
    .pReset_W_out(pResetWires[34]),
    .SC_OUT_TOP(scff_Wires[81]),
    .SC_IN_BOT(scff_Wires[80]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_8_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_8_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_8_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_8_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_8_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_8_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_8_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_8_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_8_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_8_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_8_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_8_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_8_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_8_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_8_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_8_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_8_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_8_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__3_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__3_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__3_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__3_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__3_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__3_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__3_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__3_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__3_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[96:104]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[96:104]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[96:104]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__2_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__0__3_chanx_left_out[0:29]),
    .ccff_head(sb_1__0__3_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__3_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__0__3_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__0__3_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__3_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__3_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__3_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__3_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__3_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__3_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__3_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__3_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_8_ccff_tail[0])
  );


  cbx_1__0_
  cbx_5__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[177]),
    .pReset_E_in(pResetWires[38]),
    .pReset_W_out(pResetWires[37]),
    .SC_OUT_BOT(scff_Wires[132]),
    .SC_IN_TOP(scff_Wires[131]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_7_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_7_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_7_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_7_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_7_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_7_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_7_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_7_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_7_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_7_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_7_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_7_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_7_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_7_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_7_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_7_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_7_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_7_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__4_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__4_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__4_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__4_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__4_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__4_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__4_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__4_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__4_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87:95]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87:95]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87:95]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__3_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__0__4_chanx_left_out[0:29]),
    .ccff_head(sb_1__0__4_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__4_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__0__4_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__0__4_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__4_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__4_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__4_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__4_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__4_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__4_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__4_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__4_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_7_ccff_tail[0])
  );


  cbx_1__0_
  cbx_6__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[215]),
    .pReset_E_in(pResetWires[41]),
    .pReset_W_out(pResetWires[40]),
    .SC_OUT_TOP(scff_Wires[134]),
    .SC_IN_BOT(scff_Wires[133]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_6_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_6_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_6_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_6_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_6_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_6_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_6_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_6_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_6_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_6_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_6_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_6_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_6_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_6_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_6_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_6_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_6_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_6_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__5_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__5_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__5_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__5_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__5_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__5_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__5_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__5_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__5_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78:86]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78:86]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78:86]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__4_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__0__5_chanx_left_out[0:29]),
    .ccff_head(sb_1__0__5_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__5_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__0__5_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__0__5_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__5_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__5_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__5_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__5_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__5_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__5_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__5_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__5_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_6_ccff_tail[0])
  );


  cbx_1__0_
  cbx_7__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[253]),
    .pReset_E_out(pResetWires[44]),
    .pReset_W_in(pResetWires[43]),
    .SC_OUT_BOT(scff_Wires[185]),
    .SC_IN_TOP(scff_Wires[184]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_5_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_5_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_5_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_5_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_5_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_5_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_5_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_5_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_5_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_5_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_5_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_5_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_5_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_5_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_5_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_5_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_5_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_5_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__6_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__6_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__6_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__6_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__6_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__6_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__6_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__6_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__6_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69:77]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69:77]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69:77]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__5_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__0__6_chanx_left_out[0:29]),
    .ccff_head(sb_1__0__6_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__6_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__0__6_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__0__6_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__6_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__6_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__6_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__6_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__6_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__6_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__6_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__6_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_5_ccff_tail[0])
  );


  cbx_1__0_
  cbx_8__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[291]),
    .pReset_E_out(pResetWires[47]),
    .pReset_W_in(pResetWires[46]),
    .SC_OUT_TOP(scff_Wires[187]),
    .SC_IN_BOT(scff_Wires[186]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_4_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_4_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_4_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_4_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_4_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_4_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_4_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_4_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_4_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_4_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_4_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_4_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_4_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_4_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_4_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_4_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_4_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_4_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__7_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__7_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__7_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__7_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__7_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__7_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__7_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__7_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__7_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60:68]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60:68]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60:68]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__6_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__0__7_chanx_left_out[0:29]),
    .ccff_head(sb_1__0__7_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__7_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__0__7_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__0__7_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__7_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__7_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__7_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__7_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__7_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__7_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__7_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__7_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_4_ccff_tail[0])
  );


  cbx_1__0_
  cbx_9__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[329]),
    .pReset_E_out(pResetWires[50]),
    .pReset_W_in(pResetWires[49]),
    .SC_OUT_BOT(scff_Wires[238]),
    .SC_IN_TOP(scff_Wires[237]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_3_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_3_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_3_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_3_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_3_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_3_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_3_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_3_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_3_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_3_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_3_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_3_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_3_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_3_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_3_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_3_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_3_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_3_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__8_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__8_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__8_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__8_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__8_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__8_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__8_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__8_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__8_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51:59]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51:59]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51:59]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__7_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__0__8_chanx_left_out[0:29]),
    .ccff_head(sb_1__0__8_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__8_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__0__8_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__0__8_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__8_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__8_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__8_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__8_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__8_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__8_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__8_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__8_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_3_ccff_tail[0])
  );


  cbx_1__0_
  cbx_10__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[367]),
    .pReset_E_out(pResetWires[53]),
    .pReset_W_in(pResetWires[52]),
    .SC_OUT_TOP(scff_Wires[240]),
    .SC_IN_BOT(scff_Wires[239]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_2_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_2_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_2_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_2_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_2_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_2_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_2_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_2_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_2_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_2_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_2_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_2_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_2_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_2_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_2_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_2_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_2_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_2_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__9_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__9_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__9_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__9_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__9_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__9_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__9_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__9_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__9_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42:50]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42:50]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42:50]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__8_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__0__9_chanx_left_out[0:29]),
    .ccff_head(sb_1__0__9_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__9_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__0__9_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__0__9_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__9_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__9_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__9_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__9_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__9_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__9_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__9_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__9_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_2_ccff_tail[0])
  );


  cbx_1__0_
  cbx_11__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[405]),
    .pReset_E_out(pResetWires[56]),
    .pReset_W_in(pResetWires[55]),
    .SC_OUT_BOT(scff_Wires[291]),
    .SC_IN_TOP(scff_Wires[290]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_1_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_1_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_1_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_1_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_1_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_1_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_1_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_1_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_1_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_1_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_1_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_1_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_1_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_1_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_1_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_1_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_1_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_1_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__10_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__10_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__10_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__10_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__10_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__10_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__10_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__10_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__10_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33:41]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33:41]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33:41]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__9_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__0__10_chanx_left_out[0:29]),
    .ccff_head(sb_1__0__10_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__10_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__0__10_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__0__10_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__10_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__10_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__10_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__10_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__10_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__10_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__10_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__10_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_1_ccff_tail[0])
  );


  cbx_1__0_
  cbx_12__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[443]),
    .pReset_E_out(pResetWires[59]),
    .pReset_W_in(pResetWires[58]),
    .SC_OUT_TOP(scff_Wires[293]),
    .SC_IN_BOT(scff_Wires[292]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_0_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_0_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_0_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_0_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_0_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_0_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_0_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_0_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_0_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_0_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_0_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_0_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_0_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_0_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_0_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_0_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_0_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_0_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__11_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__11_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__11_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__11_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__11_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__11_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__11_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__11_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__11_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24:32]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24:32]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24:32]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__10_chanx_right_out[0:29]),
    .chanx_right_in(sb_12__0__0_chanx_left_out[0:29]),
    .ccff_head(sb_12__0__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__11_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__0__11_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__0__11_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__11_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__11_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__11_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__11_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__11_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__11_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__11_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__11_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_0_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__1_
  (
    .clk_1_S_out(clk_1_wires[4]),
    .clk_1_N_out(clk_1_wires[3]),
    .clk_1_E_in(clk_1_wires[2]),
    .prog_clk_1_S_out(prog_clk_1_wires[4]),
    .prog_clk_1_N_out(prog_clk_1_wires[3]),
    .prog_clk_1_E_in(prog_clk_1_wires[2]),
    .prog_clk_0_N_in(prog_clk_0_wires[6]),
    .prog_clk_0_W_out(prog_clk_0_wires[4]),
    .pReset_S_out(pResetWires[63]),
    .pReset_E_in(pResetWires[62]),
    .pReset_W_out(pResetWires[61]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[0]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[0]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[0]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[0]),
    .SC_OUT_BOT(scff_Wires[23]),
    .SC_IN_TOP(scff_Wires[22]),
    .chanx_left_in(sb_0__1__0_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__0_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__0_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__0_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__0_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__0_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__0_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__0_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__0_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__0_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__0_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__0_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__0_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__0_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__0_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__0_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__0_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__0_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__0_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__0_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__0_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[11]),
    .prog_clk_0_W_out(prog_clk_0_wires[10]),
    .pReset_S_out(pResetWires[112]),
    .pReset_E_in(pResetWires[111]),
    .pReset_W_out(pResetWires[110]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[1]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[1]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[1]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[1]),
    .SC_OUT_BOT(scff_Wires[21]),
    .SC_IN_TOP(scff_Wires[20]),
    .chanx_left_in(sb_0__1__1_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__1_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__1_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__1_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__1_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__1_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__1_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__1_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__1_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__1_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__1_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__1_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__1_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__1_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__1_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__1_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__1_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__1_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__1_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__1_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__1_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__1_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__3_
  (
    .clk_1_S_out(clk_1_wires[11]),
    .clk_1_N_out(clk_1_wires[10]),
    .clk_1_E_in(clk_1_wires[9]),
    .prog_clk_1_S_out(prog_clk_1_wires[11]),
    .prog_clk_1_N_out(prog_clk_1_wires[10]),
    .prog_clk_1_E_in(prog_clk_1_wires[9]),
    .prog_clk_0_N_in(prog_clk_0_wires[16]),
    .prog_clk_0_W_out(prog_clk_0_wires[15]),
    .pReset_S_out(pResetWires[161]),
    .pReset_E_in(pResetWires[160]),
    .pReset_W_out(pResetWires[159]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[2]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[2]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[2]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[2]),
    .SC_OUT_BOT(scff_Wires[19]),
    .SC_IN_TOP(scff_Wires[18]),
    .chanx_left_in(sb_0__1__2_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__2_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__2_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__2_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__2_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__2_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__2_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__2_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__2_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__2_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__2_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__2_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__2_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__2_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__2_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__2_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__2_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__2_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__2_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__2_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__2_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__2_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[21]),
    .prog_clk_0_W_out(prog_clk_0_wires[20]),
    .pReset_S_out(pResetWires[210]),
    .pReset_E_in(pResetWires[209]),
    .pReset_W_out(pResetWires[208]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[3]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[3]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[3]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[3]),
    .SC_OUT_BOT(scff_Wires[17]),
    .SC_IN_TOP(scff_Wires[16]),
    .chanx_left_in(sb_0__1__3_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__3_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__3_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__3_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__3_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__3_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__3_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__3_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__3_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__3_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__3_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__3_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__3_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__3_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__3_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__3_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__3_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__3_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__3_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__3_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__3_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__3_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__5_
  (
    .clk_1_S_out(clk_1_wires[18]),
    .clk_1_N_out(clk_1_wires[17]),
    .clk_1_E_in(clk_1_wires[16]),
    .prog_clk_1_S_out(prog_clk_1_wires[18]),
    .prog_clk_1_N_out(prog_clk_1_wires[17]),
    .prog_clk_1_E_in(prog_clk_1_wires[16]),
    .prog_clk_0_N_in(prog_clk_0_wires[26]),
    .prog_clk_0_W_out(prog_clk_0_wires[25]),
    .pReset_S_out(pResetWires[259]),
    .pReset_E_in(pResetWires[258]),
    .pReset_W_out(pResetWires[257]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[4]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[4]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[4]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[4]),
    .SC_OUT_BOT(scff_Wires[15]),
    .SC_IN_TOP(scff_Wires[14]),
    .chanx_left_in(sb_0__1__4_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__4_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__4_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__4_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__4_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__4_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__4_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__4_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__4_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__4_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__4_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__4_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__4_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__4_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__4_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__4_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__4_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__4_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__4_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__4_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__4_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__4_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[31]),
    .prog_clk_0_W_out(prog_clk_0_wires[30]),
    .pReset_S_out(pResetWires[308]),
    .pReset_E_in(pResetWires[307]),
    .pReset_W_out(pResetWires[306]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[5]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[5]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[5]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[5]),
    .SC_OUT_BOT(scff_Wires[13]),
    .SC_IN_TOP(scff_Wires[12]),
    .chanx_left_in(sb_0__1__5_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__5_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__5_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__5_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__5_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__5_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__5_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__5_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__5_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__5_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__5_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__5_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__5_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__5_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__5_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__5_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__5_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__5_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__5_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__5_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__5_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__5_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__7_
  (
    .clk_1_S_out(clk_1_wires[25]),
    .clk_1_N_out(clk_1_wires[24]),
    .clk_1_E_in(clk_1_wires[23]),
    .prog_clk_1_S_out(prog_clk_1_wires[25]),
    .prog_clk_1_N_out(prog_clk_1_wires[24]),
    .prog_clk_1_E_in(prog_clk_1_wires[23]),
    .prog_clk_0_N_in(prog_clk_0_wires[36]),
    .prog_clk_0_W_out(prog_clk_0_wires[35]),
    .pReset_S_out(pResetWires[357]),
    .pReset_E_in(pResetWires[356]),
    .pReset_W_out(pResetWires[355]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[6]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[6]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[6]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[6]),
    .SC_OUT_BOT(scff_Wires[11]),
    .SC_IN_TOP(scff_Wires[10]),
    .chanx_left_in(sb_0__1__6_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__6_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__6_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__6_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__6_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__6_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__6_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__6_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__6_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__6_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__6_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__6_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__6_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__6_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__6_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__6_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__6_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__6_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__6_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__6_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__6_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__6_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[41]),
    .prog_clk_0_W_out(prog_clk_0_wires[40]),
    .pReset_S_out(pResetWires[406]),
    .pReset_E_in(pResetWires[405]),
    .pReset_W_out(pResetWires[404]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[7]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[7]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[7]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[7]),
    .SC_OUT_BOT(scff_Wires[9]),
    .SC_IN_TOP(scff_Wires[8]),
    .chanx_left_in(sb_0__1__7_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__7_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__7_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__7_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__7_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__7_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__7_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__7_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__7_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__7_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__7_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__7_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__7_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__7_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__7_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__7_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__7_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__7_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__7_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__7_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__7_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__7_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__9_
  (
    .clk_1_S_out(clk_1_wires[32]),
    .clk_1_N_out(clk_1_wires[31]),
    .clk_1_E_in(clk_1_wires[30]),
    .prog_clk_1_S_out(prog_clk_1_wires[32]),
    .prog_clk_1_N_out(prog_clk_1_wires[31]),
    .prog_clk_1_E_in(prog_clk_1_wires[30]),
    .prog_clk_0_N_in(prog_clk_0_wires[46]),
    .prog_clk_0_W_out(prog_clk_0_wires[45]),
    .pReset_S_out(pResetWires[455]),
    .pReset_E_in(pResetWires[454]),
    .pReset_W_out(pResetWires[453]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[8]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[8]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[8]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[8]),
    .SC_OUT_BOT(scff_Wires[7]),
    .SC_IN_TOP(scff_Wires[6]),
    .chanx_left_in(sb_0__1__8_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__8_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__8_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__8_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__8_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__8_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__8_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__8_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__8_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__8_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__8_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__8_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__8_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__8_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__8_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__8_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__8_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__8_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__8_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__8_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__8_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__8_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[51]),
    .prog_clk_0_W_out(prog_clk_0_wires[50]),
    .pReset_S_out(pResetWires[504]),
    .pReset_E_in(pResetWires[503]),
    .pReset_W_out(pResetWires[502]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[9]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[9]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[9]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[9]),
    .SC_OUT_BOT(scff_Wires[5]),
    .SC_IN_TOP(scff_Wires[4]),
    .chanx_left_in(sb_0__1__9_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__9_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__9_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__9_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__9_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__9_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__9_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__9_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__9_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__9_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__9_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__9_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__9_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__9_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__9_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__9_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__9_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__9_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__9_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__9_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__9_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__9_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__11_
  (
    .clk_1_S_out(clk_1_wires[39]),
    .clk_1_N_out(clk_1_wires[38]),
    .clk_1_E_in(clk_1_wires[37]),
    .prog_clk_1_S_out(prog_clk_1_wires[39]),
    .prog_clk_1_N_out(prog_clk_1_wires[38]),
    .prog_clk_1_E_in(prog_clk_1_wires[37]),
    .prog_clk_0_N_in(prog_clk_0_wires[56]),
    .prog_clk_0_W_out(prog_clk_0_wires[55]),
    .pReset_S_out(pResetWires[553]),
    .pReset_E_in(pResetWires[552]),
    .pReset_W_out(pResetWires[551]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[10]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[10]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[10]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[10]),
    .SC_OUT_BOT(scff_Wires[3]),
    .SC_IN_TOP(scff_Wires[2]),
    .chanx_left_in(sb_0__1__10_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__10_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__10_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__10_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__10_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__10_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__10_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__10_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__10_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__10_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__10_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__10_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__10_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__10_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__10_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__10_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__10_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__10_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__10_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__10_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__10_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__10_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__1_
  (
    .clk_1_S_out(clk_1_wires[6]),
    .clk_1_N_out(clk_1_wires[5]),
    .clk_1_W_in(clk_1_wires[1]),
    .prog_clk_1_S_out(prog_clk_1_wires[6]),
    .prog_clk_1_N_out(prog_clk_1_wires[5]),
    .prog_clk_1_W_in(prog_clk_1_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[66]),
    .pReset_S_out(pResetWires[68]),
    .pReset_E_in(pResetWires[67]),
    .pReset_W_out(pResetWires[66]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[11]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[11]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[11]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[11]),
    .SC_OUT_TOP(scff_Wires[30]),
    .SC_IN_BOT(scff_Wires[29]),
    .chanx_left_in(sb_1__1__0_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__11_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__11_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__11_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__11_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__11_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__11_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__11_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__11_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__11_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__11_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__11_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__11_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__11_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__11_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__11_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__11_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__11_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__11_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__11_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__11_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__11_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__2_
  (
    .clk_2_E_in(clk_2_wires[2]),
    .clk_2_W_out(clk_2_wires[1]),
    .prog_clk_2_E_in(prog_clk_2_wires[2]),
    .prog_clk_2_W_out(prog_clk_2_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[69]),
    .pReset_S_out(pResetWires[117]),
    .pReset_E_in(pResetWires[116]),
    .pReset_W_out(pResetWires[115]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[12]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[12]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[12]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[12]),
    .SC_OUT_TOP(scff_Wires[32]),
    .SC_IN_BOT(scff_Wires[31]),
    .chanx_left_in(sb_1__1__1_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__12_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__12_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__12_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__12_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__12_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__12_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__12_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__12_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__12_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__12_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__12_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__12_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__12_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__12_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__12_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__12_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__12_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__12_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__12_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__12_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__12_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__3_
  (
    .clk_1_S_out(clk_1_wires[13]),
    .clk_1_N_out(clk_1_wires[12]),
    .clk_1_W_in(clk_1_wires[8]),
    .prog_clk_1_S_out(prog_clk_1_wires[13]),
    .prog_clk_1_N_out(prog_clk_1_wires[12]),
    .prog_clk_1_W_in(prog_clk_1_wires[8]),
    .prog_clk_0_N_in(prog_clk_0_wires[72]),
    .pReset_S_out(pResetWires[166]),
    .pReset_E_in(pResetWires[165]),
    .pReset_W_out(pResetWires[164]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[13]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[13]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[13]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[13]),
    .SC_OUT_TOP(scff_Wires[34]),
    .SC_IN_BOT(scff_Wires[33]),
    .chanx_left_in(sb_1__1__2_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__13_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__13_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__13_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__13_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__13_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__13_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__13_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__13_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__13_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__13_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__13_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__13_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__13_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__13_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__13_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__13_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__13_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__13_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__13_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__13_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__13_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__4_
  (
    .clk_2_E_in(clk_2_wires[7]),
    .clk_2_W_out(clk_2_wires[6]),
    .prog_clk_2_E_in(prog_clk_2_wires[7]),
    .prog_clk_2_W_out(prog_clk_2_wires[6]),
    .prog_clk_0_N_in(prog_clk_0_wires[75]),
    .pReset_S_out(pResetWires[215]),
    .pReset_E_in(pResetWires[214]),
    .pReset_W_out(pResetWires[213]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[14]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[14]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[14]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[14]),
    .SC_OUT_TOP(scff_Wires[36]),
    .SC_IN_BOT(scff_Wires[35]),
    .chanx_left_in(sb_1__1__3_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__14_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__14_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__14_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__14_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__14_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__14_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__14_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__14_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__14_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__14_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__14_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__14_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__14_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__14_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__14_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__14_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__14_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__14_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__14_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__14_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__14_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__5_
  (
    .clk_1_S_out(clk_1_wires[20]),
    .clk_1_N_out(clk_1_wires[19]),
    .clk_1_W_in(clk_1_wires[15]),
    .prog_clk_1_S_out(prog_clk_1_wires[20]),
    .prog_clk_1_N_out(prog_clk_1_wires[19]),
    .prog_clk_1_W_in(prog_clk_1_wires[15]),
    .prog_clk_0_N_in(prog_clk_0_wires[78]),
    .pReset_S_out(pResetWires[264]),
    .pReset_E_in(pResetWires[263]),
    .pReset_W_out(pResetWires[262]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[15]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[15]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[15]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[15]),
    .SC_OUT_TOP(scff_Wires[38]),
    .SC_IN_BOT(scff_Wires[37]),
    .chanx_left_in(sb_1__1__4_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__15_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__15_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__15_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__15_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__15_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__15_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__15_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__15_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__15_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__15_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__15_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__15_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__15_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__15_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__15_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__15_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__15_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__15_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__15_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__15_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__15_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[81]),
    .pReset_S_out(pResetWires[313]),
    .pReset_E_in(pResetWires[312]),
    .pReset_W_out(pResetWires[311]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[16]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[16]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[16]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[16]),
    .SC_OUT_TOP(scff_Wires[40]),
    .SC_IN_BOT(scff_Wires[39]),
    .chanx_left_in(sb_1__1__5_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__16_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__16_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__16_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__16_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__16_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__16_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__16_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__16_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__16_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__16_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__16_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__16_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__16_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__16_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__16_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__16_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__16_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__16_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__16_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__16_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__16_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__7_
  (
    .clk_1_S_out(clk_1_wires[27]),
    .clk_1_N_out(clk_1_wires[26]),
    .clk_1_W_in(clk_1_wires[22]),
    .prog_clk_1_S_out(prog_clk_1_wires[27]),
    .prog_clk_1_N_out(prog_clk_1_wires[26]),
    .prog_clk_1_W_in(prog_clk_1_wires[22]),
    .prog_clk_0_N_in(prog_clk_0_wires[84]),
    .pReset_S_out(pResetWires[362]),
    .pReset_E_in(pResetWires[361]),
    .pReset_W_out(pResetWires[360]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[17]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[17]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[17]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[17]),
    .SC_OUT_TOP(scff_Wires[42]),
    .SC_IN_BOT(scff_Wires[41]),
    .chanx_left_in(sb_1__1__6_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__17_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__17_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__17_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__17_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__17_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__17_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__17_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__17_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__17_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__17_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__17_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__17_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__17_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__17_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__17_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__17_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__17_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__17_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__17_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__17_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__17_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__8_
  (
    .clk_2_E_in(clk_2_wires[14]),
    .clk_2_W_out(clk_2_wires[13]),
    .prog_clk_2_E_in(prog_clk_2_wires[14]),
    .prog_clk_2_W_out(prog_clk_2_wires[13]),
    .prog_clk_0_N_in(prog_clk_0_wires[87]),
    .pReset_S_out(pResetWires[411]),
    .pReset_E_in(pResetWires[410]),
    .pReset_W_out(pResetWires[409]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[18]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[18]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[18]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[18]),
    .SC_OUT_TOP(scff_Wires[44]),
    .SC_IN_BOT(scff_Wires[43]),
    .chanx_left_in(sb_1__1__7_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__18_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__18_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__18_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__18_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__18_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__18_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__18_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__18_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__18_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__18_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__18_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__18_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__18_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__18_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__18_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__18_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__18_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__18_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__18_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__18_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__18_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__9_
  (
    .clk_1_S_out(clk_1_wires[34]),
    .clk_1_N_out(clk_1_wires[33]),
    .clk_1_W_in(clk_1_wires[29]),
    .prog_clk_1_S_out(prog_clk_1_wires[34]),
    .prog_clk_1_N_out(prog_clk_1_wires[33]),
    .prog_clk_1_W_in(prog_clk_1_wires[29]),
    .prog_clk_0_N_in(prog_clk_0_wires[90]),
    .pReset_S_out(pResetWires[460]),
    .pReset_E_in(pResetWires[459]),
    .pReset_W_out(pResetWires[458]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[19]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[19]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[19]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[19]),
    .SC_OUT_TOP(scff_Wires[46]),
    .SC_IN_BOT(scff_Wires[45]),
    .chanx_left_in(sb_1__1__8_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__19_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__19_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__19_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__19_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__19_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__19_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__19_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__19_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__19_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__19_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__19_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__19_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__19_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__19_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__19_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__19_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__19_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__19_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__19_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__19_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__19_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__10_
  (
    .clk_2_E_in(clk_2_wires[21]),
    .clk_2_W_out(clk_2_wires[20]),
    .prog_clk_2_E_in(prog_clk_2_wires[21]),
    .prog_clk_2_W_out(prog_clk_2_wires[20]),
    .prog_clk_0_N_in(prog_clk_0_wires[93]),
    .pReset_S_out(pResetWires[509]),
    .pReset_E_in(pResetWires[508]),
    .pReset_W_out(pResetWires[507]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[20]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[20]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[20]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[20]),
    .SC_OUT_TOP(scff_Wires[48]),
    .SC_IN_BOT(scff_Wires[47]),
    .chanx_left_in(sb_1__1__9_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__20_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__20_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__20_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__20_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__20_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__20_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__20_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__20_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__20_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__20_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__20_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__20_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__20_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__20_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__20_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__20_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__20_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__20_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__20_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__20_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__20_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__11_
  (
    .clk_1_S_out(clk_1_wires[41]),
    .clk_1_N_out(clk_1_wires[40]),
    .clk_1_W_in(clk_1_wires[36]),
    .prog_clk_1_S_out(prog_clk_1_wires[41]),
    .prog_clk_1_N_out(prog_clk_1_wires[40]),
    .prog_clk_1_W_in(prog_clk_1_wires[36]),
    .prog_clk_0_N_in(prog_clk_0_wires[96]),
    .pReset_S_out(pResetWires[558]),
    .pReset_E_in(pResetWires[557]),
    .pReset_W_out(pResetWires[556]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[21]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[21]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[21]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[21]),
    .SC_OUT_TOP(scff_Wires[50]),
    .SC_IN_BOT(scff_Wires[49]),
    .chanx_left_in(sb_1__1__10_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__21_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__21_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__21_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__21_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__21_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__21_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__21_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__21_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__21_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__21_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__21_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__21_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__21_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__21_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__21_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__21_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__21_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__21_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__21_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__21_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__21_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__1_
  (
    .clk_1_S_out(clk_1_wires[46]),
    .clk_1_N_out(clk_1_wires[45]),
    .clk_1_E_in(clk_1_wires[44]),
    .prog_clk_1_S_out(prog_clk_1_wires[46]),
    .prog_clk_1_N_out(prog_clk_1_wires[45]),
    .prog_clk_1_E_in(prog_clk_1_wires[44]),
    .prog_clk_0_N_in(prog_clk_0_wires[104]),
    .pReset_S_out(pResetWires[72]),
    .pReset_E_in(pResetWires[71]),
    .pReset_W_out(pResetWires[70]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[22]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[22]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[22]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[22]),
    .SC_OUT_BOT(scff_Wires[76]),
    .SC_IN_TOP(scff_Wires[75]),
    .chanx_left_in(sb_1__1__11_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__22_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__22_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__22_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__22_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__22_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__22_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__22_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__22_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__22_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__22_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__22_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__22_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__22_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__22_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__22_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__22_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__22_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__22_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__22_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__22_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__22_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[107]),
    .pReset_S_out(pResetWires[121]),
    .pReset_E_in(pResetWires[120]),
    .pReset_W_out(pResetWires[119]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[23]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[23]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[23]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[23]),
    .SC_OUT_BOT(scff_Wires[74]),
    .SC_IN_TOP(scff_Wires[73]),
    .chanx_left_in(sb_1__1__12_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__23_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__23_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__23_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__23_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__23_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__23_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__23_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__23_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__23_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__23_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__23_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__23_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__23_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__23_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__23_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__23_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__23_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__23_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__23_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__23_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__23_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__3_
  (
    .clk_1_S_out(clk_1_wires[53]),
    .clk_1_N_out(clk_1_wires[52]),
    .clk_1_E_in(clk_1_wires[51]),
    .prog_clk_1_S_out(prog_clk_1_wires[53]),
    .prog_clk_1_N_out(prog_clk_1_wires[52]),
    .prog_clk_1_E_in(prog_clk_1_wires[51]),
    .prog_clk_0_N_in(prog_clk_0_wires[110]),
    .pReset_S_out(pResetWires[170]),
    .pReset_E_in(pResetWires[169]),
    .pReset_W_out(pResetWires[168]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[24]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[24]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[24]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[24]),
    .SC_OUT_BOT(scff_Wires[72]),
    .SC_IN_TOP(scff_Wires[71]),
    .chanx_left_in(sb_1__1__13_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__24_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__24_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__24_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__24_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__24_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__24_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__24_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__24_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__24_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__24_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__24_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__24_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__24_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__24_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__24_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__24_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__24_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__24_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__24_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__24_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__24_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[113]),
    .pReset_S_out(pResetWires[219]),
    .pReset_E_in(pResetWires[218]),
    .pReset_W_out(pResetWires[217]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[25]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[25]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[25]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[25]),
    .SC_OUT_BOT(scff_Wires[70]),
    .SC_IN_TOP(scff_Wires[69]),
    .chanx_left_in(sb_1__1__14_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__25_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__25_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__25_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__25_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__25_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__25_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__25_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__25_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__25_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__25_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__25_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__25_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__25_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__25_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__25_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__25_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__25_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__25_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__25_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__25_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__25_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__5_
  (
    .clk_1_S_out(clk_1_wires[60]),
    .clk_1_N_out(clk_1_wires[59]),
    .clk_1_E_in(clk_1_wires[58]),
    .prog_clk_1_S_out(prog_clk_1_wires[60]),
    .prog_clk_1_N_out(prog_clk_1_wires[59]),
    .prog_clk_1_E_in(prog_clk_1_wires[58]),
    .prog_clk_0_N_in(prog_clk_0_wires[116]),
    .pReset_S_out(pResetWires[268]),
    .pReset_E_in(pResetWires[267]),
    .pReset_W_out(pResetWires[266]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[26]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[26]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[26]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[26]),
    .SC_OUT_BOT(scff_Wires[68]),
    .SC_IN_TOP(scff_Wires[67]),
    .chanx_left_in(sb_1__1__15_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__26_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__26_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__26_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__26_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__26_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__26_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__26_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__26_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__26_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__26_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__26_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__26_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__26_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__26_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__26_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__26_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__26_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__26_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__26_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__26_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__26_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__6_
  (
    .clk_3_W_out(clk_3_wires[51]),
    .clk_3_E_in(clk_3_wires[50]),
    .prog_clk_3_W_out(prog_clk_3_wires[51]),
    .prog_clk_3_E_in(prog_clk_3_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[119]),
    .pReset_S_out(pResetWires[317]),
    .pReset_E_in(pResetWires[316]),
    .pReset_W_out(pResetWires[315]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[27]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[27]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[27]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[27]),
    .SC_OUT_BOT(scff_Wires[66]),
    .SC_IN_TOP(scff_Wires[65]),
    .chanx_left_in(sb_1__1__16_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__27_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__27_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__27_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__27_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__27_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__27_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__27_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__27_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__27_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__27_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__27_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__27_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__27_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__27_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__27_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__27_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__27_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__27_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__27_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__27_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__27_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__7_
  (
    .clk_1_S_out(clk_1_wires[67]),
    .clk_1_N_out(clk_1_wires[66]),
    .clk_1_E_in(clk_1_wires[65]),
    .prog_clk_1_S_out(prog_clk_1_wires[67]),
    .prog_clk_1_N_out(prog_clk_1_wires[66]),
    .prog_clk_1_E_in(prog_clk_1_wires[65]),
    .prog_clk_0_N_in(prog_clk_0_wires[122]),
    .pReset_S_out(pResetWires[366]),
    .pReset_E_in(pResetWires[365]),
    .pReset_W_out(pResetWires[364]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[28]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[28]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[28]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[28]),
    .SC_OUT_BOT(scff_Wires[64]),
    .SC_IN_TOP(scff_Wires[63]),
    .chanx_left_in(sb_1__1__17_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__28_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__28_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__28_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__28_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__28_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__28_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__28_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__28_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__28_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__28_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__28_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__28_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__28_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__28_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__28_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__28_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__28_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__28_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__28_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__28_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__28_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[125]),
    .pReset_S_out(pResetWires[415]),
    .pReset_E_in(pResetWires[414]),
    .pReset_W_out(pResetWires[413]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[29]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[29]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[29]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[29]),
    .SC_OUT_BOT(scff_Wires[62]),
    .SC_IN_TOP(scff_Wires[61]),
    .chanx_left_in(sb_1__1__18_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__29_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__29_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__29_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__29_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__29_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__29_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__29_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__29_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__29_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__29_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__29_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__29_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__29_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__29_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__29_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__29_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__29_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__29_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__29_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__29_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__29_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__9_
  (
    .clk_1_S_out(clk_1_wires[74]),
    .clk_1_N_out(clk_1_wires[73]),
    .clk_1_E_in(clk_1_wires[72]),
    .prog_clk_1_S_out(prog_clk_1_wires[74]),
    .prog_clk_1_N_out(prog_clk_1_wires[73]),
    .prog_clk_1_E_in(prog_clk_1_wires[72]),
    .prog_clk_0_N_in(prog_clk_0_wires[128]),
    .pReset_S_out(pResetWires[464]),
    .pReset_E_in(pResetWires[463]),
    .pReset_W_out(pResetWires[462]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[30]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[30]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[30]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[30]),
    .SC_OUT_BOT(scff_Wires[60]),
    .SC_IN_TOP(scff_Wires[59]),
    .chanx_left_in(sb_1__1__19_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__30_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__30_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__30_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__30_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__30_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__30_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__30_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__30_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__30_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__30_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__30_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__30_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__30_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__30_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__30_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__30_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__30_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__30_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__30_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__30_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__30_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[131]),
    .pReset_S_out(pResetWires[513]),
    .pReset_E_in(pResetWires[512]),
    .pReset_W_out(pResetWires[511]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[31]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[31]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[31]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[31]),
    .SC_OUT_BOT(scff_Wires[58]),
    .SC_IN_TOP(scff_Wires[57]),
    .chanx_left_in(sb_1__1__20_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__31_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__31_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__31_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__31_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__31_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__31_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__31_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__31_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__31_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__31_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__31_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__31_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__31_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__31_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__31_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__31_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__31_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__31_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__31_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__31_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__31_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__11_
  (
    .clk_1_S_out(clk_1_wires[81]),
    .clk_1_N_out(clk_1_wires[80]),
    .clk_1_E_in(clk_1_wires[79]),
    .prog_clk_1_S_out(prog_clk_1_wires[81]),
    .prog_clk_1_N_out(prog_clk_1_wires[80]),
    .prog_clk_1_E_in(prog_clk_1_wires[79]),
    .prog_clk_0_N_in(prog_clk_0_wires[134]),
    .pReset_S_out(pResetWires[562]),
    .pReset_E_in(pResetWires[561]),
    .pReset_W_out(pResetWires[560]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[32]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[32]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[32]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[32]),
    .SC_OUT_BOT(scff_Wires[56]),
    .SC_IN_TOP(scff_Wires[55]),
    .chanx_left_in(sb_1__1__21_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__32_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__32_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__32_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__32_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__32_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__32_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__32_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__32_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__32_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__32_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__32_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__32_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__32_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__32_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__32_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__32_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__32_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__32_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__32_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__32_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__32_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__1_
  (
    .clk_1_S_out(clk_1_wires[48]),
    .clk_1_N_out(clk_1_wires[47]),
    .clk_1_W_in(clk_1_wires[43]),
    .prog_clk_1_S_out(prog_clk_1_wires[48]),
    .prog_clk_1_N_out(prog_clk_1_wires[47]),
    .prog_clk_1_W_in(prog_clk_1_wires[43]),
    .prog_clk_0_N_in(prog_clk_0_wires[142]),
    .pReset_S_out(pResetWires[76]),
    .pReset_E_in(pResetWires[75]),
    .pReset_W_out(pResetWires[74]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[33]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[33]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[33]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[33]),
    .SC_OUT_TOP(scff_Wires[83]),
    .SC_IN_BOT(scff_Wires[82]),
    .chanx_left_in(sb_1__1__22_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__33_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__33_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__33_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__33_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__33_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__33_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__33_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__33_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__33_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__33_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__33_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__33_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__33_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__33_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__33_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__33_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__33_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__33_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__33_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__33_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__33_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__2_
  (
    .clk_2_W_out(clk_2_wires[28]),
    .clk_2_E_in(clk_2_wires[27]),
    .prog_clk_2_W_out(prog_clk_2_wires[28]),
    .prog_clk_2_E_in(prog_clk_2_wires[27]),
    .prog_clk_0_N_in(prog_clk_0_wires[145]),
    .pReset_S_out(pResetWires[125]),
    .pReset_E_in(pResetWires[124]),
    .pReset_W_out(pResetWires[123]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[34]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[34]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[34]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[34]),
    .SC_OUT_TOP(scff_Wires[85]),
    .SC_IN_BOT(scff_Wires[84]),
    .chanx_left_in(sb_1__1__23_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__34_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__34_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__34_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__34_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__34_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__34_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__34_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__34_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__34_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__34_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__34_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__34_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__34_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__34_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__34_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__34_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__34_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__34_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__34_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__34_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__34_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__3_
  (
    .clk_1_S_out(clk_1_wires[55]),
    .clk_1_N_out(clk_1_wires[54]),
    .clk_1_W_in(clk_1_wires[50]),
    .prog_clk_1_S_out(prog_clk_1_wires[55]),
    .prog_clk_1_N_out(prog_clk_1_wires[54]),
    .prog_clk_1_W_in(prog_clk_1_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[148]),
    .pReset_S_out(pResetWires[174]),
    .pReset_E_in(pResetWires[173]),
    .pReset_W_out(pResetWires[172]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[35]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[35]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[35]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[35]),
    .SC_OUT_TOP(scff_Wires[87]),
    .SC_IN_BOT(scff_Wires[86]),
    .chanx_left_in(sb_1__1__24_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__35_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__35_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__35_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__35_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__35_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__35_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__35_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__35_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__35_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__35_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__35_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__35_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__35_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__35_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__35_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__35_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__35_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__35_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__35_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__35_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__35_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__4_
  (
    .clk_2_W_out(clk_2_wires[37]),
    .clk_2_E_in(clk_2_wires[36]),
    .prog_clk_2_W_out(prog_clk_2_wires[37]),
    .prog_clk_2_E_in(prog_clk_2_wires[36]),
    .prog_clk_0_N_in(prog_clk_0_wires[151]),
    .pReset_S_out(pResetWires[223]),
    .pReset_E_in(pResetWires[222]),
    .pReset_W_out(pResetWires[221]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[36]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[36]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[36]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[36]),
    .SC_OUT_TOP(scff_Wires[89]),
    .SC_IN_BOT(scff_Wires[88]),
    .chanx_left_in(sb_1__1__25_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__36_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__36_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__36_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__36_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__36_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__36_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__36_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__36_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__36_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__36_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__36_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__36_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__36_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__36_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__36_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__36_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__36_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__36_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__36_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__36_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__36_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__5_
  (
    .clk_1_S_out(clk_1_wires[62]),
    .clk_1_N_out(clk_1_wires[61]),
    .clk_1_W_in(clk_1_wires[57]),
    .prog_clk_1_S_out(prog_clk_1_wires[62]),
    .prog_clk_1_N_out(prog_clk_1_wires[61]),
    .prog_clk_1_W_in(prog_clk_1_wires[57]),
    .prog_clk_0_N_in(prog_clk_0_wires[154]),
    .pReset_S_out(pResetWires[272]),
    .pReset_E_in(pResetWires[271]),
    .pReset_W_out(pResetWires[270]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[37]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[37]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[37]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[37]),
    .SC_OUT_TOP(scff_Wires[91]),
    .SC_IN_BOT(scff_Wires[90]),
    .chanx_left_in(sb_1__1__26_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__37_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__37_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__37_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__37_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__37_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__37_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__37_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__37_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__37_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__37_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__37_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__37_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__37_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__37_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__37_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__37_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__37_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__37_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__37_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__37_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__37_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__6_
  (
    .clk_3_W_out(clk_3_wires[47]),
    .clk_3_E_in(clk_3_wires[46]),
    .prog_clk_3_W_out(prog_clk_3_wires[47]),
    .prog_clk_3_E_in(prog_clk_3_wires[46]),
    .prog_clk_0_N_in(prog_clk_0_wires[157]),
    .pReset_S_out(pResetWires[321]),
    .pReset_E_in(pResetWires[320]),
    .pReset_W_out(pResetWires[319]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[38]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[38]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[38]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[38]),
    .SC_OUT_TOP(scff_Wires[93]),
    .SC_IN_BOT(scff_Wires[92]),
    .chanx_left_in(sb_1__1__27_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__38_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__38_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__38_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__38_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__38_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__38_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__38_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__38_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__38_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__38_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__38_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__38_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__38_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__38_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__38_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__38_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__38_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__38_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__38_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__38_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__38_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__7_
  (
    .clk_1_S_out(clk_1_wires[69]),
    .clk_1_N_out(clk_1_wires[68]),
    .clk_1_W_in(clk_1_wires[64]),
    .prog_clk_1_S_out(prog_clk_1_wires[69]),
    .prog_clk_1_N_out(prog_clk_1_wires[68]),
    .prog_clk_1_W_in(prog_clk_1_wires[64]),
    .prog_clk_0_N_in(prog_clk_0_wires[160]),
    .pReset_S_out(pResetWires[370]),
    .pReset_E_in(pResetWires[369]),
    .pReset_W_out(pResetWires[368]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[39]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[39]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[39]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[39]),
    .SC_OUT_TOP(scff_Wires[95]),
    .SC_IN_BOT(scff_Wires[94]),
    .chanx_left_in(sb_1__1__28_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__39_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__39_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__39_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__39_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__39_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__39_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__39_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__39_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__39_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__39_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__39_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__39_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__39_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__39_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__39_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__39_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__39_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__39_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__39_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__39_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__39_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__8_
  (
    .clk_2_W_out(clk_2_wires[50]),
    .clk_2_E_in(clk_2_wires[49]),
    .prog_clk_2_W_out(prog_clk_2_wires[50]),
    .prog_clk_2_E_in(prog_clk_2_wires[49]),
    .prog_clk_0_N_in(prog_clk_0_wires[163]),
    .pReset_S_out(pResetWires[419]),
    .pReset_E_in(pResetWires[418]),
    .pReset_W_out(pResetWires[417]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[40]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[40]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[40]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[40]),
    .SC_OUT_TOP(scff_Wires[97]),
    .SC_IN_BOT(scff_Wires[96]),
    .chanx_left_in(sb_1__1__29_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__40_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__40_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__40_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__40_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__40_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__40_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__40_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__40_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__40_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__40_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__40_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__40_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__40_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__40_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__40_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__40_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__40_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__40_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__40_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__40_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__40_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__9_
  (
    .clk_1_S_out(clk_1_wires[76]),
    .clk_1_N_out(clk_1_wires[75]),
    .clk_1_W_in(clk_1_wires[71]),
    .prog_clk_1_S_out(prog_clk_1_wires[76]),
    .prog_clk_1_N_out(prog_clk_1_wires[75]),
    .prog_clk_1_W_in(prog_clk_1_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[166]),
    .pReset_S_out(pResetWires[468]),
    .pReset_E_in(pResetWires[467]),
    .pReset_W_out(pResetWires[466]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[41]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[41]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[41]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[41]),
    .SC_OUT_TOP(scff_Wires[99]),
    .SC_IN_BOT(scff_Wires[98]),
    .chanx_left_in(sb_1__1__30_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__41_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__41_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__41_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__41_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__41_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__41_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__41_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__41_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__41_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__41_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__41_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__41_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__41_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__41_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__41_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__41_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__41_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__41_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__41_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__41_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__41_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__10_
  (
    .clk_2_W_out(clk_2_wires[63]),
    .clk_2_E_in(clk_2_wires[62]),
    .prog_clk_2_W_out(prog_clk_2_wires[63]),
    .prog_clk_2_E_in(prog_clk_2_wires[62]),
    .prog_clk_0_N_in(prog_clk_0_wires[169]),
    .pReset_S_out(pResetWires[517]),
    .pReset_E_in(pResetWires[516]),
    .pReset_W_out(pResetWires[515]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[42]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[42]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[42]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[42]),
    .SC_OUT_TOP(scff_Wires[101]),
    .SC_IN_BOT(scff_Wires[100]),
    .chanx_left_in(sb_1__1__31_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__42_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__42_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__42_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__42_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__42_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__42_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__42_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__42_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__42_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__42_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__42_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__42_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__42_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__42_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__42_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__42_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__42_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__42_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__42_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__42_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__42_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__11_
  (
    .clk_1_S_out(clk_1_wires[83]),
    .clk_1_N_out(clk_1_wires[82]),
    .clk_1_W_in(clk_1_wires[78]),
    .prog_clk_1_S_out(prog_clk_1_wires[83]),
    .prog_clk_1_N_out(prog_clk_1_wires[82]),
    .prog_clk_1_W_in(prog_clk_1_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[172]),
    .pReset_S_out(pResetWires[566]),
    .pReset_E_in(pResetWires[565]),
    .pReset_W_out(pResetWires[564]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[43]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[43]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[43]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[43]),
    .SC_OUT_TOP(scff_Wires[103]),
    .SC_IN_BOT(scff_Wires[102]),
    .chanx_left_in(sb_1__1__32_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__43_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__43_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__43_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__43_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__43_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__43_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__43_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__43_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__43_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__43_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__43_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__43_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__43_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__43_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__43_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__43_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__43_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__43_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__43_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__43_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__43_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__1_
  (
    .clk_1_S_out(clk_1_wires[88]),
    .clk_1_N_out(clk_1_wires[87]),
    .clk_1_E_in(clk_1_wires[86]),
    .prog_clk_1_S_out(prog_clk_1_wires[88]),
    .prog_clk_1_N_out(prog_clk_1_wires[87]),
    .prog_clk_1_E_in(prog_clk_1_wires[86]),
    .prog_clk_0_N_in(prog_clk_0_wires[180]),
    .pReset_S_out(pResetWires[80]),
    .pReset_E_in(pResetWires[79]),
    .pReset_W_out(pResetWires[78]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[44]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[44]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[44]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[44]),
    .SC_OUT_BOT(scff_Wires[129]),
    .SC_IN_TOP(scff_Wires[128]),
    .chanx_left_in(sb_1__1__33_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__44_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__44_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__44_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__44_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__44_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__44_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__44_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__44_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__44_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__44_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__44_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__44_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__44_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__44_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__44_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__44_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__44_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__44_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__44_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__44_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__44_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__2_
  (
    .clk_2_E_out(clk_2_wires[26]),
    .clk_2_W_in(clk_2_wires[25]),
    .prog_clk_2_E_out(prog_clk_2_wires[26]),
    .prog_clk_2_W_in(prog_clk_2_wires[25]),
    .prog_clk_0_N_in(prog_clk_0_wires[183]),
    .pReset_S_out(pResetWires[129]),
    .pReset_E_in(pResetWires[128]),
    .pReset_W_out(pResetWires[127]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[45]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[45]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[45]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[45]),
    .SC_OUT_BOT(scff_Wires[127]),
    .SC_IN_TOP(scff_Wires[126]),
    .chanx_left_in(sb_1__1__34_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__45_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__45_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__45_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__45_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__45_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__45_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__45_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__45_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__45_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__45_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__45_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__45_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__45_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__45_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__45_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__45_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__45_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__45_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__45_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__45_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__45_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__3_
  (
    .clk_1_S_out(clk_1_wires[95]),
    .clk_1_N_out(clk_1_wires[94]),
    .clk_1_E_in(clk_1_wires[93]),
    .prog_clk_1_S_out(prog_clk_1_wires[95]),
    .prog_clk_1_N_out(prog_clk_1_wires[94]),
    .prog_clk_1_E_in(prog_clk_1_wires[93]),
    .prog_clk_0_N_in(prog_clk_0_wires[186]),
    .pReset_S_out(pResetWires[178]),
    .pReset_E_in(pResetWires[177]),
    .pReset_W_out(pResetWires[176]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[46]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[46]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[46]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[46]),
    .SC_OUT_BOT(scff_Wires[125]),
    .SC_IN_TOP(scff_Wires[124]),
    .chanx_left_in(sb_1__1__35_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__46_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__46_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__46_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__46_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__46_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__46_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__46_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__46_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__46_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__46_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__46_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__46_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__46_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__46_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__46_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__46_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__46_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__46_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__46_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__46_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__46_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__4_
  (
    .clk_2_E_out(clk_2_wires[35]),
    .clk_2_W_in(clk_2_wires[34]),
    .prog_clk_2_E_out(prog_clk_2_wires[35]),
    .prog_clk_2_W_in(prog_clk_2_wires[34]),
    .prog_clk_0_N_in(prog_clk_0_wires[189]),
    .pReset_S_out(pResetWires[227]),
    .pReset_E_in(pResetWires[226]),
    .pReset_W_out(pResetWires[225]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[47]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[47]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[47]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[47]),
    .SC_OUT_BOT(scff_Wires[123]),
    .SC_IN_TOP(scff_Wires[122]),
    .chanx_left_in(sb_1__1__36_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__47_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__47_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__47_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__47_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__47_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__47_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__47_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__47_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__47_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__47_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__47_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__47_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__47_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__47_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__47_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__47_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__47_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__47_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__47_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__47_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__47_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__5_
  (
    .clk_1_S_out(clk_1_wires[102]),
    .clk_1_N_out(clk_1_wires[101]),
    .clk_1_E_in(clk_1_wires[100]),
    .prog_clk_1_S_out(prog_clk_1_wires[102]),
    .prog_clk_1_N_out(prog_clk_1_wires[101]),
    .prog_clk_1_E_in(prog_clk_1_wires[100]),
    .prog_clk_0_N_in(prog_clk_0_wires[192]),
    .pReset_S_out(pResetWires[276]),
    .pReset_E_in(pResetWires[275]),
    .pReset_W_out(pResetWires[274]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[48]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[48]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[48]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[48]),
    .SC_OUT_BOT(scff_Wires[121]),
    .SC_IN_TOP(scff_Wires[120]),
    .chanx_left_in(sb_1__1__37_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__48_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__48_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__48_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__48_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__48_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__48_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__48_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__48_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__48_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__48_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__48_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__48_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__48_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__48_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__48_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__48_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__48_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__48_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__48_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__48_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__48_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__6_
  (
    .clk_3_W_out(clk_3_wires[7]),
    .clk_3_E_in(clk_3_wires[6]),
    .prog_clk_3_W_out(prog_clk_3_wires[7]),
    .prog_clk_3_E_in(prog_clk_3_wires[6]),
    .prog_clk_0_N_in(prog_clk_0_wires[195]),
    .pReset_S_out(pResetWires[325]),
    .pReset_E_in(pResetWires[324]),
    .pReset_W_out(pResetWires[323]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[49]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[49]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[49]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[49]),
    .SC_OUT_BOT(scff_Wires[119]),
    .SC_IN_TOP(scff_Wires[118]),
    .chanx_left_in(sb_1__1__38_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__49_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__49_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__49_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__49_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__49_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__49_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__49_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__49_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__49_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__49_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__49_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__49_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__49_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__49_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__49_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__49_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__49_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__49_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__49_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__49_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__49_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__7_
  (
    .clk_1_S_out(clk_1_wires[109]),
    .clk_1_N_out(clk_1_wires[108]),
    .clk_1_E_in(clk_1_wires[107]),
    .prog_clk_1_S_out(prog_clk_1_wires[109]),
    .prog_clk_1_N_out(prog_clk_1_wires[108]),
    .prog_clk_1_E_in(prog_clk_1_wires[107]),
    .prog_clk_0_N_in(prog_clk_0_wires[198]),
    .pReset_S_out(pResetWires[374]),
    .pReset_E_in(pResetWires[373]),
    .pReset_W_out(pResetWires[372]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[50]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[50]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[50]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[50]),
    .SC_OUT_BOT(scff_Wires[117]),
    .SC_IN_TOP(scff_Wires[116]),
    .chanx_left_in(sb_1__1__39_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__50_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__50_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__50_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__50_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__50_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__50_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__50_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__50_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__50_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__50_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__50_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__50_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__50_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__50_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__50_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__50_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__50_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__50_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__50_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__50_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__50_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__8_
  (
    .clk_2_E_out(clk_2_wires[48]),
    .clk_2_W_in(clk_2_wires[47]),
    .prog_clk_2_E_out(prog_clk_2_wires[48]),
    .prog_clk_2_W_in(prog_clk_2_wires[47]),
    .prog_clk_0_N_in(prog_clk_0_wires[201]),
    .pReset_S_out(pResetWires[423]),
    .pReset_E_in(pResetWires[422]),
    .pReset_W_out(pResetWires[421]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[51]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[51]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[51]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[51]),
    .SC_OUT_BOT(scff_Wires[115]),
    .SC_IN_TOP(scff_Wires[114]),
    .chanx_left_in(sb_1__1__40_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__51_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__51_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__51_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__51_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__51_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__51_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__51_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__51_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__51_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__51_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__51_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__51_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__51_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__51_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__51_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__51_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__51_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__51_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__51_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__51_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__51_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__9_
  (
    .clk_1_S_out(clk_1_wires[116]),
    .clk_1_N_out(clk_1_wires[115]),
    .clk_1_E_in(clk_1_wires[114]),
    .prog_clk_1_S_out(prog_clk_1_wires[116]),
    .prog_clk_1_N_out(prog_clk_1_wires[115]),
    .prog_clk_1_E_in(prog_clk_1_wires[114]),
    .prog_clk_0_N_in(prog_clk_0_wires[204]),
    .pReset_S_out(pResetWires[472]),
    .pReset_E_in(pResetWires[471]),
    .pReset_W_out(pResetWires[470]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[52]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[52]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[52]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[52]),
    .SC_OUT_BOT(scff_Wires[113]),
    .SC_IN_TOP(scff_Wires[112]),
    .chanx_left_in(sb_1__1__41_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__52_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__52_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__52_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__52_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__52_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__52_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__52_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__52_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__52_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__52_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__52_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__52_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__52_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__52_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__52_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__52_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__52_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__52_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__52_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__52_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__52_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__10_
  (
    .clk_2_E_out(clk_2_wires[61]),
    .clk_2_W_in(clk_2_wires[60]),
    .prog_clk_2_E_out(prog_clk_2_wires[61]),
    .prog_clk_2_W_in(prog_clk_2_wires[60]),
    .prog_clk_0_N_in(prog_clk_0_wires[207]),
    .pReset_S_out(pResetWires[521]),
    .pReset_E_in(pResetWires[520]),
    .pReset_W_out(pResetWires[519]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[53]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[53]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[53]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[53]),
    .SC_OUT_BOT(scff_Wires[111]),
    .SC_IN_TOP(scff_Wires[110]),
    .chanx_left_in(sb_1__1__42_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__53_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__53_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__53_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__53_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__53_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__53_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__53_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__53_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__53_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__53_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__53_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__53_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__53_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__53_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__53_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__53_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__53_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__53_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__53_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__53_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__53_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__11_
  (
    .clk_1_S_out(clk_1_wires[123]),
    .clk_1_N_out(clk_1_wires[122]),
    .clk_1_E_in(clk_1_wires[121]),
    .prog_clk_1_S_out(prog_clk_1_wires[123]),
    .prog_clk_1_N_out(prog_clk_1_wires[122]),
    .prog_clk_1_E_in(prog_clk_1_wires[121]),
    .prog_clk_0_N_in(prog_clk_0_wires[210]),
    .pReset_S_out(pResetWires[570]),
    .pReset_E_in(pResetWires[569]),
    .pReset_W_out(pResetWires[568]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[54]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[54]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[54]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[54]),
    .SC_OUT_BOT(scff_Wires[109]),
    .SC_IN_TOP(scff_Wires[108]),
    .chanx_left_in(sb_1__1__43_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__54_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__54_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__54_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__54_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__54_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__54_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__54_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__54_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__54_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__54_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__54_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__54_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__54_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__54_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__54_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__54_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__54_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__54_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__54_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__54_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__54_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__1_
  (
    .clk_1_S_out(clk_1_wires[90]),
    .clk_1_N_out(clk_1_wires[89]),
    .clk_1_W_in(clk_1_wires[85]),
    .prog_clk_1_S_out(prog_clk_1_wires[90]),
    .prog_clk_1_N_out(prog_clk_1_wires[89]),
    .prog_clk_1_W_in(prog_clk_1_wires[85]),
    .prog_clk_0_N_in(prog_clk_0_wires[218]),
    .pReset_S_out(pResetWires[84]),
    .pReset_E_in(pResetWires[83]),
    .pReset_W_out(pResetWires[82]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[55]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[55]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[55]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[55]),
    .SC_OUT_TOP(scff_Wires[136]),
    .SC_IN_BOT(scff_Wires[135]),
    .chanx_left_in(sb_1__1__44_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__55_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__55_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__55_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__55_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__55_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__55_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__55_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__55_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__55_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__55_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__55_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__55_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__55_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__55_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__55_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__55_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__55_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__55_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__55_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__55_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__55_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[221]),
    .pReset_S_out(pResetWires[133]),
    .pReset_E_in(pResetWires[132]),
    .pReset_W_out(pResetWires[131]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[56]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[56]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[56]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[56]),
    .SC_OUT_TOP(scff_Wires[138]),
    .SC_IN_BOT(scff_Wires[137]),
    .chanx_left_in(sb_1__1__45_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__56_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__56_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__56_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__56_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__56_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__56_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__56_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__56_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__56_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__56_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__56_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__56_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__56_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__56_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__56_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__56_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__56_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__56_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__56_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__56_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__56_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__3_
  (
    .clk_1_S_out(clk_1_wires[97]),
    .clk_1_N_out(clk_1_wires[96]),
    .clk_1_W_in(clk_1_wires[92]),
    .prog_clk_1_S_out(prog_clk_1_wires[97]),
    .prog_clk_1_N_out(prog_clk_1_wires[96]),
    .prog_clk_1_W_in(prog_clk_1_wires[92]),
    .prog_clk_0_N_in(prog_clk_0_wires[224]),
    .pReset_S_out(pResetWires[182]),
    .pReset_E_in(pResetWires[181]),
    .pReset_W_out(pResetWires[180]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[57]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[57]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[57]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[57]),
    .SC_OUT_TOP(scff_Wires[140]),
    .SC_IN_BOT(scff_Wires[139]),
    .chanx_left_in(sb_1__1__46_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__57_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__57_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__57_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__57_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__57_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__57_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__57_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__57_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__57_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__57_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__57_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__57_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__57_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__57_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__57_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__57_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__57_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__57_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__57_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__57_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__57_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[227]),
    .pReset_S_out(pResetWires[231]),
    .pReset_E_in(pResetWires[230]),
    .pReset_W_out(pResetWires[229]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[58]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[58]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[58]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[58]),
    .SC_OUT_TOP(scff_Wires[142]),
    .SC_IN_BOT(scff_Wires[141]),
    .chanx_left_in(sb_1__1__47_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__58_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__58_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__58_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__58_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__58_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__58_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__58_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__58_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__58_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__58_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__58_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__58_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__58_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__58_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__58_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__58_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__58_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__58_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__58_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__58_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__58_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__5_
  (
    .clk_1_S_out(clk_1_wires[104]),
    .clk_1_N_out(clk_1_wires[103]),
    .clk_1_W_in(clk_1_wires[99]),
    .prog_clk_1_S_out(prog_clk_1_wires[104]),
    .prog_clk_1_N_out(prog_clk_1_wires[103]),
    .prog_clk_1_W_in(prog_clk_1_wires[99]),
    .prog_clk_0_N_in(prog_clk_0_wires[230]),
    .pReset_S_out(pResetWires[280]),
    .pReset_E_in(pResetWires[279]),
    .pReset_W_out(pResetWires[278]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[59]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[59]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[59]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[59]),
    .SC_OUT_TOP(scff_Wires[144]),
    .SC_IN_BOT(scff_Wires[143]),
    .chanx_left_in(sb_1__1__48_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__59_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__59_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__59_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__59_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__59_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__59_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__59_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__59_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__59_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__59_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__59_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__59_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__59_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__59_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__59_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__59_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__59_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__59_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__59_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__59_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__59_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__6_
  (
    .clk_3_W_out(clk_3_wires[3]),
    .clk_3_E_in(clk_3_wires[2]),
    .prog_clk_3_W_out(prog_clk_3_wires[3]),
    .prog_clk_3_E_in(prog_clk_3_wires[2]),
    .prog_clk_0_N_in(prog_clk_0_wires[233]),
    .pReset_S_out(pResetWires[329]),
    .pReset_E_in(pResetWires[328]),
    .pReset_W_out(pResetWires[327]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[60]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[60]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[60]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[60]),
    .SC_OUT_TOP(scff_Wires[146]),
    .SC_IN_BOT(scff_Wires[145]),
    .chanx_left_in(sb_1__1__49_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__60_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__60_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__60_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__60_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__60_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__60_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__60_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__60_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__60_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__60_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__60_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__60_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__60_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__60_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__60_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__60_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__60_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__60_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__60_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__60_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__60_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__7_
  (
    .clk_1_S_out(clk_1_wires[111]),
    .clk_1_N_out(clk_1_wires[110]),
    .clk_1_W_in(clk_1_wires[106]),
    .prog_clk_1_S_out(prog_clk_1_wires[111]),
    .prog_clk_1_N_out(prog_clk_1_wires[110]),
    .prog_clk_1_W_in(prog_clk_1_wires[106]),
    .prog_clk_0_N_in(prog_clk_0_wires[236]),
    .pReset_S_out(pResetWires[378]),
    .pReset_E_in(pResetWires[377]),
    .pReset_W_out(pResetWires[376]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[61]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[61]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[61]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[61]),
    .SC_OUT_TOP(scff_Wires[148]),
    .SC_IN_BOT(scff_Wires[147]),
    .chanx_left_in(sb_1__1__50_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__61_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__61_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__61_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__61_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__61_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__61_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__61_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__61_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__61_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__61_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__61_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__61_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__61_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__61_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__61_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__61_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__61_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__61_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__61_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__61_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__61_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[239]),
    .pReset_S_out(pResetWires[427]),
    .pReset_E_in(pResetWires[426]),
    .pReset_W_out(pResetWires[425]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[62]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[62]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[62]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[62]),
    .SC_OUT_TOP(scff_Wires[150]),
    .SC_IN_BOT(scff_Wires[149]),
    .chanx_left_in(sb_1__1__51_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__62_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__62_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__62_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__62_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__62_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__62_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__62_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__62_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__62_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__62_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__62_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__62_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__62_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__62_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__62_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__62_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__62_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__62_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__62_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__62_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__62_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__9_
  (
    .clk_1_S_out(clk_1_wires[118]),
    .clk_1_N_out(clk_1_wires[117]),
    .clk_1_W_in(clk_1_wires[113]),
    .prog_clk_1_S_out(prog_clk_1_wires[118]),
    .prog_clk_1_N_out(prog_clk_1_wires[117]),
    .prog_clk_1_W_in(prog_clk_1_wires[113]),
    .prog_clk_0_N_in(prog_clk_0_wires[242]),
    .pReset_S_out(pResetWires[476]),
    .pReset_E_in(pResetWires[475]),
    .pReset_W_out(pResetWires[474]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[63]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[63]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[63]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[63]),
    .SC_OUT_TOP(scff_Wires[152]),
    .SC_IN_BOT(scff_Wires[151]),
    .chanx_left_in(sb_1__1__52_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__63_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__63_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__63_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__63_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__63_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__63_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__63_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__63_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__63_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__63_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__63_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__63_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__63_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__63_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__63_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__63_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__63_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__63_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__63_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__63_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__63_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[245]),
    .pReset_S_out(pResetWires[525]),
    .pReset_E_in(pResetWires[524]),
    .pReset_W_out(pResetWires[523]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[64]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[64]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[64]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[64]),
    .SC_OUT_TOP(scff_Wires[154]),
    .SC_IN_BOT(scff_Wires[153]),
    .chanx_left_in(sb_1__1__53_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__64_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__64_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__64_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__64_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__64_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__64_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__64_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__64_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__64_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__64_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__64_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__64_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__64_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__64_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__64_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__64_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__64_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__64_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__64_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__64_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__64_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__11_
  (
    .clk_1_S_out(clk_1_wires[125]),
    .clk_1_N_out(clk_1_wires[124]),
    .clk_1_W_in(clk_1_wires[120]),
    .prog_clk_1_S_out(prog_clk_1_wires[125]),
    .prog_clk_1_N_out(prog_clk_1_wires[124]),
    .prog_clk_1_W_in(prog_clk_1_wires[120]),
    .prog_clk_0_N_in(prog_clk_0_wires[248]),
    .pReset_S_out(pResetWires[574]),
    .pReset_E_in(pResetWires[573]),
    .pReset_W_out(pResetWires[572]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[65]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[65]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[65]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[65]),
    .SC_OUT_TOP(scff_Wires[156]),
    .SC_IN_BOT(scff_Wires[155]),
    .chanx_left_in(sb_1__1__54_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__65_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__65_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__65_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__65_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__65_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__65_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__65_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__65_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__65_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__65_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__65_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__65_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__65_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__65_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__65_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__65_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__65_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__65_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__65_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__65_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__65_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__1_
  (
    .clk_1_S_out(clk_1_wires[130]),
    .clk_1_N_out(clk_1_wires[129]),
    .clk_1_E_in(clk_1_wires[128]),
    .prog_clk_1_S_out(prog_clk_1_wires[130]),
    .prog_clk_1_N_out(prog_clk_1_wires[129]),
    .prog_clk_1_E_in(prog_clk_1_wires[128]),
    .prog_clk_0_N_in(prog_clk_0_wires[256]),
    .pReset_S_out(pResetWires[88]),
    .pReset_E_out(pResetWires[87]),
    .pReset_W_in(pResetWires[86]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[66]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[66]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[66]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[66]),
    .SC_OUT_BOT(scff_Wires[182]),
    .SC_IN_TOP(scff_Wires[181]),
    .chanx_left_in(sb_1__1__55_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__66_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__66_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__66_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__66_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__66_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__66_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__66_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__66_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__66_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__66_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__66_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__66_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__66_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__66_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__66_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__66_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__66_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__66_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__66_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__66_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__66_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[259]),
    .pReset_S_out(pResetWires[137]),
    .pReset_E_out(pResetWires[136]),
    .pReset_W_in(pResetWires[135]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[67]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[67]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[67]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[67]),
    .SC_OUT_BOT(scff_Wires[180]),
    .SC_IN_TOP(scff_Wires[179]),
    .chanx_left_in(sb_1__1__56_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__67_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__67_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__67_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__67_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__67_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__67_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__67_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__67_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__67_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__67_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__67_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__67_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__67_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__67_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__67_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__67_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__67_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__67_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__67_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__67_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__67_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__3_
  (
    .clk_1_S_out(clk_1_wires[137]),
    .clk_1_N_out(clk_1_wires[136]),
    .clk_1_E_in(clk_1_wires[135]),
    .prog_clk_1_S_out(prog_clk_1_wires[137]),
    .prog_clk_1_N_out(prog_clk_1_wires[136]),
    .prog_clk_1_E_in(prog_clk_1_wires[135]),
    .prog_clk_0_N_in(prog_clk_0_wires[262]),
    .pReset_S_out(pResetWires[186]),
    .pReset_E_out(pResetWires[185]),
    .pReset_W_in(pResetWires[184]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[68]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[68]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[68]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[68]),
    .SC_OUT_BOT(scff_Wires[178]),
    .SC_IN_TOP(scff_Wires[177]),
    .chanx_left_in(sb_1__1__57_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__68_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__68_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__68_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__68_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__68_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__68_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__68_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__68_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__68_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__68_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__68_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__68_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__68_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__68_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__68_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__68_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__68_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__68_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__68_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__68_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__68_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[265]),
    .pReset_S_out(pResetWires[235]),
    .pReset_E_out(pResetWires[234]),
    .pReset_W_in(pResetWires[233]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[69]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[69]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[69]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[69]),
    .SC_OUT_BOT(scff_Wires[176]),
    .SC_IN_TOP(scff_Wires[175]),
    .chanx_left_in(sb_1__1__58_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__69_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__69_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__69_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__69_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__69_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__69_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__69_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__69_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__69_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__69_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__69_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__69_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__69_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__69_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__69_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__69_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__69_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__69_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__69_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__69_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__69_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__5_
  (
    .clk_1_S_out(clk_1_wires[144]),
    .clk_1_N_out(clk_1_wires[143]),
    .clk_1_E_in(clk_1_wires[142]),
    .prog_clk_1_S_out(prog_clk_1_wires[144]),
    .prog_clk_1_N_out(prog_clk_1_wires[143]),
    .prog_clk_1_E_in(prog_clk_1_wires[142]),
    .prog_clk_0_N_in(prog_clk_0_wires[268]),
    .pReset_S_out(pResetWires[284]),
    .pReset_E_out(pResetWires[283]),
    .pReset_W_in(pResetWires[282]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[70]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[70]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[70]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[70]),
    .SC_OUT_BOT(scff_Wires[174]),
    .SC_IN_TOP(scff_Wires[173]),
    .chanx_left_in(sb_1__1__59_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__70_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__70_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__70_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__70_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__70_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__70_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__70_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__70_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__70_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__70_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__70_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__70_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__70_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__70_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__70_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__70_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__70_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__70_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__70_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__70_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__70_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__6_
  (
    .clk_3_E_out(clk_3_wires[1]),
    .clk_3_W_in(clk_3_wires[0]),
    .prog_clk_3_E_out(prog_clk_3_wires[1]),
    .prog_clk_3_W_in(prog_clk_3_wires[0]),
    .prog_clk_0_N_in(prog_clk_0_wires[271]),
    .pReset_S_out(pResetWires[333]),
    .pReset_E_out(pResetWires[332]),
    .pReset_W_in(pResetWires[331]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[71]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[71]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[71]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[71]),
    .SC_OUT_BOT(scff_Wires[172]),
    .SC_IN_TOP(scff_Wires[171]),
    .chanx_left_in(sb_1__1__60_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__71_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__71_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__71_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__71_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__71_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__71_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__71_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__71_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__71_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__71_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__71_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__71_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__71_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__71_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__71_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__71_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__71_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__71_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__71_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__71_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__71_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__7_
  (
    .clk_1_S_out(clk_1_wires[151]),
    .clk_1_N_out(clk_1_wires[150]),
    .clk_1_E_in(clk_1_wires[149]),
    .prog_clk_1_S_out(prog_clk_1_wires[151]),
    .prog_clk_1_N_out(prog_clk_1_wires[150]),
    .prog_clk_1_E_in(prog_clk_1_wires[149]),
    .prog_clk_0_N_in(prog_clk_0_wires[274]),
    .pReset_S_out(pResetWires[382]),
    .pReset_E_out(pResetWires[381]),
    .pReset_W_in(pResetWires[380]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[72]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[72]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[72]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[72]),
    .SC_OUT_BOT(scff_Wires[170]),
    .SC_IN_TOP(scff_Wires[169]),
    .chanx_left_in(sb_1__1__61_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__72_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__72_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__72_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__72_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__72_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__72_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__72_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__72_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__72_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__72_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__72_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__72_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__72_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__72_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__72_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__72_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__72_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__72_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__72_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__72_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__72_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[277]),
    .pReset_S_out(pResetWires[431]),
    .pReset_E_out(pResetWires[430]),
    .pReset_W_in(pResetWires[429]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[73]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[73]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[73]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[73]),
    .SC_OUT_BOT(scff_Wires[168]),
    .SC_IN_TOP(scff_Wires[167]),
    .chanx_left_in(sb_1__1__62_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__73_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__73_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__73_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__73_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__73_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__73_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__73_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__73_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__73_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__73_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__73_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__73_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__73_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__73_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__73_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__73_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__73_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__73_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__73_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__73_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__73_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__9_
  (
    .clk_1_S_out(clk_1_wires[158]),
    .clk_1_N_out(clk_1_wires[157]),
    .clk_1_E_in(clk_1_wires[156]),
    .prog_clk_1_S_out(prog_clk_1_wires[158]),
    .prog_clk_1_N_out(prog_clk_1_wires[157]),
    .prog_clk_1_E_in(prog_clk_1_wires[156]),
    .prog_clk_0_N_in(prog_clk_0_wires[280]),
    .pReset_S_out(pResetWires[480]),
    .pReset_E_out(pResetWires[479]),
    .pReset_W_in(pResetWires[478]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[74]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[74]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[74]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[74]),
    .SC_OUT_BOT(scff_Wires[166]),
    .SC_IN_TOP(scff_Wires[165]),
    .chanx_left_in(sb_1__1__63_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__74_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__74_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__74_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__74_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__74_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__74_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__74_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__74_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__74_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__74_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__74_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__74_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__74_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__74_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__74_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__74_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__74_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__74_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__74_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__74_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__74_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[283]),
    .pReset_S_out(pResetWires[529]),
    .pReset_E_out(pResetWires[528]),
    .pReset_W_in(pResetWires[527]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[75]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[75]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[75]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[75]),
    .SC_OUT_BOT(scff_Wires[164]),
    .SC_IN_TOP(scff_Wires[163]),
    .chanx_left_in(sb_1__1__64_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__75_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__75_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__75_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__75_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__75_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__75_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__75_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__75_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__75_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__75_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__75_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__75_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__75_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__75_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__75_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__75_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__75_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__75_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__75_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__75_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__75_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__11_
  (
    .clk_1_S_out(clk_1_wires[165]),
    .clk_1_N_out(clk_1_wires[164]),
    .clk_1_E_in(clk_1_wires[163]),
    .prog_clk_1_S_out(prog_clk_1_wires[165]),
    .prog_clk_1_N_out(prog_clk_1_wires[164]),
    .prog_clk_1_E_in(prog_clk_1_wires[163]),
    .prog_clk_0_N_in(prog_clk_0_wires[286]),
    .pReset_S_out(pResetWires[578]),
    .pReset_E_out(pResetWires[577]),
    .pReset_W_in(pResetWires[576]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[76]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[76]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[76]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[76]),
    .SC_OUT_BOT(scff_Wires[162]),
    .SC_IN_TOP(scff_Wires[161]),
    .chanx_left_in(sb_1__1__65_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__76_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__76_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__76_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__76_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__76_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__76_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__76_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__76_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__76_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__76_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__76_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__76_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__76_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__76_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__76_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__76_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__76_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__76_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__76_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__76_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__76_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__1_
  (
    .clk_1_S_out(clk_1_wires[132]),
    .clk_1_N_out(clk_1_wires[131]),
    .clk_1_W_in(clk_1_wires[127]),
    .prog_clk_1_S_out(prog_clk_1_wires[132]),
    .prog_clk_1_N_out(prog_clk_1_wires[131]),
    .prog_clk_1_W_in(prog_clk_1_wires[127]),
    .prog_clk_0_N_in(prog_clk_0_wires[294]),
    .pReset_S_out(pResetWires[92]),
    .pReset_E_out(pResetWires[91]),
    .pReset_W_in(pResetWires[90]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[77]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[77]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[77]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[77]),
    .SC_OUT_TOP(scff_Wires[189]),
    .SC_IN_BOT(scff_Wires[188]),
    .chanx_left_in(sb_1__1__66_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__77_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__77_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__77_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__77_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__77_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__77_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__77_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__77_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__77_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__77_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__77_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__77_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__77_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__77_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__77_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__77_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__77_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__77_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__77_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__77_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__77_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__2_
  (
    .clk_2_W_out(clk_2_wires[72]),
    .clk_2_E_in(clk_2_wires[71]),
    .prog_clk_2_W_out(prog_clk_2_wires[72]),
    .prog_clk_2_E_in(prog_clk_2_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[297]),
    .pReset_S_out(pResetWires[141]),
    .pReset_E_out(pResetWires[140]),
    .pReset_W_in(pResetWires[139]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[78]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[78]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[78]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[78]),
    .SC_OUT_TOP(scff_Wires[191]),
    .SC_IN_BOT(scff_Wires[190]),
    .chanx_left_in(sb_1__1__67_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__78_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__78_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__78_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__78_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__78_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__78_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__78_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__78_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__78_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__78_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__78_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__78_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__78_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__78_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__78_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__78_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__78_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__78_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__78_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__78_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__78_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__3_
  (
    .clk_1_S_out(clk_1_wires[139]),
    .clk_1_N_out(clk_1_wires[138]),
    .clk_1_W_in(clk_1_wires[134]),
    .prog_clk_1_S_out(prog_clk_1_wires[139]),
    .prog_clk_1_N_out(prog_clk_1_wires[138]),
    .prog_clk_1_W_in(prog_clk_1_wires[134]),
    .prog_clk_0_N_in(prog_clk_0_wires[300]),
    .pReset_S_out(pResetWires[190]),
    .pReset_E_out(pResetWires[189]),
    .pReset_W_in(pResetWires[188]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[79]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[79]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[79]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[79]),
    .SC_OUT_TOP(scff_Wires[193]),
    .SC_IN_BOT(scff_Wires[192]),
    .chanx_left_in(sb_1__1__68_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__79_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__79_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__79_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__79_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__79_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__79_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__79_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__79_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__79_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__79_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__79_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__79_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__79_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__79_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__79_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__79_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__79_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__79_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__79_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__79_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__79_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__4_
  (
    .clk_2_W_out(clk_2_wires[81]),
    .clk_2_E_in(clk_2_wires[80]),
    .prog_clk_2_W_out(prog_clk_2_wires[81]),
    .prog_clk_2_E_in(prog_clk_2_wires[80]),
    .prog_clk_0_N_in(prog_clk_0_wires[303]),
    .pReset_S_out(pResetWires[239]),
    .pReset_E_out(pResetWires[238]),
    .pReset_W_in(pResetWires[237]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[80]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[80]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[80]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[80]),
    .SC_OUT_TOP(scff_Wires[195]),
    .SC_IN_BOT(scff_Wires[194]),
    .chanx_left_in(sb_1__1__69_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__80_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__80_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__80_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__80_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__80_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__80_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__80_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__80_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__80_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__80_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__80_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__80_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__80_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__80_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__80_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__80_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__80_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__80_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__80_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__80_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__80_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__5_
  (
    .clk_1_S_out(clk_1_wires[146]),
    .clk_1_N_out(clk_1_wires[145]),
    .clk_1_W_in(clk_1_wires[141]),
    .prog_clk_1_S_out(prog_clk_1_wires[146]),
    .prog_clk_1_N_out(prog_clk_1_wires[145]),
    .prog_clk_1_W_in(prog_clk_1_wires[141]),
    .prog_clk_0_N_in(prog_clk_0_wires[306]),
    .pReset_S_out(pResetWires[288]),
    .pReset_E_out(pResetWires[287]),
    .pReset_W_in(pResetWires[286]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[81]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[81]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[81]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[81]),
    .SC_OUT_TOP(scff_Wires[197]),
    .SC_IN_BOT(scff_Wires[196]),
    .chanx_left_in(sb_1__1__70_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__81_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__81_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__81_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__81_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__81_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__81_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__81_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__81_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__81_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__81_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__81_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__81_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__81_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__81_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__81_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__81_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__81_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__81_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__81_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__81_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__81_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__6_
  (
    .clk_3_E_out(clk_3_wires[5]),
    .clk_3_W_in(clk_3_wires[4]),
    .prog_clk_3_E_out(prog_clk_3_wires[5]),
    .prog_clk_3_W_in(prog_clk_3_wires[4]),
    .prog_clk_0_N_in(prog_clk_0_wires[309]),
    .pReset_S_out(pResetWires[337]),
    .pReset_E_out(pResetWires[336]),
    .pReset_W_in(pResetWires[335]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[82]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[82]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[82]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[82]),
    .SC_OUT_TOP(scff_Wires[199]),
    .SC_IN_BOT(scff_Wires[198]),
    .chanx_left_in(sb_1__1__71_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__82_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__82_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__82_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__82_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__82_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__82_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__82_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__82_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__82_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__82_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__82_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__82_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__82_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__82_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__82_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__82_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__82_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__82_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__82_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__82_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__82_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__7_
  (
    .clk_1_S_out(clk_1_wires[153]),
    .clk_1_N_out(clk_1_wires[152]),
    .clk_1_W_in(clk_1_wires[148]),
    .prog_clk_1_S_out(prog_clk_1_wires[153]),
    .prog_clk_1_N_out(prog_clk_1_wires[152]),
    .prog_clk_1_W_in(prog_clk_1_wires[148]),
    .prog_clk_0_N_in(prog_clk_0_wires[312]),
    .pReset_S_out(pResetWires[386]),
    .pReset_E_out(pResetWires[385]),
    .pReset_W_in(pResetWires[384]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[83]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[83]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[83]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[83]),
    .SC_OUT_TOP(scff_Wires[201]),
    .SC_IN_BOT(scff_Wires[200]),
    .chanx_left_in(sb_1__1__72_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__83_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__83_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__83_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__83_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__83_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__83_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__83_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__83_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__83_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__83_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__83_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__83_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__83_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__83_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__83_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__83_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__83_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__83_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__83_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__83_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__83_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__8_
  (
    .clk_2_W_out(clk_2_wires[94]),
    .clk_2_E_in(clk_2_wires[93]),
    .prog_clk_2_W_out(prog_clk_2_wires[94]),
    .prog_clk_2_E_in(prog_clk_2_wires[93]),
    .prog_clk_0_N_in(prog_clk_0_wires[315]),
    .pReset_S_out(pResetWires[435]),
    .pReset_E_out(pResetWires[434]),
    .pReset_W_in(pResetWires[433]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[84]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[84]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[84]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[84]),
    .SC_OUT_TOP(scff_Wires[203]),
    .SC_IN_BOT(scff_Wires[202]),
    .chanx_left_in(sb_1__1__73_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__84_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__84_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__84_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__84_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__84_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__84_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__84_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__84_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__84_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__84_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__84_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__84_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__84_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__84_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__84_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__84_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__84_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__84_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__84_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__84_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__84_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__9_
  (
    .clk_1_S_out(clk_1_wires[160]),
    .clk_1_N_out(clk_1_wires[159]),
    .clk_1_W_in(clk_1_wires[155]),
    .prog_clk_1_S_out(prog_clk_1_wires[160]),
    .prog_clk_1_N_out(prog_clk_1_wires[159]),
    .prog_clk_1_W_in(prog_clk_1_wires[155]),
    .prog_clk_0_N_in(prog_clk_0_wires[318]),
    .pReset_S_out(pResetWires[484]),
    .pReset_E_out(pResetWires[483]),
    .pReset_W_in(pResetWires[482]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[85]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[85]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[85]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[85]),
    .SC_OUT_TOP(scff_Wires[205]),
    .SC_IN_BOT(scff_Wires[204]),
    .chanx_left_in(sb_1__1__74_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__85_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__85_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__85_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__85_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__85_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__85_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__85_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__85_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__85_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__85_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__85_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__85_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__85_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__85_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__85_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__85_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__85_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__85_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__85_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__85_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__85_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__10_
  (
    .clk_2_W_out(clk_2_wires[107]),
    .clk_2_E_in(clk_2_wires[106]),
    .prog_clk_2_W_out(prog_clk_2_wires[107]),
    .prog_clk_2_E_in(prog_clk_2_wires[106]),
    .prog_clk_0_N_in(prog_clk_0_wires[321]),
    .pReset_S_out(pResetWires[533]),
    .pReset_E_out(pResetWires[532]),
    .pReset_W_in(pResetWires[531]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[86]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[86]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[86]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[86]),
    .SC_OUT_TOP(scff_Wires[207]),
    .SC_IN_BOT(scff_Wires[206]),
    .chanx_left_in(sb_1__1__75_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__86_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__86_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__86_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__86_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__86_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__86_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__86_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__86_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__86_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__86_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__86_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__86_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__86_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__86_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__86_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__86_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__86_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__86_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__86_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__86_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__86_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__11_
  (
    .clk_1_S_out(clk_1_wires[167]),
    .clk_1_N_out(clk_1_wires[166]),
    .clk_1_W_in(clk_1_wires[162]),
    .prog_clk_1_S_out(prog_clk_1_wires[167]),
    .prog_clk_1_N_out(prog_clk_1_wires[166]),
    .prog_clk_1_W_in(prog_clk_1_wires[162]),
    .prog_clk_0_N_in(prog_clk_0_wires[324]),
    .pReset_S_out(pResetWires[582]),
    .pReset_E_out(pResetWires[581]),
    .pReset_W_in(pResetWires[580]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[87]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[87]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[87]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[87]),
    .SC_OUT_TOP(scff_Wires[209]),
    .SC_IN_BOT(scff_Wires[208]),
    .chanx_left_in(sb_1__1__76_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__87_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__87_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__87_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__87_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__87_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__87_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__87_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__87_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__87_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__87_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__87_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__87_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__87_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__87_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__87_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__87_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__87_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__87_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__87_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__87_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__87_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__1_
  (
    .clk_1_S_out(clk_1_wires[172]),
    .clk_1_N_out(clk_1_wires[171]),
    .clk_1_E_in(clk_1_wires[170]),
    .prog_clk_1_S_out(prog_clk_1_wires[172]),
    .prog_clk_1_N_out(prog_clk_1_wires[171]),
    .prog_clk_1_E_in(prog_clk_1_wires[170]),
    .prog_clk_0_N_in(prog_clk_0_wires[332]),
    .pReset_S_out(pResetWires[96]),
    .pReset_E_out(pResetWires[95]),
    .pReset_W_in(pResetWires[94]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[88]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[88]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[88]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[88]),
    .SC_OUT_BOT(scff_Wires[235]),
    .SC_IN_TOP(scff_Wires[234]),
    .chanx_left_in(sb_1__1__77_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__88_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__88_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__88_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__88_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__88_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__88_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__88_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__88_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__88_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__88_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__88_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__88_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__88_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__88_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__88_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__88_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__88_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__88_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__88_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__88_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__88_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__2_
  (
    .clk_2_E_out(clk_2_wires[70]),
    .clk_2_W_in(clk_2_wires[69]),
    .prog_clk_2_E_out(prog_clk_2_wires[70]),
    .prog_clk_2_W_in(prog_clk_2_wires[69]),
    .prog_clk_0_N_in(prog_clk_0_wires[335]),
    .pReset_S_out(pResetWires[145]),
    .pReset_E_out(pResetWires[144]),
    .pReset_W_in(pResetWires[143]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[89]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[89]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[89]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[89]),
    .SC_OUT_BOT(scff_Wires[233]),
    .SC_IN_TOP(scff_Wires[232]),
    .chanx_left_in(sb_1__1__78_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__89_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__89_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__89_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__89_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__89_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__89_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__89_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__89_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__89_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__89_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__89_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__89_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__89_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__89_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__89_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__89_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__89_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__89_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__89_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__89_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__89_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__3_
  (
    .clk_1_S_out(clk_1_wires[179]),
    .clk_1_N_out(clk_1_wires[178]),
    .clk_1_E_in(clk_1_wires[177]),
    .prog_clk_1_S_out(prog_clk_1_wires[179]),
    .prog_clk_1_N_out(prog_clk_1_wires[178]),
    .prog_clk_1_E_in(prog_clk_1_wires[177]),
    .prog_clk_0_N_in(prog_clk_0_wires[338]),
    .pReset_S_out(pResetWires[194]),
    .pReset_E_out(pResetWires[193]),
    .pReset_W_in(pResetWires[192]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[90]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[90]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[90]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[90]),
    .SC_OUT_BOT(scff_Wires[231]),
    .SC_IN_TOP(scff_Wires[230]),
    .chanx_left_in(sb_1__1__79_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__90_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__90_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__90_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__90_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__90_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__90_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__90_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__90_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__90_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__90_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__90_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__90_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__90_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__90_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__90_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__90_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__90_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__90_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__90_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__90_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__90_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__4_
  (
    .clk_2_E_out(clk_2_wires[79]),
    .clk_2_W_in(clk_2_wires[78]),
    .prog_clk_2_E_out(prog_clk_2_wires[79]),
    .prog_clk_2_W_in(prog_clk_2_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[341]),
    .pReset_S_out(pResetWires[243]),
    .pReset_E_out(pResetWires[242]),
    .pReset_W_in(pResetWires[241]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[91]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[91]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[91]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[91]),
    .SC_OUT_BOT(scff_Wires[229]),
    .SC_IN_TOP(scff_Wires[228]),
    .chanx_left_in(sb_1__1__80_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__91_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__91_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__91_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__91_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__91_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__91_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__91_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__91_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__91_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__91_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__91_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__91_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__91_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__91_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__91_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__91_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__91_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__91_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__91_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__91_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__91_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__5_
  (
    .clk_1_S_out(clk_1_wires[186]),
    .clk_1_N_out(clk_1_wires[185]),
    .clk_1_E_in(clk_1_wires[184]),
    .prog_clk_1_S_out(prog_clk_1_wires[186]),
    .prog_clk_1_N_out(prog_clk_1_wires[185]),
    .prog_clk_1_E_in(prog_clk_1_wires[184]),
    .prog_clk_0_N_in(prog_clk_0_wires[344]),
    .pReset_S_out(pResetWires[292]),
    .pReset_E_out(pResetWires[291]),
    .pReset_W_in(pResetWires[290]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[92]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[92]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[92]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[92]),
    .SC_OUT_BOT(scff_Wires[227]),
    .SC_IN_TOP(scff_Wires[226]),
    .chanx_left_in(sb_1__1__81_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__92_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__92_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__92_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__92_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__92_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__92_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__92_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__92_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__92_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__92_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__92_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__92_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__92_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__92_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__92_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__92_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__92_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__92_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__92_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__92_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__92_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__6_
  (
    .clk_3_E_out(clk_3_wires[45]),
    .clk_3_W_in(clk_3_wires[44]),
    .prog_clk_3_E_out(prog_clk_3_wires[45]),
    .prog_clk_3_W_in(prog_clk_3_wires[44]),
    .prog_clk_0_N_in(prog_clk_0_wires[347]),
    .pReset_S_out(pResetWires[341]),
    .pReset_E_out(pResetWires[340]),
    .pReset_W_in(pResetWires[339]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[93]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[93]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[93]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[93]),
    .SC_OUT_BOT(scff_Wires[225]),
    .SC_IN_TOP(scff_Wires[224]),
    .chanx_left_in(sb_1__1__82_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__93_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__93_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__93_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__93_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__93_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__93_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__93_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__93_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__93_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__93_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__93_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__93_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__93_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__93_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__93_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__93_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__93_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__93_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__93_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__93_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__93_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__7_
  (
    .clk_1_S_out(clk_1_wires[193]),
    .clk_1_N_out(clk_1_wires[192]),
    .clk_1_E_in(clk_1_wires[191]),
    .prog_clk_1_S_out(prog_clk_1_wires[193]),
    .prog_clk_1_N_out(prog_clk_1_wires[192]),
    .prog_clk_1_E_in(prog_clk_1_wires[191]),
    .prog_clk_0_N_in(prog_clk_0_wires[350]),
    .pReset_S_out(pResetWires[390]),
    .pReset_E_out(pResetWires[389]),
    .pReset_W_in(pResetWires[388]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[94]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[94]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[94]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[94]),
    .SC_OUT_BOT(scff_Wires[223]),
    .SC_IN_TOP(scff_Wires[222]),
    .chanx_left_in(sb_1__1__83_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__94_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__94_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__94_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__94_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__94_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__94_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__94_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__94_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__94_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__94_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__94_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__94_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__94_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__94_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__94_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__94_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__94_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__94_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__94_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__94_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__94_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__8_
  (
    .clk_2_E_out(clk_2_wires[92]),
    .clk_2_W_in(clk_2_wires[91]),
    .prog_clk_2_E_out(prog_clk_2_wires[92]),
    .prog_clk_2_W_in(prog_clk_2_wires[91]),
    .prog_clk_0_N_in(prog_clk_0_wires[353]),
    .pReset_S_out(pResetWires[439]),
    .pReset_E_out(pResetWires[438]),
    .pReset_W_in(pResetWires[437]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[95]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[95]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[95]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[95]),
    .SC_OUT_BOT(scff_Wires[221]),
    .SC_IN_TOP(scff_Wires[220]),
    .chanx_left_in(sb_1__1__84_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__95_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__95_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__95_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__95_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__95_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__95_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__95_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__95_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__95_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__95_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__95_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__95_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__95_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__95_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__95_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__95_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__95_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__95_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__95_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__95_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__95_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__9_
  (
    .clk_1_S_out(clk_1_wires[200]),
    .clk_1_N_out(clk_1_wires[199]),
    .clk_1_E_in(clk_1_wires[198]),
    .prog_clk_1_S_out(prog_clk_1_wires[200]),
    .prog_clk_1_N_out(prog_clk_1_wires[199]),
    .prog_clk_1_E_in(prog_clk_1_wires[198]),
    .prog_clk_0_N_in(prog_clk_0_wires[356]),
    .pReset_S_out(pResetWires[488]),
    .pReset_E_out(pResetWires[487]),
    .pReset_W_in(pResetWires[486]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[96]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[96]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[96]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[96]),
    .SC_OUT_BOT(scff_Wires[219]),
    .SC_IN_TOP(scff_Wires[218]),
    .chanx_left_in(sb_1__1__85_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__96_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__96_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__96_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__96_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__96_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__96_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__96_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__96_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__96_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__96_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__96_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__96_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__96_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__96_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__96_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__96_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__96_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__96_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__96_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__96_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__96_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__10_
  (
    .clk_2_E_out(clk_2_wires[105]),
    .clk_2_W_in(clk_2_wires[104]),
    .prog_clk_2_E_out(prog_clk_2_wires[105]),
    .prog_clk_2_W_in(prog_clk_2_wires[104]),
    .prog_clk_0_N_in(prog_clk_0_wires[359]),
    .pReset_S_out(pResetWires[537]),
    .pReset_E_out(pResetWires[536]),
    .pReset_W_in(pResetWires[535]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[97]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[97]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[97]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[97]),
    .SC_OUT_BOT(scff_Wires[217]),
    .SC_IN_TOP(scff_Wires[216]),
    .chanx_left_in(sb_1__1__86_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__97_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__97_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__97_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__97_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__97_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__97_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__97_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__97_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__97_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__97_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__97_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__97_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__97_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__97_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__97_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__97_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__97_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__97_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__97_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__97_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__97_ccff_tail[0])
  );


  cbx_1__1_
  cbx_9__11_
  (
    .clk_1_S_out(clk_1_wires[207]),
    .clk_1_N_out(clk_1_wires[206]),
    .clk_1_E_in(clk_1_wires[205]),
    .prog_clk_1_S_out(prog_clk_1_wires[207]),
    .prog_clk_1_N_out(prog_clk_1_wires[206]),
    .prog_clk_1_E_in(prog_clk_1_wires[205]),
    .prog_clk_0_N_in(prog_clk_0_wires[362]),
    .pReset_S_out(pResetWires[586]),
    .pReset_E_out(pResetWires[585]),
    .pReset_W_in(pResetWires[584]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[98]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[98]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[98]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[98]),
    .SC_OUT_BOT(scff_Wires[215]),
    .SC_IN_TOP(scff_Wires[214]),
    .chanx_left_in(sb_1__1__87_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__98_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__98_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__98_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__98_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__98_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__98_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__98_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__98_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__98_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__98_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__98_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__98_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__98_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__98_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__98_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__98_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__98_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__98_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__98_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__98_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__98_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__1_
  (
    .clk_1_S_out(clk_1_wires[174]),
    .clk_1_N_out(clk_1_wires[173]),
    .clk_1_W_in(clk_1_wires[169]),
    .prog_clk_1_S_out(prog_clk_1_wires[174]),
    .prog_clk_1_N_out(prog_clk_1_wires[173]),
    .prog_clk_1_W_in(prog_clk_1_wires[169]),
    .prog_clk_0_N_in(prog_clk_0_wires[370]),
    .pReset_S_out(pResetWires[100]),
    .pReset_E_out(pResetWires[99]),
    .pReset_W_in(pResetWires[98]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[99]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[99]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[99]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[99]),
    .SC_OUT_TOP(scff_Wires[242]),
    .SC_IN_BOT(scff_Wires[241]),
    .chanx_left_in(sb_1__1__88_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__99_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__99_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__99_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__99_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__99_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__99_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__99_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__99_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__99_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__99_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__99_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__99_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__99_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__99_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__99_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__99_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__99_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__99_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__99_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__99_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__99_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[373]),
    .pReset_S_out(pResetWires[149]),
    .pReset_E_out(pResetWires[148]),
    .pReset_W_in(pResetWires[147]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[100]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[100]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[100]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[100]),
    .SC_OUT_TOP(scff_Wires[244]),
    .SC_IN_BOT(scff_Wires[243]),
    .chanx_left_in(sb_1__1__89_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__100_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__100_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__100_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__100_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__100_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__100_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__100_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__100_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__100_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__100_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__100_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__100_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__100_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__100_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__100_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__100_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__100_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__100_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__100_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__100_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__100_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__3_
  (
    .clk_1_S_out(clk_1_wires[181]),
    .clk_1_N_out(clk_1_wires[180]),
    .clk_1_W_in(clk_1_wires[176]),
    .prog_clk_1_S_out(prog_clk_1_wires[181]),
    .prog_clk_1_N_out(prog_clk_1_wires[180]),
    .prog_clk_1_W_in(prog_clk_1_wires[176]),
    .prog_clk_0_N_in(prog_clk_0_wires[376]),
    .pReset_S_out(pResetWires[198]),
    .pReset_E_out(pResetWires[197]),
    .pReset_W_in(pResetWires[196]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[101]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[101]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[101]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[101]),
    .SC_OUT_TOP(scff_Wires[246]),
    .SC_IN_BOT(scff_Wires[245]),
    .chanx_left_in(sb_1__1__90_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__101_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__101_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__101_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__101_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__101_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__101_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__101_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__101_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__101_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__101_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__101_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__101_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__101_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__101_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__101_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__101_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__101_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__101_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__101_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__101_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__101_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[379]),
    .pReset_S_out(pResetWires[247]),
    .pReset_E_out(pResetWires[246]),
    .pReset_W_in(pResetWires[245]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[102]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[102]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[102]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[102]),
    .SC_OUT_TOP(scff_Wires[248]),
    .SC_IN_BOT(scff_Wires[247]),
    .chanx_left_in(sb_1__1__91_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__102_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__102_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__102_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__102_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__102_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__102_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__102_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__102_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__102_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__102_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__102_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__102_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__102_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__102_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__102_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__102_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__102_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__102_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__102_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__102_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__102_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__5_
  (
    .clk_1_S_out(clk_1_wires[188]),
    .clk_1_N_out(clk_1_wires[187]),
    .clk_1_W_in(clk_1_wires[183]),
    .prog_clk_1_S_out(prog_clk_1_wires[188]),
    .prog_clk_1_N_out(prog_clk_1_wires[187]),
    .prog_clk_1_W_in(prog_clk_1_wires[183]),
    .prog_clk_0_N_in(prog_clk_0_wires[382]),
    .pReset_S_out(pResetWires[296]),
    .pReset_E_out(pResetWires[295]),
    .pReset_W_in(pResetWires[294]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[103]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[103]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[103]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[103]),
    .SC_OUT_TOP(scff_Wires[250]),
    .SC_IN_BOT(scff_Wires[249]),
    .chanx_left_in(sb_1__1__92_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__103_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__103_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__103_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__103_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__103_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__103_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__103_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__103_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__103_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__103_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__103_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__103_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__103_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__103_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__103_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__103_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__103_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__103_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__103_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__103_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__103_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__6_
  (
    .clk_3_E_out(clk_3_wires[49]),
    .clk_3_W_in(clk_3_wires[48]),
    .prog_clk_3_E_out(prog_clk_3_wires[49]),
    .prog_clk_3_W_in(prog_clk_3_wires[48]),
    .prog_clk_0_N_in(prog_clk_0_wires[385]),
    .pReset_S_out(pResetWires[345]),
    .pReset_E_out(pResetWires[344]),
    .pReset_W_in(pResetWires[343]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[104]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[104]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[104]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[104]),
    .SC_OUT_TOP(scff_Wires[252]),
    .SC_IN_BOT(scff_Wires[251]),
    .chanx_left_in(sb_1__1__93_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__104_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__104_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__104_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__104_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__104_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__104_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__104_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__104_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__104_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__104_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__104_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__104_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__104_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__104_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__104_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__104_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__104_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__104_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__104_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__104_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__104_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__7_
  (
    .clk_1_S_out(clk_1_wires[195]),
    .clk_1_N_out(clk_1_wires[194]),
    .clk_1_W_in(clk_1_wires[190]),
    .prog_clk_1_S_out(prog_clk_1_wires[195]),
    .prog_clk_1_N_out(prog_clk_1_wires[194]),
    .prog_clk_1_W_in(prog_clk_1_wires[190]),
    .prog_clk_0_N_in(prog_clk_0_wires[388]),
    .pReset_S_out(pResetWires[394]),
    .pReset_E_out(pResetWires[393]),
    .pReset_W_in(pResetWires[392]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[105]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[105]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[105]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[105]),
    .SC_OUT_TOP(scff_Wires[254]),
    .SC_IN_BOT(scff_Wires[253]),
    .chanx_left_in(sb_1__1__94_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__105_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__105_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__105_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__105_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__105_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__105_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__105_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__105_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__105_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__105_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__105_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__105_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__105_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__105_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__105_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__105_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__105_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__105_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__105_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__105_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__105_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[391]),
    .pReset_S_out(pResetWires[443]),
    .pReset_E_out(pResetWires[442]),
    .pReset_W_in(pResetWires[441]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[106]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[106]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[106]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[106]),
    .SC_OUT_TOP(scff_Wires[256]),
    .SC_IN_BOT(scff_Wires[255]),
    .chanx_left_in(sb_1__1__95_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__106_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__106_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__106_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__106_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__106_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__106_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__106_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__106_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__106_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__106_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__106_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__106_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__106_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__106_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__106_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__106_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__106_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__106_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__106_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__106_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__106_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__9_
  (
    .clk_1_S_out(clk_1_wires[202]),
    .clk_1_N_out(clk_1_wires[201]),
    .clk_1_W_in(clk_1_wires[197]),
    .prog_clk_1_S_out(prog_clk_1_wires[202]),
    .prog_clk_1_N_out(prog_clk_1_wires[201]),
    .prog_clk_1_W_in(prog_clk_1_wires[197]),
    .prog_clk_0_N_in(prog_clk_0_wires[394]),
    .pReset_S_out(pResetWires[492]),
    .pReset_E_out(pResetWires[491]),
    .pReset_W_in(pResetWires[490]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[107]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[107]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[107]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[107]),
    .SC_OUT_TOP(scff_Wires[258]),
    .SC_IN_BOT(scff_Wires[257]),
    .chanx_left_in(sb_1__1__96_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__107_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__107_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__107_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__107_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__107_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__107_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__107_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__107_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__107_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__107_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__107_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__107_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__107_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__107_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__107_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__107_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__107_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__107_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__107_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__107_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__107_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[397]),
    .pReset_S_out(pResetWires[541]),
    .pReset_E_out(pResetWires[540]),
    .pReset_W_in(pResetWires[539]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[108]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[108]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[108]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[108]),
    .SC_OUT_TOP(scff_Wires[260]),
    .SC_IN_BOT(scff_Wires[259]),
    .chanx_left_in(sb_1__1__97_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__108_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__108_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__108_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__108_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__108_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__108_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__108_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__108_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__108_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__108_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__108_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__108_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__108_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__108_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__108_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__108_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__108_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__108_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__108_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__108_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__108_ccff_tail[0])
  );


  cbx_1__1_
  cbx_10__11_
  (
    .clk_1_S_out(clk_1_wires[209]),
    .clk_1_N_out(clk_1_wires[208]),
    .clk_1_W_in(clk_1_wires[204]),
    .prog_clk_1_S_out(prog_clk_1_wires[209]),
    .prog_clk_1_N_out(prog_clk_1_wires[208]),
    .prog_clk_1_W_in(prog_clk_1_wires[204]),
    .prog_clk_0_N_in(prog_clk_0_wires[400]),
    .pReset_S_out(pResetWires[590]),
    .pReset_E_out(pResetWires[589]),
    .pReset_W_in(pResetWires[588]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[109]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[109]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[109]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[109]),
    .SC_OUT_TOP(scff_Wires[262]),
    .SC_IN_BOT(scff_Wires[261]),
    .chanx_left_in(sb_1__1__98_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__109_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__109_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__109_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__109_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__109_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__109_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__109_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__109_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__109_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__109_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__109_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__109_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__109_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__109_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__109_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__109_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__109_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__109_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__109_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__109_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__109_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__1_
  (
    .clk_1_S_out(clk_1_wires[214]),
    .clk_1_N_out(clk_1_wires[213]),
    .clk_1_E_in(clk_1_wires[212]),
    .prog_clk_1_S_out(prog_clk_1_wires[214]),
    .prog_clk_1_N_out(prog_clk_1_wires[213]),
    .prog_clk_1_E_in(prog_clk_1_wires[212]),
    .prog_clk_0_N_in(prog_clk_0_wires[408]),
    .pReset_S_out(pResetWires[104]),
    .pReset_E_out(pResetWires[103]),
    .pReset_W_in(pResetWires[102]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[110]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[110]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[110]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[110]),
    .SC_OUT_BOT(scff_Wires[288]),
    .SC_IN_TOP(scff_Wires[287]),
    .chanx_left_in(sb_1__1__99_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__110_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__110_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__110_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__110_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__110_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__110_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__110_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__110_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__110_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__110_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__110_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__110_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__110_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__110_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__110_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__110_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__110_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__110_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__110_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__110_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__110_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__2_
  (
    .clk_2_W_in(clk_2_wires[114]),
    .clk_2_E_out(clk_2_wires[113]),
    .prog_clk_2_W_in(prog_clk_2_wires[114]),
    .prog_clk_2_E_out(prog_clk_2_wires[113]),
    .prog_clk_0_N_in(prog_clk_0_wires[411]),
    .pReset_S_out(pResetWires[153]),
    .pReset_E_out(pResetWires[152]),
    .pReset_W_in(pResetWires[151]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[111]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[111]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[111]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[111]),
    .SC_OUT_BOT(scff_Wires[286]),
    .SC_IN_TOP(scff_Wires[285]),
    .chanx_left_in(sb_1__1__100_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__111_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__111_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__111_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__111_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__111_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__111_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__111_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__111_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__111_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__111_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__111_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__111_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__111_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__111_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__111_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__111_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__111_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__111_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__111_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__111_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__111_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__3_
  (
    .clk_1_S_out(clk_1_wires[221]),
    .clk_1_N_out(clk_1_wires[220]),
    .clk_1_E_in(clk_1_wires[219]),
    .prog_clk_1_S_out(prog_clk_1_wires[221]),
    .prog_clk_1_N_out(prog_clk_1_wires[220]),
    .prog_clk_1_E_in(prog_clk_1_wires[219]),
    .prog_clk_0_N_in(prog_clk_0_wires[414]),
    .pReset_S_out(pResetWires[202]),
    .pReset_E_out(pResetWires[201]),
    .pReset_W_in(pResetWires[200]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[112]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[112]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[112]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[112]),
    .SC_OUT_BOT(scff_Wires[284]),
    .SC_IN_TOP(scff_Wires[283]),
    .chanx_left_in(sb_1__1__101_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__112_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__112_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__112_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__112_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__112_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__112_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__112_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__112_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__112_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__112_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__112_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__112_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__112_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__112_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__112_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__112_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__112_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__112_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__112_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__112_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__112_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__4_
  (
    .clk_2_W_in(clk_2_wires[119]),
    .clk_2_E_out(clk_2_wires[118]),
    .prog_clk_2_W_in(prog_clk_2_wires[119]),
    .prog_clk_2_E_out(prog_clk_2_wires[118]),
    .prog_clk_0_N_in(prog_clk_0_wires[417]),
    .pReset_S_out(pResetWires[251]),
    .pReset_E_out(pResetWires[250]),
    .pReset_W_in(pResetWires[249]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[113]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[113]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[113]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[113]),
    .SC_OUT_BOT(scff_Wires[282]),
    .SC_IN_TOP(scff_Wires[281]),
    .chanx_left_in(sb_1__1__102_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__113_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__113_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__113_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__113_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__113_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__113_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__113_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__113_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__113_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__113_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__113_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__113_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__113_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__113_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__113_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__113_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__113_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__113_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__113_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__113_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__113_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__5_
  (
    .clk_1_S_out(clk_1_wires[228]),
    .clk_1_N_out(clk_1_wires[227]),
    .clk_1_E_in(clk_1_wires[226]),
    .prog_clk_1_S_out(prog_clk_1_wires[228]),
    .prog_clk_1_N_out(prog_clk_1_wires[227]),
    .prog_clk_1_E_in(prog_clk_1_wires[226]),
    .prog_clk_0_N_in(prog_clk_0_wires[420]),
    .pReset_S_out(pResetWires[300]),
    .pReset_E_out(pResetWires[299]),
    .pReset_W_in(pResetWires[298]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[114]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[114]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[114]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[114]),
    .SC_OUT_BOT(scff_Wires[280]),
    .SC_IN_TOP(scff_Wires[279]),
    .chanx_left_in(sb_1__1__103_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__114_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__114_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__114_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__114_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__114_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__114_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__114_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__114_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__114_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__114_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__114_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__114_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__114_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__114_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__114_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__114_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__114_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__114_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__114_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__114_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__114_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[423]),
    .pReset_S_out(pResetWires[349]),
    .pReset_E_out(pResetWires[348]),
    .pReset_W_in(pResetWires[347]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[115]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[115]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[115]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[115]),
    .SC_OUT_BOT(scff_Wires[278]),
    .SC_IN_TOP(scff_Wires[277]),
    .chanx_left_in(sb_1__1__104_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__115_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__115_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__115_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__115_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__115_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__115_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__115_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__115_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__115_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__115_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__115_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__115_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__115_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__115_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__115_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__115_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__115_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__115_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__115_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__115_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__115_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__7_
  (
    .clk_1_S_out(clk_1_wires[235]),
    .clk_1_N_out(clk_1_wires[234]),
    .clk_1_E_in(clk_1_wires[233]),
    .prog_clk_1_S_out(prog_clk_1_wires[235]),
    .prog_clk_1_N_out(prog_clk_1_wires[234]),
    .prog_clk_1_E_in(prog_clk_1_wires[233]),
    .prog_clk_0_N_in(prog_clk_0_wires[426]),
    .pReset_S_out(pResetWires[398]),
    .pReset_E_out(pResetWires[397]),
    .pReset_W_in(pResetWires[396]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[116]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[116]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[116]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[116]),
    .SC_OUT_BOT(scff_Wires[276]),
    .SC_IN_TOP(scff_Wires[275]),
    .chanx_left_in(sb_1__1__105_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__116_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__116_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__116_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__116_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__116_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__116_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__116_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__116_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__116_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__116_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__116_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__116_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__116_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__116_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__116_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__116_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__116_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__116_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__116_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__116_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__116_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__8_
  (
    .clk_2_W_in(clk_2_wires[126]),
    .clk_2_E_out(clk_2_wires[125]),
    .prog_clk_2_W_in(prog_clk_2_wires[126]),
    .prog_clk_2_E_out(prog_clk_2_wires[125]),
    .prog_clk_0_N_in(prog_clk_0_wires[429]),
    .pReset_S_out(pResetWires[447]),
    .pReset_E_out(pResetWires[446]),
    .pReset_W_in(pResetWires[445]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[117]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[117]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[117]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[117]),
    .SC_OUT_BOT(scff_Wires[274]),
    .SC_IN_TOP(scff_Wires[273]),
    .chanx_left_in(sb_1__1__106_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__117_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__117_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__117_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__117_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__117_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__117_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__117_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__117_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__117_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__117_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__117_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__117_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__117_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__117_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__117_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__117_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__117_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__117_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__117_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__117_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__117_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__9_
  (
    .clk_1_S_out(clk_1_wires[242]),
    .clk_1_N_out(clk_1_wires[241]),
    .clk_1_E_in(clk_1_wires[240]),
    .prog_clk_1_S_out(prog_clk_1_wires[242]),
    .prog_clk_1_N_out(prog_clk_1_wires[241]),
    .prog_clk_1_E_in(prog_clk_1_wires[240]),
    .prog_clk_0_N_in(prog_clk_0_wires[432]),
    .pReset_S_out(pResetWires[496]),
    .pReset_E_out(pResetWires[495]),
    .pReset_W_in(pResetWires[494]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[118]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[118]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[118]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[118]),
    .SC_OUT_BOT(scff_Wires[272]),
    .SC_IN_TOP(scff_Wires[271]),
    .chanx_left_in(sb_1__1__107_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__118_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__118_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__118_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__118_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__118_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__118_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__118_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__118_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__118_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__118_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__118_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__118_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__118_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__118_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__118_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__118_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__118_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__118_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__118_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__118_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__118_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__10_
  (
    .clk_2_W_in(clk_2_wires[133]),
    .clk_2_E_out(clk_2_wires[132]),
    .prog_clk_2_W_in(prog_clk_2_wires[133]),
    .prog_clk_2_E_out(prog_clk_2_wires[132]),
    .prog_clk_0_N_in(prog_clk_0_wires[435]),
    .pReset_S_out(pResetWires[545]),
    .pReset_E_out(pResetWires[544]),
    .pReset_W_in(pResetWires[543]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[119]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[119]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[119]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[119]),
    .SC_OUT_BOT(scff_Wires[270]),
    .SC_IN_TOP(scff_Wires[269]),
    .chanx_left_in(sb_1__1__108_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__119_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__119_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__119_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__119_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__119_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__119_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__119_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__119_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__119_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__119_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__119_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__119_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__119_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__119_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__119_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__119_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__119_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__119_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__119_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__119_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__119_ccff_tail[0])
  );


  cbx_1__1_
  cbx_11__11_
  (
    .clk_1_S_out(clk_1_wires[249]),
    .clk_1_N_out(clk_1_wires[248]),
    .clk_1_E_in(clk_1_wires[247]),
    .prog_clk_1_S_out(prog_clk_1_wires[249]),
    .prog_clk_1_N_out(prog_clk_1_wires[248]),
    .prog_clk_1_E_in(prog_clk_1_wires[247]),
    .prog_clk_0_N_in(prog_clk_0_wires[438]),
    .pReset_S_out(pResetWires[594]),
    .pReset_E_out(pResetWires[593]),
    .pReset_W_in(pResetWires[592]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[120]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[120]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[120]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[120]),
    .SC_OUT_BOT(scff_Wires[268]),
    .SC_IN_TOP(scff_Wires[267]),
    .chanx_left_in(sb_1__1__109_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__1__120_chanx_left_out[0:29]),
    .ccff_head(sb_1__1__120_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__120_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__120_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__120_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__120_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__120_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__120_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__120_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__120_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__120_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__120_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__120_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__120_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__120_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__120_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__120_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__120_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__120_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__120_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__120_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__1_
  (
    .clk_1_S_out(clk_1_wires[216]),
    .clk_1_N_out(clk_1_wires[215]),
    .clk_1_W_in(clk_1_wires[211]),
    .prog_clk_1_S_out(prog_clk_1_wires[216]),
    .prog_clk_1_N_out(prog_clk_1_wires[215]),
    .prog_clk_1_W_in(prog_clk_1_wires[211]),
    .prog_clk_0_N_in(prog_clk_0_wires[446]),
    .pReset_S_out(pResetWires[108]),
    .pReset_E_out(pResetWires[107]),
    .pReset_W_in(pResetWires[106]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[121]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[121]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[121]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[121]),
    .SC_OUT_TOP(scff_Wires[295]),
    .SC_IN_BOT(scff_Wires[294]),
    .chanx_left_in(sb_1__1__110_chanx_right_out[0:29]),
    .chanx_right_in(sb_12__1__0_chanx_left_out[0:29]),
    .ccff_head(sb_12__1__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__121_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__121_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__121_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__121_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__121_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__121_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__121_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__121_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__121_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__121_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__121_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__121_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__121_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__121_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__121_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__121_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__121_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__121_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__121_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[449]),
    .pReset_S_out(pResetWires[157]),
    .pReset_E_out(pResetWires[156]),
    .pReset_W_in(pResetWires[155]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[122]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[122]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[122]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[122]),
    .SC_OUT_TOP(scff_Wires[297]),
    .SC_IN_BOT(scff_Wires[296]),
    .chanx_left_in(sb_1__1__111_chanx_right_out[0:29]),
    .chanx_right_in(sb_12__1__1_chanx_left_out[0:29]),
    .ccff_head(sb_12__1__1_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__122_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__122_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__122_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__122_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__122_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__122_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__122_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__122_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__122_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__122_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__122_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__122_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__122_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__122_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__122_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__122_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__122_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__122_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__122_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__3_
  (
    .clk_1_S_out(clk_1_wires[223]),
    .clk_1_N_out(clk_1_wires[222]),
    .clk_1_W_in(clk_1_wires[218]),
    .prog_clk_1_S_out(prog_clk_1_wires[223]),
    .prog_clk_1_N_out(prog_clk_1_wires[222]),
    .prog_clk_1_W_in(prog_clk_1_wires[218]),
    .prog_clk_0_N_in(prog_clk_0_wires[452]),
    .pReset_S_out(pResetWires[206]),
    .pReset_E_out(pResetWires[205]),
    .pReset_W_in(pResetWires[204]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[123]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[123]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[123]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[123]),
    .SC_OUT_TOP(scff_Wires[299]),
    .SC_IN_BOT(scff_Wires[298]),
    .chanx_left_in(sb_1__1__112_chanx_right_out[0:29]),
    .chanx_right_in(sb_12__1__2_chanx_left_out[0:29]),
    .ccff_head(sb_12__1__2_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__123_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__123_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__123_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__123_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__123_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__123_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__123_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__123_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__123_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__123_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__123_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__123_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__123_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__123_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__123_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__123_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__123_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__123_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__123_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[455]),
    .pReset_S_out(pResetWires[255]),
    .pReset_E_out(pResetWires[254]),
    .pReset_W_in(pResetWires[253]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[124]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[124]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[124]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[124]),
    .SC_OUT_TOP(scff_Wires[301]),
    .SC_IN_BOT(scff_Wires[300]),
    .chanx_left_in(sb_1__1__113_chanx_right_out[0:29]),
    .chanx_right_in(sb_12__1__3_chanx_left_out[0:29]),
    .ccff_head(sb_12__1__3_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__124_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__124_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__124_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__124_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__124_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__124_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__124_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__124_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__124_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__124_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__124_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__124_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__124_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__124_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__124_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__124_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__124_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__124_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__124_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__5_
  (
    .clk_1_S_out(clk_1_wires[230]),
    .clk_1_N_out(clk_1_wires[229]),
    .clk_1_W_in(clk_1_wires[225]),
    .prog_clk_1_S_out(prog_clk_1_wires[230]),
    .prog_clk_1_N_out(prog_clk_1_wires[229]),
    .prog_clk_1_W_in(prog_clk_1_wires[225]),
    .prog_clk_0_N_in(prog_clk_0_wires[458]),
    .pReset_S_out(pResetWires[304]),
    .pReset_E_out(pResetWires[303]),
    .pReset_W_in(pResetWires[302]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[125]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[125]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[125]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[125]),
    .SC_OUT_TOP(scff_Wires[303]),
    .SC_IN_BOT(scff_Wires[302]),
    .chanx_left_in(sb_1__1__114_chanx_right_out[0:29]),
    .chanx_right_in(sb_12__1__4_chanx_left_out[0:29]),
    .ccff_head(sb_12__1__4_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__125_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__125_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__125_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__125_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__125_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__125_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__125_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__125_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__125_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__125_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__125_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__125_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__125_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__125_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__125_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__125_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__125_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__125_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__125_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[461]),
    .pReset_S_out(pResetWires[353]),
    .pReset_E_out(pResetWires[352]),
    .pReset_W_in(pResetWires[351]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[126]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[126]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[126]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[126]),
    .SC_OUT_TOP(scff_Wires[305]),
    .SC_IN_BOT(scff_Wires[304]),
    .chanx_left_in(sb_1__1__115_chanx_right_out[0:29]),
    .chanx_right_in(sb_12__1__5_chanx_left_out[0:29]),
    .ccff_head(sb_12__1__5_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__126_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__126_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__126_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__126_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__126_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__126_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__126_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__126_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__126_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__126_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__126_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__126_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__126_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__126_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__126_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__126_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__126_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__126_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__126_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__7_
  (
    .clk_1_S_out(clk_1_wires[237]),
    .clk_1_N_out(clk_1_wires[236]),
    .clk_1_W_in(clk_1_wires[232]),
    .prog_clk_1_S_out(prog_clk_1_wires[237]),
    .prog_clk_1_N_out(prog_clk_1_wires[236]),
    .prog_clk_1_W_in(prog_clk_1_wires[232]),
    .prog_clk_0_N_in(prog_clk_0_wires[464]),
    .pReset_S_out(pResetWires[402]),
    .pReset_E_out(pResetWires[401]),
    .pReset_W_in(pResetWires[400]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[127]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[127]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[127]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[127]),
    .SC_OUT_TOP(scff_Wires[307]),
    .SC_IN_BOT(scff_Wires[306]),
    .chanx_left_in(sb_1__1__116_chanx_right_out[0:29]),
    .chanx_right_in(sb_12__1__6_chanx_left_out[0:29]),
    .ccff_head(sb_12__1__6_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__127_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__127_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__127_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__127_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__127_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__127_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__127_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__127_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__127_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__127_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__127_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__127_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__127_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__127_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__127_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__127_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__127_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__127_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__127_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__8_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[467]),
    .pReset_S_out(pResetWires[451]),
    .pReset_E_out(pResetWires[450]),
    .pReset_W_in(pResetWires[449]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[128]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[128]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[128]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[128]),
    .SC_OUT_TOP(scff_Wires[309]),
    .SC_IN_BOT(scff_Wires[308]),
    .chanx_left_in(sb_1__1__117_chanx_right_out[0:29]),
    .chanx_right_in(sb_12__1__7_chanx_left_out[0:29]),
    .ccff_head(sb_12__1__7_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__128_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__128_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__128_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__128_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__128_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__128_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__128_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__128_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__128_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__128_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__128_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__128_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__128_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__128_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__128_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__128_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__128_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__128_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__128_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__9_
  (
    .clk_1_S_out(clk_1_wires[244]),
    .clk_1_N_out(clk_1_wires[243]),
    .clk_1_W_in(clk_1_wires[239]),
    .prog_clk_1_S_out(prog_clk_1_wires[244]),
    .prog_clk_1_N_out(prog_clk_1_wires[243]),
    .prog_clk_1_W_in(prog_clk_1_wires[239]),
    .prog_clk_0_N_in(prog_clk_0_wires[470]),
    .pReset_S_out(pResetWires[500]),
    .pReset_E_out(pResetWires[499]),
    .pReset_W_in(pResetWires[498]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[129]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[129]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[129]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[129]),
    .SC_OUT_TOP(scff_Wires[311]),
    .SC_IN_BOT(scff_Wires[310]),
    .chanx_left_in(sb_1__1__118_chanx_right_out[0:29]),
    .chanx_right_in(sb_12__1__8_chanx_left_out[0:29]),
    .ccff_head(sb_12__1__8_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__129_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__129_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__129_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__129_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__129_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__129_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__129_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__129_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__129_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__129_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__129_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__129_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__129_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__129_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__129_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__129_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__129_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__129_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__129_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__10_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[473]),
    .pReset_S_out(pResetWires[549]),
    .pReset_E_out(pResetWires[548]),
    .pReset_W_in(pResetWires[547]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[130]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[130]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[130]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[130]),
    .SC_OUT_TOP(scff_Wires[313]),
    .SC_IN_BOT(scff_Wires[312]),
    .chanx_left_in(sb_1__1__119_chanx_right_out[0:29]),
    .chanx_right_in(sb_12__1__9_chanx_left_out[0:29]),
    .ccff_head(sb_12__1__9_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__130_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__130_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__130_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__130_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__130_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__130_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__130_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__130_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__130_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__130_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__130_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__130_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__130_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__130_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__130_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__130_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__130_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__130_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__130_ccff_tail[0])
  );


  cbx_1__1_
  cbx_12__11_
  (
    .clk_1_S_out(clk_1_wires[251]),
    .clk_1_N_out(clk_1_wires[250]),
    .clk_1_W_in(clk_1_wires[246]),
    .prog_clk_1_S_out(prog_clk_1_wires[251]),
    .prog_clk_1_N_out(prog_clk_1_wires[250]),
    .prog_clk_1_W_in(prog_clk_1_wires[246]),
    .prog_clk_0_N_in(prog_clk_0_wires[476]),
    .pReset_S_out(pResetWires[598]),
    .pReset_E_out(pResetWires[597]),
    .pReset_W_in(pResetWires[596]),
    .COUT_FEEDTHROUGH(cout_feedthrough_wires[131]),
    .CIN_FEEDTHROUGH(cin_feedthrough_wires[131]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[131]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[131]),
    .SC_OUT_TOP(scff_Wires[315]),
    .SC_IN_BOT(scff_Wires[314]),
    .chanx_left_in(sb_1__1__120_chanx_right_out[0:29]),
    .chanx_right_in(sb_12__1__10_chanx_left_out[0:29]),
    .ccff_head(sb_12__1__10_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__131_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__1__131_chanx_right_out[0:29]),
    .bottom_grid_pin_0_(cbx_1__1__131_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__131_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__131_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__131_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__131_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__131_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__131_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__131_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__131_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__131_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__131_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__131_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__131_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__131_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__131_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__131_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__131_ccff_tail[0])
  );


  cbx_1__2_
  cbx_1__12_
  (
    .prog_clk_0_W_out(prog_clk_0_wires[62]),
    .prog_clk_0_S_in(prog_clk_0_wires[59]),
    .pReset_S_out(pResetWires[602]),
    .pReset_E_in(pResetWires[601]),
    .pReset_W_out(pResetWires[600]),
    .SC_OUT_BOT(scff_Wires[1]),
    .SC_IN_TOP(scff_Wires[0]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_0_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_0_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__0_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_0__12__0_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__12__0_chanx_left_out[0:29]),
    .ccff_head(sb_1__12__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__0_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__12__0_chanx_right_out[0:29]),
    .top_grid_pin_0_(cbx_1__12__0_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__0_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__0_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__0_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__0_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__0_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__0_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__0_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__0_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__0_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__0_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__0_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__0_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__0_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__0_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__0_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__0_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_0_ccff_tail[0])
  );


  cbx_1__2_
  cbx_2__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[99]),
    .pReset_S_out(pResetWires[606]),
    .pReset_E_in(pResetWires[605]),
    .pReset_W_out(pResetWires[604]),
    .SC_OUT_TOP(scff_Wires[52]),
    .SC_IN_BOT(scff_Wires[51]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_1_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_1_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__1_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__0_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__12__1_chanx_left_out[0:29]),
    .ccff_head(sb_1__12__1_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__1_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__12__1_chanx_right_out[0:29]),
    .top_grid_pin_0_(cbx_1__12__1_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__1_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__1_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__1_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__1_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__1_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__1_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__1_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__1_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__1_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__1_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__1_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__1_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__1_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__1_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__1_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__1_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_1_ccff_tail[0])
  );


  cbx_1__2_
  cbx_3__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[137]),
    .pReset_S_out(pResetWires[609]),
    .pReset_E_in(pResetWires[608]),
    .pReset_W_out(pResetWires[607]),
    .SC_OUT_BOT(scff_Wires[54]),
    .SC_IN_TOP(scff_Wires[53]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_2_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_2_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__2_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__1_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__12__2_chanx_left_out[0:29]),
    .ccff_head(sb_1__12__2_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__2_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__12__2_chanx_right_out[0:29]),
    .top_grid_pin_0_(cbx_1__12__2_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__2_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__2_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__2_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__2_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__2_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__2_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__2_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__2_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__2_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__2_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__2_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__2_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__2_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__2_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__2_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__2_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_2_ccff_tail[0])
  );


  cbx_1__2_
  cbx_4__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[175]),
    .pReset_S_out(pResetWires[612]),
    .pReset_E_in(pResetWires[611]),
    .pReset_W_out(pResetWires[610]),
    .SC_OUT_TOP(scff_Wires[105]),
    .SC_IN_BOT(scff_Wires[104]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_3_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_3_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__3_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__2_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__12__3_chanx_left_out[0:29]),
    .ccff_head(sb_1__12__3_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__3_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__12__3_chanx_right_out[0:29]),
    .top_grid_pin_0_(cbx_1__12__3_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__3_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__3_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__3_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__3_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__3_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__3_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__3_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__3_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__3_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__3_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__3_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__3_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__3_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__3_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__3_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__3_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_3_ccff_tail[0])
  );


  cbx_1__2_
  cbx_5__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[213]),
    .pReset_S_out(pResetWires[615]),
    .pReset_E_in(pResetWires[614]),
    .pReset_W_out(pResetWires[613]),
    .SC_OUT_BOT(scff_Wires[107]),
    .SC_IN_TOP(scff_Wires[106]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_4_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_4_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__4_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__3_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__12__4_chanx_left_out[0:29]),
    .ccff_head(sb_1__12__4_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__4_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__12__4_chanx_right_out[0:29]),
    .top_grid_pin_0_(cbx_1__12__4_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__4_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__4_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__4_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__4_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__4_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__4_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__4_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__4_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__4_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__4_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__4_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__4_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__4_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__4_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__4_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__4_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_4_ccff_tail[0])
  );


  cbx_1__2_
  cbx_6__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[251]),
    .pReset_S_out(pResetWires[618]),
    .pReset_E_in(pResetWires[617]),
    .pReset_W_out(pResetWires[616]),
    .SC_OUT_TOP(scff_Wires[158]),
    .SC_IN_BOT(scff_Wires[157]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_5_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_5_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__5_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__4_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__12__5_chanx_left_out[0:29]),
    .ccff_head(sb_1__12__5_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__5_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__12__5_chanx_right_out[0:29]),
    .top_grid_pin_0_(cbx_1__12__5_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__5_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__5_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__5_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__5_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__5_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__5_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__5_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__5_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__5_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__5_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__5_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__5_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__5_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__5_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__5_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__5_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_5_ccff_tail[0])
  );


  cbx_1__2_
  cbx_7__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[289]),
    .pReset_S_out(pResetWires[621]),
    .pReset_E_out(pResetWires[620]),
    .pReset_W_in(pResetWires[619]),
    .SC_OUT_BOT(scff_Wires[160]),
    .SC_IN_TOP(scff_Wires[159]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_6_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_6_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__6_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__5_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__12__6_chanx_left_out[0:29]),
    .ccff_head(sb_1__12__6_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__6_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__12__6_chanx_right_out[0:29]),
    .top_grid_pin_0_(cbx_1__12__6_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__6_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__6_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__6_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__6_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__6_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__6_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__6_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__6_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__6_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__6_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__6_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__6_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__6_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__6_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__6_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__6_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_6_ccff_tail[0])
  );


  cbx_1__2_
  cbx_8__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[327]),
    .pReset_S_out(pResetWires[624]),
    .pReset_E_out(pResetWires[623]),
    .pReset_W_in(pResetWires[622]),
    .SC_OUT_TOP(scff_Wires[211]),
    .SC_IN_BOT(scff_Wires[210]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_7_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_7_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__7_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__6_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__12__7_chanx_left_out[0:29]),
    .ccff_head(sb_1__12__7_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__7_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__12__7_chanx_right_out[0:29]),
    .top_grid_pin_0_(cbx_1__12__7_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__7_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__7_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__7_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__7_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__7_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__7_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__7_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__7_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__7_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__7_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__7_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__7_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__7_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__7_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__7_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__7_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_7_ccff_tail[0])
  );


  cbx_1__2_
  cbx_9__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[365]),
    .pReset_S_out(pResetWires[627]),
    .pReset_E_out(pResetWires[626]),
    .pReset_W_in(pResetWires[625]),
    .SC_OUT_BOT(scff_Wires[213]),
    .SC_IN_TOP(scff_Wires[212]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_8_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_8_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__8_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__7_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__12__8_chanx_left_out[0:29]),
    .ccff_head(sb_1__12__8_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__8_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__12__8_chanx_right_out[0:29]),
    .top_grid_pin_0_(cbx_1__12__8_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__8_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__8_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__8_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__8_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__8_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__8_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__8_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__8_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__8_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__8_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__8_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__8_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__8_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__8_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__8_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__8_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_8_ccff_tail[0])
  );


  cbx_1__2_
  cbx_10__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[403]),
    .pReset_S_out(pResetWires[630]),
    .pReset_E_out(pResetWires[629]),
    .pReset_W_in(pResetWires[628]),
    .SC_OUT_TOP(scff_Wires[264]),
    .SC_IN_BOT(scff_Wires[263]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_9_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_9_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__9_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__8_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__12__9_chanx_left_out[0:29]),
    .ccff_head(sb_1__12__9_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__9_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__12__9_chanx_right_out[0:29]),
    .top_grid_pin_0_(cbx_1__12__9_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__9_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__9_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__9_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__9_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__9_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__9_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__9_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__9_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__9_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__9_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__9_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__9_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__9_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__9_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__9_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__9_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_9_ccff_tail[0])
  );


  cbx_1__2_
  cbx_11__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[441]),
    .pReset_S_out(pResetWires[633]),
    .pReset_E_out(pResetWires[632]),
    .pReset_W_in(pResetWires[631]),
    .SC_OUT_BOT(scff_Wires[266]),
    .SC_IN_TOP(scff_Wires[265]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_10_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_10_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__10_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__9_chanx_right_out[0:29]),
    .chanx_right_in(sb_1__12__10_chanx_left_out[0:29]),
    .ccff_head(sb_1__12__10_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__10_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__12__10_chanx_right_out[0:29]),
    .top_grid_pin_0_(cbx_1__12__10_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__10_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__10_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__10_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__10_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__10_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__10_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__10_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__10_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__10_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__10_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__10_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__10_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__10_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__10_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__10_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__10_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_10_ccff_tail[0])
  );


  cbx_1__2_
  cbx_12__12_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[479]),
    .pReset_S_out(pResetWires[636]),
    .pReset_E_out(pResetWires[635]),
    .pReset_W_in(pResetWires[634]),
    .SC_OUT_TOP(scff_Wires[317]),
    .SC_IN_BOT(scff_Wires[316]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_11_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_11_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__12__11_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__12__10_chanx_right_out[0:29]),
    .chanx_right_in(sb_12__12__0_chanx_left_out[0:29]),
    .ccff_head(sb_12__12__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__12__11_chanx_left_out[0:29]),
    .chanx_right_out(cbx_1__12__11_chanx_right_out[0:29]),
    .top_grid_pin_0_(cbx_1__12__11_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__12__11_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__12__11_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__12__11_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__12__11_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__12__11_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__12__11_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__12__11_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__12__11_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__12__11_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__12__11_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__12__11_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__12__11_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__12__11_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__12__11_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__12__11_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__12__11_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_11_ccff_tail[0])
  );


  cby_0__1_
  cby_0__1_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[3]),
    .pReset_N_in(pResetWires[64]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_0_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_0_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__0_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[132]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[132]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[132]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__0__0_chany_top_out[0:29]),
    .chany_top_in(sb_0__1__0_chany_bottom_out[0:29]),
    .ccff_head(sb_0__1__0_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__0_chany_bottom_out[0:29]),
    .chany_top_out(cby_0__1__0_chany_top_out[0:29]),
    .left_grid_pin_0_(cby_0__1__0_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_0_ccff_tail[0])
  );


  cby_0__1_
  cby_0__2_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[9]),
    .pReset_N_in(pResetWires[113]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_1_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_1_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__1_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[133]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[133]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[133]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__0_chany_top_out[0:29]),
    .chany_top_in(sb_0__1__1_chany_bottom_out[0:29]),
    .ccff_head(sb_0__1__1_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__1_chany_bottom_out[0:29]),
    .chany_top_out(cby_0__1__1_chany_top_out[0:29]),
    .left_grid_pin_0_(cby_0__1__1_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_1_ccff_tail[0])
  );


  cby_0__1_
  cby_0__3_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[14]),
    .pReset_N_in(pResetWires[162]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_2_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_2_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__2_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[134]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[134]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[134]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__1_chany_top_out[0:29]),
    .chany_top_in(sb_0__1__2_chany_bottom_out[0:29]),
    .ccff_head(sb_0__1__2_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__2_chany_bottom_out[0:29]),
    .chany_top_out(cby_0__1__2_chany_top_out[0:29]),
    .left_grid_pin_0_(cby_0__1__2_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_2_ccff_tail[0])
  );


  cby_0__1_
  cby_0__4_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[19]),
    .pReset_N_in(pResetWires[211]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_3_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_3_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__3_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[135]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[135]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[135]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__2_chany_top_out[0:29]),
    .chany_top_in(sb_0__1__3_chany_bottom_out[0:29]),
    .ccff_head(sb_0__1__3_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__3_chany_bottom_out[0:29]),
    .chany_top_out(cby_0__1__3_chany_top_out[0:29]),
    .left_grid_pin_0_(cby_0__1__3_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_3_ccff_tail[0])
  );


  cby_0__1_
  cby_0__5_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[24]),
    .pReset_N_in(pResetWires[260]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_4_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_4_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__4_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[136]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[136]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[136]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__3_chany_top_out[0:29]),
    .chany_top_in(sb_0__1__4_chany_bottom_out[0:29]),
    .ccff_head(sb_0__1__4_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__4_chany_bottom_out[0:29]),
    .chany_top_out(cby_0__1__4_chany_top_out[0:29]),
    .left_grid_pin_0_(cby_0__1__4_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_4_ccff_tail[0])
  );


  cby_0__1_
  cby_0__6_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[29]),
    .pReset_N_in(pResetWires[309]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_5_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_5_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__5_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[137]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[137]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[137]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__4_chany_top_out[0:29]),
    .chany_top_in(sb_0__1__5_chany_bottom_out[0:29]),
    .ccff_head(sb_0__1__5_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__5_chany_bottom_out[0:29]),
    .chany_top_out(cby_0__1__5_chany_top_out[0:29]),
    .left_grid_pin_0_(cby_0__1__5_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_5_ccff_tail[0])
  );


  cby_0__1_
  cby_0__7_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[34]),
    .pReset_N_in(pResetWires[358]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_6_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_6_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__6_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[138]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[138]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[138]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__5_chany_top_out[0:29]),
    .chany_top_in(sb_0__1__6_chany_bottom_out[0:29]),
    .ccff_head(sb_0__1__6_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__6_chany_bottom_out[0:29]),
    .chany_top_out(cby_0__1__6_chany_top_out[0:29]),
    .left_grid_pin_0_(cby_0__1__6_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_6_ccff_tail[0])
  );


  cby_0__1_
  cby_0__8_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[39]),
    .pReset_N_in(pResetWires[407]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_7_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_7_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__7_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[139]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[139]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[139]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__6_chany_top_out[0:29]),
    .chany_top_in(sb_0__1__7_chany_bottom_out[0:29]),
    .ccff_head(sb_0__1__7_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__7_chany_bottom_out[0:29]),
    .chany_top_out(cby_0__1__7_chany_top_out[0:29]),
    .left_grid_pin_0_(cby_0__1__7_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_7_ccff_tail[0])
  );


  cby_0__1_
  cby_0__9_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[44]),
    .pReset_N_in(pResetWires[456]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_8_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_8_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__8_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[140]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[140]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[140]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__7_chany_top_out[0:29]),
    .chany_top_in(sb_0__1__8_chany_bottom_out[0:29]),
    .ccff_head(sb_0__1__8_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__8_chany_bottom_out[0:29]),
    .chany_top_out(cby_0__1__8_chany_top_out[0:29]),
    .left_grid_pin_0_(cby_0__1__8_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_8_ccff_tail[0])
  );


  cby_0__1_
  cby_0__10_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[49]),
    .pReset_N_in(pResetWires[505]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_9_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_9_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__9_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[141]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[141]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[141]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__8_chany_top_out[0:29]),
    .chany_top_in(sb_0__1__9_chany_bottom_out[0:29]),
    .ccff_head(sb_0__1__9_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__9_chany_bottom_out[0:29]),
    .chany_top_out(cby_0__1__9_chany_top_out[0:29]),
    .left_grid_pin_0_(cby_0__1__9_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_9_ccff_tail[0])
  );


  cby_0__1_
  cby_0__11_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[54]),
    .pReset_N_in(pResetWires[554]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_10_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_10_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__10_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[142]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[142]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[142]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__9_chany_top_out[0:29]),
    .chany_top_in(sb_0__1__10_chany_bottom_out[0:29]),
    .ccff_head(sb_0__1__10_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__10_chany_bottom_out[0:29]),
    .chany_top_out(cby_0__1__10_chany_top_out[0:29]),
    .left_grid_pin_0_(cby_0__1__10_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_10_ccff_tail[0])
  );


  cby_0__1_
  cby_0__12_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[61]),
    .pReset_N_in(pResetWires[603]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_11_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_11_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__11_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[143]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[143]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[143]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__10_chany_top_out[0:29]),
    .chany_top_in(sb_0__12__0_chany_bottom_out[0:29]),
    .ccff_head(sb_0__12__0_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__11_chany_bottom_out[0:29]),
    .chany_top_out(cby_0__1__11_chany_top_out[0:29]),
    .left_grid_pin_0_(cby_0__1__11_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_11_ccff_tail[0])
  );


  cby_1__1_
  cby_1__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[2]),
    .prog_clk_0_W_in(prog_clk_0_wires[1]),
    .Reset_E_in(ResetWires[26]),
    .Reset_W_out(ResetWires[24]),
    .pReset_S_in(pResetWires[27]),
    .Test_en_E_in(Test_enWires[26]),
    .Test_en_W_out(Test_enWires[24]),
    .chany_bottom_in(sb_1__0__0_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__0_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_0_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__0_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__0_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__0_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__0_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__0_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__0_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__0_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__0_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__0_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__0_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__0_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__0_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__0_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__0_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__0_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__0_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__0_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__0_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__0_ccff_tail[0])
  );


  cby_1__1_
  cby_1__2_
  (
    .clk_2_S_out(clk_2_wires[4]),
    .clk_2_N_in(clk_2_wires[3]),
    .prog_clk_2_S_out(prog_clk_2_wires[4]),
    .prog_clk_2_N_in(prog_clk_2_wires[3]),
    .prog_clk_0_S_out(prog_clk_0_wires[8]),
    .prog_clk_0_W_in(prog_clk_0_wires[7]),
    .Reset_E_in(ResetWires[48]),
    .Reset_W_out(ResetWires[46]),
    .pReset_S_in(pResetWires[65]),
    .Test_en_E_in(Test_enWires[48]),
    .Test_en_W_out(Test_enWires[46]),
    .chany_bottom_in(sb_1__1__0_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__1_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_1_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__1_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__1_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__1_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__1_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__1_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__1_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__1_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__1_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__1_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__1_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__1_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__1_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__1_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__1_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__1_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__1_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__1_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__1_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__1_ccff_tail[0])
  );


  cby_1__1_
  cby_1__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[13]),
    .prog_clk_0_W_in(prog_clk_0_wires[12]),
    .Reset_E_in(ResetWires[70]),
    .Reset_W_out(ResetWires[68]),
    .pReset_S_in(pResetWires[114]),
    .Test_en_E_in(Test_enWires[70]),
    .Test_en_W_out(Test_enWires[68]),
    .chany_bottom_in(sb_1__1__1_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__2_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_2_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__2_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__2_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__2_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__2_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__2_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__2_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__2_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__2_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__2_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__2_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__2_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__2_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__2_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__2_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__2_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__2_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__2_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__2_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__2_ccff_tail[0])
  );


  cby_1__1_
  cby_1__4_
  (
    .clk_2_S_out(clk_2_wires[11]),
    .clk_2_N_in(clk_2_wires[10]),
    .prog_clk_2_S_out(prog_clk_2_wires[11]),
    .prog_clk_2_N_in(prog_clk_2_wires[10]),
    .prog_clk_0_S_out(prog_clk_0_wires[18]),
    .prog_clk_0_W_in(prog_clk_0_wires[17]),
    .Reset_E_in(ResetWires[92]),
    .Reset_W_out(ResetWires[90]),
    .pReset_S_in(pResetWires[163]),
    .Test_en_E_in(Test_enWires[92]),
    .Test_en_W_out(Test_enWires[90]),
    .chany_bottom_in(sb_1__1__2_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__3_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_3_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__3_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__3_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__3_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__3_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__3_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__3_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__3_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__3_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__3_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__3_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__3_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__3_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__3_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__3_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__3_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__3_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__3_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__3_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__3_ccff_tail[0])
  );


  cby_1__1_
  cby_1__5_
  (
    .clk_2_N_out(clk_2_wires[9]),
    .clk_2_S_in(clk_2_wires[8]),
    .prog_clk_2_N_out(prog_clk_2_wires[9]),
    .prog_clk_2_S_in(prog_clk_2_wires[8]),
    .prog_clk_0_S_out(prog_clk_0_wires[23]),
    .prog_clk_0_W_in(prog_clk_0_wires[22]),
    .Reset_E_in(ResetWires[114]),
    .Reset_W_out(ResetWires[112]),
    .pReset_S_in(pResetWires[212]),
    .Test_en_E_in(Test_enWires[114]),
    .Test_en_W_out(Test_enWires[112]),
    .chany_bottom_in(sb_1__1__3_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__4_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_4_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__4_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__4_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__4_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__4_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__4_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__4_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__4_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__4_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__4_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__4_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__4_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__4_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__4_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__4_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__4_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__4_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__4_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__4_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__4_ccff_tail[0])
  );


  cby_1__1_
  cby_1__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[28]),
    .prog_clk_0_W_in(prog_clk_0_wires[27]),
    .Reset_E_in(ResetWires[136]),
    .Reset_W_out(ResetWires[134]),
    .pReset_S_in(pResetWires[261]),
    .Test_en_E_in(Test_enWires[136]),
    .Test_en_W_out(Test_enWires[134]),
    .chany_bottom_in(sb_1__1__4_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__5_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_5_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__5_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__5_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__5_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__5_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__5_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__5_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__5_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__5_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__5_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__5_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__5_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__5_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__5_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__5_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__5_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__5_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__5_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__5_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__5_ccff_tail[0])
  );


  cby_1__1_
  cby_1__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[33]),
    .prog_clk_0_W_in(prog_clk_0_wires[32]),
    .Reset_E_in(ResetWires[158]),
    .Reset_W_out(ResetWires[156]),
    .pReset_S_in(pResetWires[310]),
    .Test_en_E_in(Test_enWires[158]),
    .Test_en_W_out(Test_enWires[156]),
    .chany_bottom_in(sb_1__1__5_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__6_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_6_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__6_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__6_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__6_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__6_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__6_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__6_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__6_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__6_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__6_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__6_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__6_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__6_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__6_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__6_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__6_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__6_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__6_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__6_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__6_ccff_tail[0])
  );


  cby_1__1_
  cby_1__8_
  (
    .clk_2_S_out(clk_2_wires[18]),
    .clk_2_N_in(clk_2_wires[17]),
    .prog_clk_2_S_out(prog_clk_2_wires[18]),
    .prog_clk_2_N_in(prog_clk_2_wires[17]),
    .prog_clk_0_S_out(prog_clk_0_wires[38]),
    .prog_clk_0_W_in(prog_clk_0_wires[37]),
    .Reset_E_in(ResetWires[180]),
    .Reset_W_out(ResetWires[178]),
    .pReset_S_in(pResetWires[359]),
    .Test_en_E_in(Test_enWires[180]),
    .Test_en_W_out(Test_enWires[178]),
    .chany_bottom_in(sb_1__1__6_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__7_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_7_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__7_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__7_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__7_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__7_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__7_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__7_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__7_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__7_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__7_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__7_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__7_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__7_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__7_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__7_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__7_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__7_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__7_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__7_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__7_ccff_tail[0])
  );


  cby_1__1_
  cby_1__9_
  (
    .clk_2_N_out(clk_2_wires[16]),
    .clk_2_S_in(clk_2_wires[15]),
    .prog_clk_2_N_out(prog_clk_2_wires[16]),
    .prog_clk_2_S_in(prog_clk_2_wires[15]),
    .prog_clk_0_S_out(prog_clk_0_wires[43]),
    .prog_clk_0_W_in(prog_clk_0_wires[42]),
    .Reset_E_in(ResetWires[202]),
    .Reset_W_out(ResetWires[200]),
    .pReset_S_in(pResetWires[408]),
    .Test_en_E_in(Test_enWires[202]),
    .Test_en_W_out(Test_enWires[200]),
    .chany_bottom_in(sb_1__1__7_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__8_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_8_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__8_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__8_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__8_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__8_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__8_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__8_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__8_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__8_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__8_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__8_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__8_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__8_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__8_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__8_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__8_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__8_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__8_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__8_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__8_ccff_tail[0])
  );


  cby_1__1_
  cby_1__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[48]),
    .prog_clk_0_W_in(prog_clk_0_wires[47]),
    .Reset_E_in(ResetWires[224]),
    .Reset_W_out(ResetWires[222]),
    .pReset_S_in(pResetWires[457]),
    .Test_en_E_in(Test_enWires[224]),
    .Test_en_W_out(Test_enWires[222]),
    .chany_bottom_in(sb_1__1__8_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__9_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_9_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__9_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__9_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__9_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__9_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__9_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__9_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__9_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__9_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__9_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__9_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__9_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__9_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__9_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__9_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__9_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__9_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__9_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__9_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__9_ccff_tail[0])
  );


  cby_1__1_
  cby_1__11_
  (
    .clk_2_N_out(clk_2_wires[23]),
    .clk_2_S_in(clk_2_wires[22]),
    .prog_clk_2_N_out(prog_clk_2_wires[23]),
    .prog_clk_2_S_in(prog_clk_2_wires[22]),
    .prog_clk_0_S_out(prog_clk_0_wires[53]),
    .prog_clk_0_W_in(prog_clk_0_wires[52]),
    .Reset_E_in(ResetWires[246]),
    .Reset_W_out(ResetWires[244]),
    .pReset_S_in(pResetWires[506]),
    .Test_en_E_in(Test_enWires[246]),
    .Test_en_W_out(Test_enWires[244]),
    .chany_bottom_in(sb_1__1__9_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__10_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_10_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__10_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__10_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__10_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__10_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__10_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__10_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__10_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__10_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__10_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__10_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__10_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__10_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__10_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__10_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__10_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__10_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__10_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__10_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__10_ccff_tail[0])
  );


  cby_1__1_
  cby_1__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[60]),
    .prog_clk_0_S_out(prog_clk_0_wires[58]),
    .prog_clk_0_W_in(prog_clk_0_wires[57]),
    .Reset_E_in(ResetWires[268]),
    .Reset_W_out(ResetWires[266]),
    .pReset_S_in(pResetWires[555]),
    .Test_en_E_in(Test_enWires[268]),
    .Test_en_W_out(Test_enWires[266]),
    .chany_bottom_in(sb_1__1__10_chany_top_out[0:29]),
    .chany_top_in(sb_1__12__0_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_11_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__11_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__11_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__11_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__11_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__11_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__11_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__11_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__11_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__11_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__11_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__11_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__11_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__11_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__11_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__11_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__11_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__11_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__11_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__11_ccff_tail[0])
  );


  cby_1__1_
  cby_2__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[65]),
    .prog_clk_0_W_in(prog_clk_0_wires[64]),
    .Reset_E_in(ResetWires[28]),
    .Reset_W_out(ResetWires[25]),
    .pReset_S_in(pResetWires[30]),
    .Test_en_E_in(Test_enWires[28]),
    .Test_en_W_out(Test_enWires[25]),
    .chany_bottom_in(sb_1__0__1_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__11_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_12_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__12_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__12_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__12_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__12_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__12_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__12_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__12_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__12_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__12_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__12_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__12_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__12_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__12_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__12_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__12_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__12_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__12_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__12_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__12_ccff_tail[0])
  );


  cby_1__1_
  cby_2__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[68]),
    .prog_clk_0_W_in(prog_clk_0_wires[67]),
    .Reset_E_in(ResetWires[50]),
    .Reset_W_out(ResetWires[47]),
    .pReset_S_in(pResetWires[69]),
    .Test_en_E_in(Test_enWires[50]),
    .Test_en_W_out(Test_enWires[47]),
    .chany_bottom_in(sb_1__1__11_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__12_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_13_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__13_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__13_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__13_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__13_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__13_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__13_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__13_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__13_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__13_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__13_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__13_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__13_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__13_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__13_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__13_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__13_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__13_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__13_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__13_ccff_tail[0])
  );


  cby_1__1_
  cby_2__3_
  (
    .clk_3_S_out(clk_3_wires[69]),
    .clk_3_N_in(clk_3_wires[68]),
    .prog_clk_3_S_out(prog_clk_3_wires[69]),
    .prog_clk_3_N_in(prog_clk_3_wires[68]),
    .prog_clk_0_S_out(prog_clk_0_wires[71]),
    .prog_clk_0_W_in(prog_clk_0_wires[70]),
    .Reset_E_in(ResetWires[72]),
    .Reset_W_out(ResetWires[69]),
    .pReset_S_in(pResetWires[118]),
    .Test_en_E_in(Test_enWires[72]),
    .Test_en_W_out(Test_enWires[69]),
    .chany_bottom_in(sb_1__1__12_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__13_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_14_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__14_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__14_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__14_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__14_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__14_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__14_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__14_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__14_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__14_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__14_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__14_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__14_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__14_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__14_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__14_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__14_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__14_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__14_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__14_ccff_tail[0])
  );


  cby_1__1_
  cby_2__4_
  (
    .clk_3_S_out(clk_3_wires[65]),
    .clk_3_N_in(clk_3_wires[64]),
    .prog_clk_3_S_out(prog_clk_3_wires[65]),
    .prog_clk_3_N_in(prog_clk_3_wires[64]),
    .prog_clk_0_S_out(prog_clk_0_wires[74]),
    .prog_clk_0_W_in(prog_clk_0_wires[73]),
    .Reset_E_in(ResetWires[94]),
    .Reset_W_out(ResetWires[91]),
    .pReset_S_in(pResetWires[167]),
    .Test_en_E_in(Test_enWires[94]),
    .Test_en_W_out(Test_enWires[91]),
    .chany_bottom_in(sb_1__1__13_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__14_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_15_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__15_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__15_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__15_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__15_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__15_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__15_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__15_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__15_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__15_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__15_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__15_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__15_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__15_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__15_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__15_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__15_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__15_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__15_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__15_ccff_tail[0])
  );


  cby_1__1_
  cby_2__5_
  (
    .clk_3_S_out(clk_3_wires[59]),
    .clk_3_N_in(clk_3_wires[58]),
    .prog_clk_3_S_out(prog_clk_3_wires[59]),
    .prog_clk_3_N_in(prog_clk_3_wires[58]),
    .prog_clk_0_S_out(prog_clk_0_wires[77]),
    .prog_clk_0_W_in(prog_clk_0_wires[76]),
    .Reset_E_in(ResetWires[116]),
    .Reset_W_out(ResetWires[113]),
    .pReset_S_in(pResetWires[216]),
    .Test_en_E_in(Test_enWires[116]),
    .Test_en_W_out(Test_enWires[113]),
    .chany_bottom_in(sb_1__1__14_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__15_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_16_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__16_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__16_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__16_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__16_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__16_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__16_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__16_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__16_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__16_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__16_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__16_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__16_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__16_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__16_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__16_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__16_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__16_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__16_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__16_ccff_tail[0])
  );


  cby_1__1_
  cby_2__6_
  (
    .clk_3_S_out(clk_3_wires[55]),
    .clk_3_N_in(clk_3_wires[54]),
    .prog_clk_3_S_out(prog_clk_3_wires[55]),
    .prog_clk_3_N_in(prog_clk_3_wires[54]),
    .prog_clk_0_S_out(prog_clk_0_wires[80]),
    .prog_clk_0_W_in(prog_clk_0_wires[79]),
    .Reset_E_in(ResetWires[138]),
    .Reset_W_out(ResetWires[135]),
    .pReset_S_in(pResetWires[265]),
    .Test_en_E_in(Test_enWires[138]),
    .Test_en_W_out(Test_enWires[135]),
    .chany_bottom_in(sb_1__1__15_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__16_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_17_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__17_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__17_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__17_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__17_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__17_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__17_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__17_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__17_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__17_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__17_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__17_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__17_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__17_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__17_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__17_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__17_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__17_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__17_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__17_ccff_tail[0])
  );


  cby_1__1_
  cby_2__7_
  (
    .clk_3_N_out(clk_3_wires[53]),
    .clk_3_S_in(clk_3_wires[52]),
    .prog_clk_3_N_out(prog_clk_3_wires[53]),
    .prog_clk_3_S_in(prog_clk_3_wires[52]),
    .prog_clk_0_S_out(prog_clk_0_wires[83]),
    .prog_clk_0_W_in(prog_clk_0_wires[82]),
    .Reset_E_in(ResetWires[160]),
    .Reset_W_out(ResetWires[157]),
    .pReset_S_in(pResetWires[314]),
    .Test_en_E_in(Test_enWires[160]),
    .Test_en_W_out(Test_enWires[157]),
    .chany_bottom_in(sb_1__1__16_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__17_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_18_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__18_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__18_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__18_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__18_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__18_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__18_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__18_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__18_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__18_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__18_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__18_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__18_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__18_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__18_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__18_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__18_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__18_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__18_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__18_ccff_tail[0])
  );


  cby_1__1_
  cby_2__8_
  (
    .clk_3_N_out(clk_3_wires[57]),
    .clk_3_S_in(clk_3_wires[56]),
    .prog_clk_3_N_out(prog_clk_3_wires[57]),
    .prog_clk_3_S_in(prog_clk_3_wires[56]),
    .prog_clk_0_S_out(prog_clk_0_wires[86]),
    .prog_clk_0_W_in(prog_clk_0_wires[85]),
    .Reset_E_in(ResetWires[182]),
    .Reset_W_out(ResetWires[179]),
    .pReset_S_in(pResetWires[363]),
    .Test_en_E_in(Test_enWires[182]),
    .Test_en_W_out(Test_enWires[179]),
    .chany_bottom_in(sb_1__1__17_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__18_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_19_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__19_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__19_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__19_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__19_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__19_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__19_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__19_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__19_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__19_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__19_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__19_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__19_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__19_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__19_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__19_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__19_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__19_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__19_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__19_ccff_tail[0])
  );


  cby_1__1_
  cby_2__9_
  (
    .clk_3_N_out(clk_3_wires[63]),
    .clk_3_S_in(clk_3_wires[62]),
    .prog_clk_3_N_out(prog_clk_3_wires[63]),
    .prog_clk_3_S_in(prog_clk_3_wires[62]),
    .prog_clk_0_S_out(prog_clk_0_wires[89]),
    .prog_clk_0_W_in(prog_clk_0_wires[88]),
    .Reset_E_in(ResetWires[204]),
    .Reset_W_out(ResetWires[201]),
    .pReset_S_in(pResetWires[412]),
    .Test_en_E_in(Test_enWires[204]),
    .Test_en_W_out(Test_enWires[201]),
    .chany_bottom_in(sb_1__1__18_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__19_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_20_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__20_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__20_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__20_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__20_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__20_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__20_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__20_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__20_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__20_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__20_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__20_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__20_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__20_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__20_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__20_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__20_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__20_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__20_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__20_ccff_tail[0])
  );


  cby_1__1_
  cby_2__10_
  (
    .clk_3_N_out(clk_3_wires[67]),
    .clk_3_S_in(clk_3_wires[66]),
    .prog_clk_3_N_out(prog_clk_3_wires[67]),
    .prog_clk_3_S_in(prog_clk_3_wires[66]),
    .prog_clk_0_S_out(prog_clk_0_wires[92]),
    .prog_clk_0_W_in(prog_clk_0_wires[91]),
    .Reset_E_in(ResetWires[226]),
    .Reset_W_out(ResetWires[223]),
    .pReset_S_in(pResetWires[461]),
    .Test_en_E_in(Test_enWires[226]),
    .Test_en_W_out(Test_enWires[223]),
    .chany_bottom_in(sb_1__1__19_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__20_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_21_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__21_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__21_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__21_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__21_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__21_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__21_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__21_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__21_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__21_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__21_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__21_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__21_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__21_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__21_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__21_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__21_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__21_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__21_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__21_ccff_tail[0])
  );


  cby_1__1_
  cby_2__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[95]),
    .prog_clk_0_W_in(prog_clk_0_wires[94]),
    .Reset_E_in(ResetWires[248]),
    .Reset_W_out(ResetWires[245]),
    .pReset_S_in(pResetWires[510]),
    .Test_en_E_in(Test_enWires[248]),
    .Test_en_W_out(Test_enWires[245]),
    .chany_bottom_in(sb_1__1__20_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__21_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_22_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__22_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__22_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__22_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__22_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__22_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__22_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__22_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__22_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__22_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__22_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__22_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__22_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__22_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__22_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__22_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__22_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__22_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__22_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__22_ccff_tail[0])
  );


  cby_1__1_
  cby_2__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[100]),
    .prog_clk_0_S_out(prog_clk_0_wires[98]),
    .prog_clk_0_W_in(prog_clk_0_wires[97]),
    .Reset_E_in(ResetWires[270]),
    .Reset_W_out(ResetWires[267]),
    .pReset_S_in(pResetWires[559]),
    .Test_en_E_in(Test_enWires[270]),
    .Test_en_W_out(Test_enWires[267]),
    .chany_bottom_in(sb_1__1__21_chany_top_out[0:29]),
    .chany_top_in(sb_1__12__1_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_23_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__23_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__23_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__23_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__23_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__23_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__23_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__23_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__23_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__23_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__23_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__23_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__23_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__23_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__23_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__23_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__23_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__23_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__23_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__23_ccff_tail[0])
  );


  cby_1__1_
  cby_3__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[103]),
    .prog_clk_0_W_in(prog_clk_0_wires[102]),
    .Reset_E_in(ResetWires[30]),
    .Reset_W_out(ResetWires[27]),
    .pReset_S_in(pResetWires[33]),
    .Test_en_E_in(Test_enWires[30]),
    .Test_en_W_out(Test_enWires[27]),
    .chany_bottom_in(sb_1__0__2_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__22_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_24_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__24_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__24_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__24_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__24_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__24_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__24_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__24_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__24_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__24_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__24_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__24_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__24_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__24_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__24_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__24_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__24_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__24_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__24_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__24_ccff_tail[0])
  );


  cby_1__1_
  cby_3__2_
  (
    .clk_2_S_out(clk_2_wires[30]),
    .clk_2_N_in(clk_2_wires[29]),
    .prog_clk_2_S_out(prog_clk_2_wires[30]),
    .prog_clk_2_N_in(prog_clk_2_wires[29]),
    .prog_clk_0_S_out(prog_clk_0_wires[106]),
    .prog_clk_0_W_in(prog_clk_0_wires[105]),
    .Reset_E_in(ResetWires[52]),
    .Reset_W_out(ResetWires[49]),
    .pReset_S_in(pResetWires[73]),
    .Test_en_E_in(Test_enWires[52]),
    .Test_en_W_out(Test_enWires[49]),
    .chany_bottom_in(sb_1__1__22_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__23_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_25_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__25_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__25_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__25_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__25_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__25_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__25_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__25_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__25_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__25_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__25_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__25_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__25_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__25_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__25_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__25_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__25_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__25_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__25_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__25_ccff_tail[0])
  );


  cby_1__1_
  cby_3__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[109]),
    .prog_clk_0_W_in(prog_clk_0_wires[108]),
    .Reset_E_in(ResetWires[74]),
    .Reset_W_out(ResetWires[71]),
    .pReset_S_in(pResetWires[122]),
    .Test_en_E_in(Test_enWires[74]),
    .Test_en_W_out(Test_enWires[71]),
    .chany_bottom_in(sb_1__1__23_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__24_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_26_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__26_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__26_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__26_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__26_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__26_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__26_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__26_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__26_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__26_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__26_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__26_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__26_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__26_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__26_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__26_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__26_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__26_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__26_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__26_ccff_tail[0])
  );


  cby_1__1_
  cby_3__4_
  (
    .clk_2_S_out(clk_2_wires[41]),
    .clk_2_N_in(clk_2_wires[40]),
    .prog_clk_2_S_out(prog_clk_2_wires[41]),
    .prog_clk_2_N_in(prog_clk_2_wires[40]),
    .prog_clk_0_S_out(prog_clk_0_wires[112]),
    .prog_clk_0_W_in(prog_clk_0_wires[111]),
    .Reset_E_in(ResetWires[96]),
    .Reset_W_out(ResetWires[93]),
    .pReset_S_in(pResetWires[171]),
    .Test_en_E_in(Test_enWires[96]),
    .Test_en_W_out(Test_enWires[93]),
    .chany_bottom_in(sb_1__1__24_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__25_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_27_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__27_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__27_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__27_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__27_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__27_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__27_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__27_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__27_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__27_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__27_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__27_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__27_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__27_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__27_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__27_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__27_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__27_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__27_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__27_ccff_tail[0])
  );


  cby_1__1_
  cby_3__5_
  (
    .clk_2_N_out(clk_2_wires[39]),
    .clk_2_S_in(clk_2_wires[38]),
    .prog_clk_2_N_out(prog_clk_2_wires[39]),
    .prog_clk_2_S_in(prog_clk_2_wires[38]),
    .prog_clk_0_S_out(prog_clk_0_wires[115]),
    .prog_clk_0_W_in(prog_clk_0_wires[114]),
    .Reset_E_in(ResetWires[118]),
    .Reset_W_out(ResetWires[115]),
    .pReset_S_in(pResetWires[220]),
    .Test_en_E_in(Test_enWires[118]),
    .Test_en_W_out(Test_enWires[115]),
    .chany_bottom_in(sb_1__1__25_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__26_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_28_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__28_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__28_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__28_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__28_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__28_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__28_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__28_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__28_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__28_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__28_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__28_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__28_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__28_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__28_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__28_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__28_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__28_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__28_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__28_ccff_tail[0])
  );


  cby_1__1_
  cby_3__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[118]),
    .prog_clk_0_W_in(prog_clk_0_wires[117]),
    .Reset_E_in(ResetWires[140]),
    .Reset_W_out(ResetWires[137]),
    .pReset_S_in(pResetWires[269]),
    .Test_en_E_in(Test_enWires[140]),
    .Test_en_W_out(Test_enWires[137]),
    .chany_bottom_in(sb_1__1__26_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__27_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_29_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__29_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__29_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__29_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__29_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__29_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__29_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__29_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__29_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__29_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__29_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__29_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__29_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__29_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__29_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__29_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__29_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__29_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__29_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__29_ccff_tail[0])
  );


  cby_1__1_
  cby_3__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[121]),
    .prog_clk_0_W_in(prog_clk_0_wires[120]),
    .Reset_E_in(ResetWires[162]),
    .Reset_W_out(ResetWires[159]),
    .pReset_S_in(pResetWires[318]),
    .Test_en_E_in(Test_enWires[162]),
    .Test_en_W_out(Test_enWires[159]),
    .chany_bottom_in(sb_1__1__27_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__28_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_30_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__30_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__30_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__30_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__30_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__30_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__30_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__30_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__30_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__30_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__30_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__30_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__30_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__30_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__30_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__30_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__30_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__30_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__30_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__30_ccff_tail[0])
  );


  cby_1__1_
  cby_3__8_
  (
    .clk_2_S_out(clk_2_wires[54]),
    .clk_2_N_in(clk_2_wires[53]),
    .prog_clk_2_S_out(prog_clk_2_wires[54]),
    .prog_clk_2_N_in(prog_clk_2_wires[53]),
    .prog_clk_0_S_out(prog_clk_0_wires[124]),
    .prog_clk_0_W_in(prog_clk_0_wires[123]),
    .Reset_E_in(ResetWires[184]),
    .Reset_W_out(ResetWires[181]),
    .pReset_S_in(pResetWires[367]),
    .Test_en_E_in(Test_enWires[184]),
    .Test_en_W_out(Test_enWires[181]),
    .chany_bottom_in(sb_1__1__28_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__29_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_31_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__31_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__31_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__31_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__31_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__31_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__31_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__31_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__31_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__31_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__31_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__31_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__31_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__31_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__31_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__31_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__31_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__31_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__31_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__31_ccff_tail[0])
  );


  cby_1__1_
  cby_3__9_
  (
    .clk_2_N_out(clk_2_wires[52]),
    .clk_2_S_in(clk_2_wires[51]),
    .prog_clk_2_N_out(prog_clk_2_wires[52]),
    .prog_clk_2_S_in(prog_clk_2_wires[51]),
    .prog_clk_0_S_out(prog_clk_0_wires[127]),
    .prog_clk_0_W_in(prog_clk_0_wires[126]),
    .Reset_E_in(ResetWires[206]),
    .Reset_W_out(ResetWires[203]),
    .pReset_S_in(pResetWires[416]),
    .Test_en_E_in(Test_enWires[206]),
    .Test_en_W_out(Test_enWires[203]),
    .chany_bottom_in(sb_1__1__29_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__30_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_32_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__32_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__32_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__32_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__32_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__32_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__32_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__32_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__32_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__32_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__32_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__32_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__32_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__32_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__32_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__32_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__32_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__32_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__32_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__32_ccff_tail[0])
  );


  cby_1__1_
  cby_3__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[130]),
    .prog_clk_0_W_in(prog_clk_0_wires[129]),
    .Reset_E_in(ResetWires[228]),
    .Reset_W_out(ResetWires[225]),
    .pReset_S_in(pResetWires[465]),
    .Test_en_E_in(Test_enWires[228]),
    .Test_en_W_out(Test_enWires[225]),
    .chany_bottom_in(sb_1__1__30_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__31_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_33_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__33_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__33_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__33_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__33_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__33_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__33_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__33_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__33_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__33_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__33_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__33_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__33_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__33_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__33_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__33_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__33_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__33_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__33_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__33_ccff_tail[0])
  );


  cby_1__1_
  cby_3__11_
  (
    .clk_2_N_out(clk_2_wires[65]),
    .clk_2_S_in(clk_2_wires[64]),
    .prog_clk_2_N_out(prog_clk_2_wires[65]),
    .prog_clk_2_S_in(prog_clk_2_wires[64]),
    .prog_clk_0_S_out(prog_clk_0_wires[133]),
    .prog_clk_0_W_in(prog_clk_0_wires[132]),
    .Reset_E_in(ResetWires[250]),
    .Reset_W_out(ResetWires[247]),
    .pReset_S_in(pResetWires[514]),
    .Test_en_E_in(Test_enWires[250]),
    .Test_en_W_out(Test_enWires[247]),
    .chany_bottom_in(sb_1__1__31_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__32_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_34_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__34_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__34_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__34_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__34_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__34_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__34_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__34_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__34_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__34_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__34_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__34_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__34_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__34_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__34_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__34_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__34_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__34_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__34_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__34_ccff_tail[0])
  );


  cby_1__1_
  cby_3__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[138]),
    .prog_clk_0_S_out(prog_clk_0_wires[136]),
    .prog_clk_0_W_in(prog_clk_0_wires[135]),
    .Reset_E_in(ResetWires[272]),
    .Reset_W_out(ResetWires[269]),
    .pReset_S_in(pResetWires[563]),
    .Test_en_E_in(Test_enWires[272]),
    .Test_en_W_out(Test_enWires[269]),
    .chany_bottom_in(sb_1__1__32_chany_top_out[0:29]),
    .chany_top_in(sb_1__12__2_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_35_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__35_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__35_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__35_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__35_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__35_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__35_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__35_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__35_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__35_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__35_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__35_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__35_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__35_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__35_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__35_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__35_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__35_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__35_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__35_ccff_tail[0])
  );


  cby_1__1_
  cby_4__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[141]),
    .prog_clk_0_W_in(prog_clk_0_wires[140]),
    .Reset_E_in(ResetWires[32]),
    .Reset_W_out(ResetWires[29]),
    .pReset_S_in(pResetWires[36]),
    .Test_en_E_in(Test_enWires[32]),
    .Test_en_W_out(Test_enWires[29]),
    .chany_bottom_in(sb_1__0__3_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__33_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_36_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__36_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__36_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__36_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__36_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__36_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__36_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__36_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__36_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__36_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__36_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__36_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__36_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__36_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__36_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__36_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__36_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__36_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__36_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__36_ccff_tail[0])
  );


  cby_1__1_
  cby_4__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[144]),
    .prog_clk_0_W_in(prog_clk_0_wires[143]),
    .Reset_E_in(ResetWires[54]),
    .Reset_W_out(ResetWires[51]),
    .pReset_S_in(pResetWires[77]),
    .Test_en_E_in(Test_enWires[54]),
    .Test_en_W_out(Test_enWires[51]),
    .chany_bottom_in(sb_1__1__33_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__34_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_37_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__37_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__37_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__37_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__37_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__37_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__37_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__37_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__37_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__37_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__37_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__37_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__37_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__37_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__37_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__37_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__37_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__37_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__37_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__37_ccff_tail[0])
  );


  cby_1__1_
  cby_4__3_
  (
    .clk_3_S_out(clk_3_wires[25]),
    .clk_3_N_in(clk_3_wires[24]),
    .prog_clk_3_S_out(prog_clk_3_wires[25]),
    .prog_clk_3_N_in(prog_clk_3_wires[24]),
    .prog_clk_0_S_out(prog_clk_0_wires[147]),
    .prog_clk_0_W_in(prog_clk_0_wires[146]),
    .Reset_E_in(ResetWires[76]),
    .Reset_W_out(ResetWires[73]),
    .pReset_S_in(pResetWires[126]),
    .Test_en_E_in(Test_enWires[76]),
    .Test_en_W_out(Test_enWires[73]),
    .chany_bottom_in(sb_1__1__34_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__35_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_38_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__38_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__38_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__38_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__38_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__38_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__38_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__38_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__38_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__38_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__38_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__38_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__38_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__38_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__38_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__38_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__38_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__38_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__38_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__38_ccff_tail[0])
  );


  cby_1__1_
  cby_4__4_
  (
    .clk_3_S_out(clk_3_wires[21]),
    .clk_3_N_in(clk_3_wires[20]),
    .prog_clk_3_S_out(prog_clk_3_wires[21]),
    .prog_clk_3_N_in(prog_clk_3_wires[20]),
    .prog_clk_0_S_out(prog_clk_0_wires[150]),
    .prog_clk_0_W_in(prog_clk_0_wires[149]),
    .Reset_E_in(ResetWires[98]),
    .Reset_W_out(ResetWires[95]),
    .pReset_S_in(pResetWires[175]),
    .Test_en_E_in(Test_enWires[98]),
    .Test_en_W_out(Test_enWires[95]),
    .chany_bottom_in(sb_1__1__35_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__36_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_39_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__39_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__39_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__39_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__39_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__39_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__39_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__39_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__39_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__39_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__39_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__39_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__39_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__39_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__39_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__39_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__39_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__39_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__39_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__39_ccff_tail[0])
  );


  cby_1__1_
  cby_4__5_
  (
    .clk_3_S_out(clk_3_wires[15]),
    .clk_3_N_in(clk_3_wires[14]),
    .prog_clk_3_S_out(prog_clk_3_wires[15]),
    .prog_clk_3_N_in(prog_clk_3_wires[14]),
    .prog_clk_0_S_out(prog_clk_0_wires[153]),
    .prog_clk_0_W_in(prog_clk_0_wires[152]),
    .Reset_E_in(ResetWires[120]),
    .Reset_W_out(ResetWires[117]),
    .pReset_S_in(pResetWires[224]),
    .Test_en_E_in(Test_enWires[120]),
    .Test_en_W_out(Test_enWires[117]),
    .chany_bottom_in(sb_1__1__36_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__37_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_40_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__40_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__40_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__40_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__40_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__40_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__40_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__40_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__40_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__40_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__40_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__40_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__40_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__40_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__40_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__40_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__40_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__40_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__40_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__40_ccff_tail[0])
  );


  cby_1__1_
  cby_4__6_
  (
    .clk_3_S_out(clk_3_wires[11]),
    .clk_3_N_in(clk_3_wires[10]),
    .prog_clk_3_S_out(prog_clk_3_wires[11]),
    .prog_clk_3_N_in(prog_clk_3_wires[10]),
    .prog_clk_0_S_out(prog_clk_0_wires[156]),
    .prog_clk_0_W_in(prog_clk_0_wires[155]),
    .Reset_E_in(ResetWires[142]),
    .Reset_W_out(ResetWires[139]),
    .pReset_S_in(pResetWires[273]),
    .Test_en_E_in(Test_enWires[142]),
    .Test_en_W_out(Test_enWires[139]),
    .chany_bottom_in(sb_1__1__37_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__38_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_41_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__41_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__41_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__41_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__41_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__41_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__41_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__41_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__41_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__41_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__41_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__41_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__41_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__41_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__41_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__41_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__41_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__41_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__41_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__41_ccff_tail[0])
  );


  cby_1__1_
  cby_4__7_
  (
    .clk_3_N_out(clk_3_wires[9]),
    .clk_3_S_in(clk_3_wires[8]),
    .prog_clk_3_N_out(prog_clk_3_wires[9]),
    .prog_clk_3_S_in(prog_clk_3_wires[8]),
    .prog_clk_0_S_out(prog_clk_0_wires[159]),
    .prog_clk_0_W_in(prog_clk_0_wires[158]),
    .Reset_E_in(ResetWires[164]),
    .Reset_W_out(ResetWires[161]),
    .pReset_S_in(pResetWires[322]),
    .Test_en_E_in(Test_enWires[164]),
    .Test_en_W_out(Test_enWires[161]),
    .chany_bottom_in(sb_1__1__38_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__39_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_42_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__42_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__42_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__42_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__42_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__42_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__42_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__42_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__42_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__42_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__42_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__42_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__42_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__42_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__42_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__42_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__42_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__42_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__42_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__42_ccff_tail[0])
  );


  cby_1__1_
  cby_4__8_
  (
    .clk_3_N_out(clk_3_wires[13]),
    .clk_3_S_in(clk_3_wires[12]),
    .prog_clk_3_N_out(prog_clk_3_wires[13]),
    .prog_clk_3_S_in(prog_clk_3_wires[12]),
    .prog_clk_0_S_out(prog_clk_0_wires[162]),
    .prog_clk_0_W_in(prog_clk_0_wires[161]),
    .Reset_E_in(ResetWires[186]),
    .Reset_W_out(ResetWires[183]),
    .pReset_S_in(pResetWires[371]),
    .Test_en_E_in(Test_enWires[186]),
    .Test_en_W_out(Test_enWires[183]),
    .chany_bottom_in(sb_1__1__39_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__40_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_43_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__43_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__43_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__43_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__43_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__43_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__43_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__43_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__43_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__43_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__43_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__43_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__43_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__43_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__43_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__43_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__43_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__43_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__43_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__43_ccff_tail[0])
  );


  cby_1__1_
  cby_4__9_
  (
    .clk_3_N_out(clk_3_wires[19]),
    .clk_3_S_in(clk_3_wires[18]),
    .prog_clk_3_N_out(prog_clk_3_wires[19]),
    .prog_clk_3_S_in(prog_clk_3_wires[18]),
    .prog_clk_0_S_out(prog_clk_0_wires[165]),
    .prog_clk_0_W_in(prog_clk_0_wires[164]),
    .Reset_E_in(ResetWires[208]),
    .Reset_W_out(ResetWires[205]),
    .pReset_S_in(pResetWires[420]),
    .Test_en_E_in(Test_enWires[208]),
    .Test_en_W_out(Test_enWires[205]),
    .chany_bottom_in(sb_1__1__40_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__41_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_44_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__44_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__44_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__44_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__44_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__44_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__44_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__44_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__44_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__44_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__44_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__44_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__44_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__44_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__44_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__44_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__44_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__44_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__44_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__44_ccff_tail[0])
  );


  cby_1__1_
  cby_4__10_
  (
    .clk_3_N_out(clk_3_wires[23]),
    .clk_3_S_in(clk_3_wires[22]),
    .prog_clk_3_N_out(prog_clk_3_wires[23]),
    .prog_clk_3_S_in(prog_clk_3_wires[22]),
    .prog_clk_0_S_out(prog_clk_0_wires[168]),
    .prog_clk_0_W_in(prog_clk_0_wires[167]),
    .Reset_E_in(ResetWires[230]),
    .Reset_W_out(ResetWires[227]),
    .pReset_S_in(pResetWires[469]),
    .Test_en_E_in(Test_enWires[230]),
    .Test_en_W_out(Test_enWires[227]),
    .chany_bottom_in(sb_1__1__41_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__42_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_45_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__45_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__45_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__45_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__45_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__45_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__45_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__45_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__45_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__45_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__45_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__45_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__45_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__45_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__45_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__45_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__45_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__45_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__45_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__45_ccff_tail[0])
  );


  cby_1__1_
  cby_4__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[171]),
    .prog_clk_0_W_in(prog_clk_0_wires[170]),
    .Reset_E_in(ResetWires[252]),
    .Reset_W_out(ResetWires[249]),
    .pReset_S_in(pResetWires[518]),
    .Test_en_E_in(Test_enWires[252]),
    .Test_en_W_out(Test_enWires[249]),
    .chany_bottom_in(sb_1__1__42_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__43_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_46_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__46_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__46_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__46_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__46_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__46_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__46_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__46_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__46_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__46_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__46_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__46_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__46_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__46_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__46_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__46_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__46_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__46_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__46_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__46_ccff_tail[0])
  );


  cby_1__1_
  cby_4__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[176]),
    .prog_clk_0_S_out(prog_clk_0_wires[174]),
    .prog_clk_0_W_in(prog_clk_0_wires[173]),
    .Reset_E_in(ResetWires[274]),
    .Reset_W_out(ResetWires[271]),
    .pReset_S_in(pResetWires[567]),
    .Test_en_E_in(Test_enWires[274]),
    .Test_en_W_out(Test_enWires[271]),
    .chany_bottom_in(sb_1__1__43_chany_top_out[0:29]),
    .chany_top_in(sb_1__12__3_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_47_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__47_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__47_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__47_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__47_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__47_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__47_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__47_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__47_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__47_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__47_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__47_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__47_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__47_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__47_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__47_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__47_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__47_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__47_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__47_ccff_tail[0])
  );


  cby_1__1_
  cby_5__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[179]),
    .prog_clk_0_W_in(prog_clk_0_wires[178]),
    .Reset_E_in(ResetWires[34]),
    .Reset_W_out(ResetWires[31]),
    .pReset_S_in(pResetWires[39]),
    .Test_en_E_in(Test_enWires[34]),
    .Test_en_W_out(Test_enWires[31]),
    .chany_bottom_in(sb_1__0__4_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__44_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_48_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__48_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__48_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__48_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__48_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__48_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__48_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__48_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__48_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__48_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__48_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__48_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__48_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__48_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__48_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__48_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__48_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__48_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__48_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__48_ccff_tail[0])
  );


  cby_1__1_
  cby_5__2_
  (
    .clk_2_S_out(clk_2_wires[32]),
    .clk_2_N_in(clk_2_wires[31]),
    .prog_clk_2_S_out(prog_clk_2_wires[32]),
    .prog_clk_2_N_in(prog_clk_2_wires[31]),
    .prog_clk_0_S_out(prog_clk_0_wires[182]),
    .prog_clk_0_W_in(prog_clk_0_wires[181]),
    .Reset_E_in(ResetWires[56]),
    .Reset_W_out(ResetWires[53]),
    .pReset_S_in(pResetWires[81]),
    .Test_en_E_in(Test_enWires[56]),
    .Test_en_W_out(Test_enWires[53]),
    .chany_bottom_in(sb_1__1__44_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__45_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_49_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__49_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__49_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__49_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__49_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__49_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__49_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__49_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__49_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__49_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__49_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__49_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__49_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__49_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__49_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__49_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__49_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__49_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__49_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__49_ccff_tail[0])
  );


  cby_1__1_
  cby_5__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[185]),
    .prog_clk_0_W_in(prog_clk_0_wires[184]),
    .Reset_E_in(ResetWires[78]),
    .Reset_W_out(ResetWires[75]),
    .pReset_S_in(pResetWires[130]),
    .Test_en_E_in(Test_enWires[78]),
    .Test_en_W_out(Test_enWires[75]),
    .chany_bottom_in(sb_1__1__45_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__46_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_50_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__50_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__50_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__50_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__50_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__50_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__50_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__50_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__50_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__50_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__50_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__50_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__50_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__50_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__50_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__50_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__50_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__50_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__50_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__50_ccff_tail[0])
  );


  cby_1__1_
  cby_5__4_
  (
    .clk_2_S_out(clk_2_wires[45]),
    .clk_2_N_in(clk_2_wires[44]),
    .prog_clk_2_S_out(prog_clk_2_wires[45]),
    .prog_clk_2_N_in(prog_clk_2_wires[44]),
    .prog_clk_0_S_out(prog_clk_0_wires[188]),
    .prog_clk_0_W_in(prog_clk_0_wires[187]),
    .Reset_E_in(ResetWires[100]),
    .Reset_W_out(ResetWires[97]),
    .pReset_S_in(pResetWires[179]),
    .Test_en_E_in(Test_enWires[100]),
    .Test_en_W_out(Test_enWires[97]),
    .chany_bottom_in(sb_1__1__46_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__47_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_51_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__51_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__51_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__51_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__51_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__51_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__51_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__51_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__51_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__51_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__51_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__51_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__51_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__51_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__51_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__51_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__51_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__51_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__51_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__51_ccff_tail[0])
  );


  cby_1__1_
  cby_5__5_
  (
    .clk_2_N_out(clk_2_wires[43]),
    .clk_2_S_in(clk_2_wires[42]),
    .prog_clk_2_N_out(prog_clk_2_wires[43]),
    .prog_clk_2_S_in(prog_clk_2_wires[42]),
    .prog_clk_0_S_out(prog_clk_0_wires[191]),
    .prog_clk_0_W_in(prog_clk_0_wires[190]),
    .Reset_E_in(ResetWires[122]),
    .Reset_W_out(ResetWires[119]),
    .pReset_S_in(pResetWires[228]),
    .Test_en_E_in(Test_enWires[122]),
    .Test_en_W_out(Test_enWires[119]),
    .chany_bottom_in(sb_1__1__47_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__48_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_52_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__52_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__52_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__52_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__52_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__52_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__52_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__52_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__52_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__52_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__52_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__52_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__52_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__52_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__52_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__52_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__52_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__52_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__52_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__52_ccff_tail[0])
  );


  cby_1__1_
  cby_5__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[194]),
    .prog_clk_0_W_in(prog_clk_0_wires[193]),
    .Reset_E_in(ResetWires[144]),
    .Reset_W_out(ResetWires[141]),
    .pReset_S_in(pResetWires[277]),
    .Test_en_E_in(Test_enWires[144]),
    .Test_en_W_out(Test_enWires[141]),
    .chany_bottom_in(sb_1__1__48_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__49_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_53_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__53_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__53_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__53_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__53_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__53_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__53_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__53_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__53_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__53_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__53_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__53_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__53_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__53_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__53_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__53_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__53_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__53_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__53_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__53_ccff_tail[0])
  );


  cby_1__1_
  cby_5__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[197]),
    .prog_clk_0_W_in(prog_clk_0_wires[196]),
    .Reset_E_in(ResetWires[166]),
    .Reset_W_out(ResetWires[163]),
    .pReset_S_in(pResetWires[326]),
    .Test_en_E_in(Test_enWires[166]),
    .Test_en_W_out(Test_enWires[163]),
    .chany_bottom_in(sb_1__1__49_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__50_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_54_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__54_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__54_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__54_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__54_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__54_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__54_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__54_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__54_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__54_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__54_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__54_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__54_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__54_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__54_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__54_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__54_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__54_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__54_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__54_ccff_tail[0])
  );


  cby_1__1_
  cby_5__8_
  (
    .clk_2_S_out(clk_2_wires[58]),
    .clk_2_N_in(clk_2_wires[57]),
    .prog_clk_2_S_out(prog_clk_2_wires[58]),
    .prog_clk_2_N_in(prog_clk_2_wires[57]),
    .prog_clk_0_S_out(prog_clk_0_wires[200]),
    .prog_clk_0_W_in(prog_clk_0_wires[199]),
    .Reset_E_in(ResetWires[188]),
    .Reset_W_out(ResetWires[185]),
    .pReset_S_in(pResetWires[375]),
    .Test_en_E_in(Test_enWires[188]),
    .Test_en_W_out(Test_enWires[185]),
    .chany_bottom_in(sb_1__1__50_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__51_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_55_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__55_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__55_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__55_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__55_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__55_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__55_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__55_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__55_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__55_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__55_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__55_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__55_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__55_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__55_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__55_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__55_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__55_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__55_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__55_ccff_tail[0])
  );


  cby_1__1_
  cby_5__9_
  (
    .clk_2_N_out(clk_2_wires[56]),
    .clk_2_S_in(clk_2_wires[55]),
    .prog_clk_2_N_out(prog_clk_2_wires[56]),
    .prog_clk_2_S_in(prog_clk_2_wires[55]),
    .prog_clk_0_S_out(prog_clk_0_wires[203]),
    .prog_clk_0_W_in(prog_clk_0_wires[202]),
    .Reset_E_in(ResetWires[210]),
    .Reset_W_out(ResetWires[207]),
    .pReset_S_in(pResetWires[424]),
    .Test_en_E_in(Test_enWires[210]),
    .Test_en_W_out(Test_enWires[207]),
    .chany_bottom_in(sb_1__1__51_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__52_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_56_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__56_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__56_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__56_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__56_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__56_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__56_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__56_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__56_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__56_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__56_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__56_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__56_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__56_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__56_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__56_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__56_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__56_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__56_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__56_ccff_tail[0])
  );


  cby_1__1_
  cby_5__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[206]),
    .prog_clk_0_W_in(prog_clk_0_wires[205]),
    .Reset_E_in(ResetWires[232]),
    .Reset_W_out(ResetWires[229]),
    .pReset_S_in(pResetWires[473]),
    .Test_en_E_in(Test_enWires[232]),
    .Test_en_W_out(Test_enWires[229]),
    .chany_bottom_in(sb_1__1__52_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__53_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_57_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__57_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__57_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__57_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__57_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__57_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__57_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__57_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__57_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__57_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__57_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__57_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__57_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__57_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__57_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__57_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__57_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__57_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__57_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__57_ccff_tail[0])
  );


  cby_1__1_
  cby_5__11_
  (
    .clk_2_N_out(clk_2_wires[67]),
    .clk_2_S_in(clk_2_wires[66]),
    .prog_clk_2_N_out(prog_clk_2_wires[67]),
    .prog_clk_2_S_in(prog_clk_2_wires[66]),
    .prog_clk_0_S_out(prog_clk_0_wires[209]),
    .prog_clk_0_W_in(prog_clk_0_wires[208]),
    .Reset_E_in(ResetWires[254]),
    .Reset_W_out(ResetWires[251]),
    .pReset_S_in(pResetWires[522]),
    .Test_en_E_in(Test_enWires[254]),
    .Test_en_W_out(Test_enWires[251]),
    .chany_bottom_in(sb_1__1__53_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__54_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_58_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__58_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__58_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__58_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__58_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__58_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__58_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__58_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__58_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__58_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__58_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__58_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__58_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__58_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__58_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__58_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__58_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__58_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__58_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__58_ccff_tail[0])
  );


  cby_1__1_
  cby_5__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[214]),
    .prog_clk_0_S_out(prog_clk_0_wires[212]),
    .prog_clk_0_W_in(prog_clk_0_wires[211]),
    .Reset_E_in(ResetWires[276]),
    .Reset_W_out(ResetWires[273]),
    .pReset_S_in(pResetWires[571]),
    .Test_en_E_in(Test_enWires[276]),
    .Test_en_W_out(Test_enWires[273]),
    .chany_bottom_in(sb_1__1__54_chany_top_out[0:29]),
    .chany_top_in(sb_1__12__4_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_59_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__59_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__59_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__59_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__59_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__59_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__59_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__59_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__59_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__59_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__59_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__59_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__59_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__59_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__59_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__59_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__59_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__59_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__59_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__59_ccff_tail[0])
  );


  cby_1__1_
  cby_6__1_
  (
    .clk_3_S_in(clk_3_wires[90]),
    .clk_3_N_out(clk_3_wires[89]),
    .prog_clk_3_S_in(prog_clk_3_wires[90]),
    .prog_clk_3_N_out(prog_clk_3_wires[89]),
    .prog_clk_0_S_out(prog_clk_0_wires[217]),
    .prog_clk_0_W_in(prog_clk_0_wires[216]),
    .Reset_E_out(ResetWires[35]),
    .Reset_W_out(ResetWires[33]),
    .Reset_N_out(ResetWires[2]),
    .Reset_S_in(ResetWires[1]),
    .pReset_N_out(pResetWires[2]),
    .pReset_S_in(pResetWires[42]),
    .Test_en_E_out(Test_enWires[35]),
    .Test_en_W_out(Test_enWires[33]),
    .Test_en_N_out(Test_enWires[2]),
    .Test_en_S_in(Test_enWires[1]),
    .chany_bottom_in(sb_1__0__5_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__55_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_60_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__60_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__60_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__60_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__60_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__60_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__60_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__60_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__60_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__60_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__60_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__60_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__60_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__60_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__60_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__60_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__60_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__60_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__60_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__60_ccff_tail[0])
  );


  cby_1__1_
  cby_6__2_
  (
    .clk_3_S_in(clk_3_wires[92]),
    .clk_3_N_out(clk_3_wires[91]),
    .prog_clk_3_S_in(prog_clk_3_wires[92]),
    .prog_clk_3_N_out(prog_clk_3_wires[91]),
    .prog_clk_0_S_out(prog_clk_0_wires[220]),
    .prog_clk_0_W_in(prog_clk_0_wires[219]),
    .Reset_E_out(ResetWires[57]),
    .Reset_W_out(ResetWires[55]),
    .Reset_N_out(ResetWires[4]),
    .Reset_S_in(ResetWires[3]),
    .pReset_N_out(pResetWires[4]),
    .pReset_S_in(pResetWires[85]),
    .Test_en_E_out(Test_enWires[57]),
    .Test_en_W_out(Test_enWires[55]),
    .Test_en_N_out(Test_enWires[4]),
    .Test_en_S_in(Test_enWires[3]),
    .chany_bottom_in(sb_1__1__55_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__56_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_61_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__61_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__61_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__61_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__61_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__61_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__61_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__61_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__61_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__61_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__61_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__61_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__61_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__61_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__61_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__61_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__61_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__61_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__61_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__61_ccff_tail[0])
  );


  cby_1__1_
  cby_6__3_
  (
    .clk_3_S_in(clk_3_wires[94]),
    .clk_3_N_out(clk_3_wires[93]),
    .prog_clk_3_S_in(prog_clk_3_wires[94]),
    .prog_clk_3_N_out(prog_clk_3_wires[93]),
    .prog_clk_0_S_out(prog_clk_0_wires[223]),
    .prog_clk_0_W_in(prog_clk_0_wires[222]),
    .Reset_E_out(ResetWires[79]),
    .Reset_W_out(ResetWires[77]),
    .Reset_N_out(ResetWires[6]),
    .Reset_S_in(ResetWires[5]),
    .pReset_N_out(pResetWires[6]),
    .pReset_S_in(pResetWires[134]),
    .Test_en_E_out(Test_enWires[79]),
    .Test_en_W_out(Test_enWires[77]),
    .Test_en_N_out(Test_enWires[6]),
    .Test_en_S_in(Test_enWires[5]),
    .chany_bottom_in(sb_1__1__56_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__57_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_62_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__62_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__62_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__62_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__62_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__62_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__62_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__62_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__62_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__62_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__62_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__62_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__62_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__62_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__62_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__62_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__62_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__62_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__62_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__62_ccff_tail[0])
  );


  cby_1__1_
  cby_6__4_
  (
    .clk_3_S_in(clk_3_wires[96]),
    .clk_3_N_out(clk_3_wires[95]),
    .prog_clk_3_S_in(prog_clk_3_wires[96]),
    .prog_clk_3_N_out(prog_clk_3_wires[95]),
    .prog_clk_0_S_out(prog_clk_0_wires[226]),
    .prog_clk_0_W_in(prog_clk_0_wires[225]),
    .Reset_E_out(ResetWires[101]),
    .Reset_W_out(ResetWires[99]),
    .Reset_N_out(ResetWires[8]),
    .Reset_S_in(ResetWires[7]),
    .pReset_N_out(pResetWires[8]),
    .pReset_S_in(pResetWires[183]),
    .Test_en_E_out(Test_enWires[101]),
    .Test_en_W_out(Test_enWires[99]),
    .Test_en_N_out(Test_enWires[8]),
    .Test_en_S_in(Test_enWires[7]),
    .chany_bottom_in(sb_1__1__57_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__58_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_63_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__63_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__63_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__63_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__63_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__63_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__63_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__63_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__63_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__63_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__63_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__63_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__63_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__63_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__63_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__63_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__63_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__63_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__63_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__63_ccff_tail[0])
  );


  cby_1__1_
  cby_6__5_
  (
    .clk_3_S_in(clk_3_wires[98]),
    .clk_3_N_out(clk_3_wires[97]),
    .prog_clk_3_S_in(prog_clk_3_wires[98]),
    .prog_clk_3_N_out(prog_clk_3_wires[97]),
    .prog_clk_0_S_out(prog_clk_0_wires[229]),
    .prog_clk_0_W_in(prog_clk_0_wires[228]),
    .Reset_E_out(ResetWires[123]),
    .Reset_W_out(ResetWires[121]),
    .Reset_N_out(ResetWires[10]),
    .Reset_S_in(ResetWires[9]),
    .pReset_N_out(pResetWires[10]),
    .pReset_S_in(pResetWires[232]),
    .Test_en_E_out(Test_enWires[123]),
    .Test_en_W_out(Test_enWires[121]),
    .Test_en_N_out(Test_enWires[10]),
    .Test_en_S_in(Test_enWires[9]),
    .chany_bottom_in(sb_1__1__58_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__59_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_64_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__64_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__64_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__64_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__64_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__64_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__64_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__64_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__64_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__64_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__64_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__64_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__64_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__64_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__64_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__64_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__64_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__64_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__64_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__64_ccff_tail[0])
  );


  cby_1__1_
  cby_6__6_
  (
    .clk_3_S_in(clk_3_wires[100]),
    .clk_3_N_out(clk_3_wires[99]),
    .prog_clk_3_S_in(prog_clk_3_wires[100]),
    .prog_clk_3_N_out(prog_clk_3_wires[99]),
    .prog_clk_0_S_out(prog_clk_0_wires[232]),
    .prog_clk_0_W_in(prog_clk_0_wires[231]),
    .Reset_E_out(ResetWires[145]),
    .Reset_W_out(ResetWires[143]),
    .Reset_N_out(ResetWires[12]),
    .Reset_S_in(ResetWires[11]),
    .pReset_N_out(pResetWires[12]),
    .pReset_S_in(pResetWires[281]),
    .Test_en_E_out(Test_enWires[145]),
    .Test_en_W_out(Test_enWires[143]),
    .Test_en_N_out(Test_enWires[12]),
    .Test_en_S_in(Test_enWires[11]),
    .chany_bottom_in(sb_1__1__59_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__60_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_65_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__65_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__65_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__65_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__65_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__65_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__65_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__65_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__65_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__65_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__65_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__65_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__65_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__65_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__65_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__65_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__65_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__65_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__65_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__65_ccff_tail[0])
  );


  cby_1__1_
  cby_6__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[235]),
    .prog_clk_0_W_in(prog_clk_0_wires[234]),
    .Reset_E_out(ResetWires[167]),
    .Reset_W_out(ResetWires[165]),
    .Reset_N_out(ResetWires[14]),
    .Reset_S_in(ResetWires[13]),
    .pReset_N_out(pResetWires[14]),
    .pReset_S_in(pResetWires[330]),
    .Test_en_E_out(Test_enWires[167]),
    .Test_en_W_out(Test_enWires[165]),
    .Test_en_N_out(Test_enWires[14]),
    .Test_en_S_in(Test_enWires[13]),
    .chany_bottom_in(sb_1__1__60_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__61_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_66_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__66_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__66_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__66_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__66_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__66_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__66_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__66_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__66_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__66_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__66_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__66_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__66_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__66_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__66_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__66_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__66_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__66_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__66_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__66_ccff_tail[0])
  );


  cby_1__1_
  cby_6__8_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[238]),
    .prog_clk_0_W_in(prog_clk_0_wires[237]),
    .Reset_E_out(ResetWires[189]),
    .Reset_W_out(ResetWires[187]),
    .Reset_N_out(ResetWires[16]),
    .Reset_S_in(ResetWires[15]),
    .pReset_N_out(pResetWires[16]),
    .pReset_S_in(pResetWires[379]),
    .Test_en_E_out(Test_enWires[189]),
    .Test_en_W_out(Test_enWires[187]),
    .Test_en_N_out(Test_enWires[16]),
    .Test_en_S_in(Test_enWires[15]),
    .chany_bottom_in(sb_1__1__61_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__62_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_67_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__67_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__67_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__67_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__67_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__67_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__67_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__67_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__67_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__67_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__67_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__67_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__67_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__67_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__67_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__67_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__67_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__67_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__67_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__67_ccff_tail[0])
  );


  cby_1__1_
  cby_6__9_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[241]),
    .prog_clk_0_W_in(prog_clk_0_wires[240]),
    .Reset_E_out(ResetWires[211]),
    .Reset_W_out(ResetWires[209]),
    .Reset_N_out(ResetWires[18]),
    .Reset_S_in(ResetWires[17]),
    .pReset_N_out(pResetWires[18]),
    .pReset_S_in(pResetWires[428]),
    .Test_en_E_out(Test_enWires[211]),
    .Test_en_W_out(Test_enWires[209]),
    .Test_en_N_out(Test_enWires[18]),
    .Test_en_S_in(Test_enWires[17]),
    .chany_bottom_in(sb_1__1__62_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__63_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_68_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__68_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__68_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__68_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__68_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__68_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__68_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__68_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__68_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__68_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__68_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__68_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__68_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__68_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__68_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__68_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__68_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__68_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__68_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__68_ccff_tail[0])
  );


  cby_1__1_
  cby_6__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[244]),
    .prog_clk_0_W_in(prog_clk_0_wires[243]),
    .Reset_E_out(ResetWires[233]),
    .Reset_W_out(ResetWires[231]),
    .Reset_N_out(ResetWires[20]),
    .Reset_S_in(ResetWires[19]),
    .pReset_N_out(pResetWires[20]),
    .pReset_S_in(pResetWires[477]),
    .Test_en_E_out(Test_enWires[233]),
    .Test_en_W_out(Test_enWires[231]),
    .Test_en_N_out(Test_enWires[20]),
    .Test_en_S_in(Test_enWires[19]),
    .chany_bottom_in(sb_1__1__63_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__64_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_69_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__69_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__69_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__69_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__69_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__69_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__69_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__69_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__69_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__69_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__69_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__69_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__69_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__69_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__69_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__69_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__69_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__69_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__69_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__69_ccff_tail[0])
  );


  cby_1__1_
  cby_6__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[247]),
    .prog_clk_0_W_in(prog_clk_0_wires[246]),
    .Reset_E_out(ResetWires[255]),
    .Reset_W_out(ResetWires[253]),
    .Reset_N_out(ResetWires[22]),
    .Reset_S_in(ResetWires[21]),
    .pReset_N_out(pResetWires[22]),
    .pReset_S_in(pResetWires[526]),
    .Test_en_E_out(Test_enWires[255]),
    .Test_en_W_out(Test_enWires[253]),
    .Test_en_N_out(Test_enWires[22]),
    .Test_en_S_in(Test_enWires[21]),
    .chany_bottom_in(sb_1__1__64_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__65_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_70_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__70_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__70_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__70_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__70_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__70_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__70_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__70_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__70_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__70_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__70_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__70_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__70_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__70_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__70_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__70_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__70_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__70_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__70_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__70_ccff_tail[0])
  );


  cby_1__1_
  cby_6__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[252]),
    .prog_clk_0_S_out(prog_clk_0_wires[250]),
    .prog_clk_0_W_in(prog_clk_0_wires[249]),
    .Reset_E_out(ResetWires[277]),
    .Reset_W_out(ResetWires[275]),
    .Reset_S_in(ResetWires[23]),
    .pReset_N_out(pResetWires[24]),
    .pReset_S_in(pResetWires[575]),
    .Test_en_E_out(Test_enWires[277]),
    .Test_en_W_out(Test_enWires[275]),
    .Test_en_S_in(Test_enWires[23]),
    .chany_bottom_in(sb_1__1__65_chany_top_out[0:29]),
    .chany_top_in(sb_1__12__5_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_71_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__71_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__71_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__71_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__71_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__71_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__71_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__71_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__71_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__71_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__71_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__71_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__71_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__71_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__71_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__71_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__71_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__71_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__71_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__71_ccff_tail[0])
  );


  cby_1__1_
  cby_7__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[255]),
    .prog_clk_0_W_in(prog_clk_0_wires[254]),
    .Reset_E_out(ResetWires[37]),
    .Reset_W_in(ResetWires[36]),
    .pReset_S_in(pResetWires[45]),
    .Test_en_E_out(Test_enWires[37]),
    .Test_en_W_in(Test_enWires[36]),
    .chany_bottom_in(sb_1__0__6_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__66_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_72_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__72_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__72_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__72_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__72_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__72_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__72_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__72_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__72_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__72_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__72_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__72_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__72_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__72_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__72_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__72_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__72_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__72_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__72_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__72_ccff_tail[0])
  );


  cby_1__1_
  cby_7__2_
  (
    .clk_2_S_out(clk_2_wires[74]),
    .clk_2_N_in(clk_2_wires[73]),
    .prog_clk_2_S_out(prog_clk_2_wires[74]),
    .prog_clk_2_N_in(prog_clk_2_wires[73]),
    .prog_clk_0_S_out(prog_clk_0_wires[258]),
    .prog_clk_0_W_in(prog_clk_0_wires[257]),
    .Reset_E_out(ResetWires[59]),
    .Reset_W_in(ResetWires[58]),
    .pReset_S_in(pResetWires[89]),
    .Test_en_E_out(Test_enWires[59]),
    .Test_en_W_in(Test_enWires[58]),
    .chany_bottom_in(sb_1__1__66_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__67_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_73_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__73_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__73_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__73_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__73_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__73_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__73_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__73_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__73_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__73_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__73_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__73_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__73_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__73_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__73_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__73_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__73_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__73_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__73_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__73_ccff_tail[0])
  );


  cby_1__1_
  cby_7__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[261]),
    .prog_clk_0_W_in(prog_clk_0_wires[260]),
    .Reset_E_out(ResetWires[81]),
    .Reset_W_in(ResetWires[80]),
    .pReset_S_in(pResetWires[138]),
    .Test_en_E_out(Test_enWires[81]),
    .Test_en_W_in(Test_enWires[80]),
    .chany_bottom_in(sb_1__1__67_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__68_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_74_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__74_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__74_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__74_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__74_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__74_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__74_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__74_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__74_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__74_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__74_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__74_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__74_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__74_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__74_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__74_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__74_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__74_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__74_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__74_ccff_tail[0])
  );


  cby_1__1_
  cby_7__4_
  (
    .clk_2_S_out(clk_2_wires[85]),
    .clk_2_N_in(clk_2_wires[84]),
    .prog_clk_2_S_out(prog_clk_2_wires[85]),
    .prog_clk_2_N_in(prog_clk_2_wires[84]),
    .prog_clk_0_S_out(prog_clk_0_wires[264]),
    .prog_clk_0_W_in(prog_clk_0_wires[263]),
    .Reset_E_out(ResetWires[103]),
    .Reset_W_in(ResetWires[102]),
    .pReset_S_in(pResetWires[187]),
    .Test_en_E_out(Test_enWires[103]),
    .Test_en_W_in(Test_enWires[102]),
    .chany_bottom_in(sb_1__1__68_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__69_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_75_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__75_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__75_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__75_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__75_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__75_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__75_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__75_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__75_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__75_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__75_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__75_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__75_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__75_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__75_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__75_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__75_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__75_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__75_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__75_ccff_tail[0])
  );


  cby_1__1_
  cby_7__5_
  (
    .clk_2_N_out(clk_2_wires[83]),
    .clk_2_S_in(clk_2_wires[82]),
    .prog_clk_2_N_out(prog_clk_2_wires[83]),
    .prog_clk_2_S_in(prog_clk_2_wires[82]),
    .prog_clk_0_S_out(prog_clk_0_wires[267]),
    .prog_clk_0_W_in(prog_clk_0_wires[266]),
    .Reset_E_out(ResetWires[125]),
    .Reset_W_in(ResetWires[124]),
    .pReset_S_in(pResetWires[236]),
    .Test_en_E_out(Test_enWires[125]),
    .Test_en_W_in(Test_enWires[124]),
    .chany_bottom_in(sb_1__1__69_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__70_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_76_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__76_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__76_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__76_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__76_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__76_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__76_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__76_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__76_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__76_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__76_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__76_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__76_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__76_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__76_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__76_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__76_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__76_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__76_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__76_ccff_tail[0])
  );


  cby_1__1_
  cby_7__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[270]),
    .prog_clk_0_W_in(prog_clk_0_wires[269]),
    .Reset_E_out(ResetWires[147]),
    .Reset_W_in(ResetWires[146]),
    .pReset_S_in(pResetWires[285]),
    .Test_en_E_out(Test_enWires[147]),
    .Test_en_W_in(Test_enWires[146]),
    .chany_bottom_in(sb_1__1__70_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__71_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_77_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__77_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__77_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__77_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__77_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__77_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__77_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__77_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__77_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__77_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__77_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__77_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__77_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__77_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__77_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__77_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__77_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__77_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__77_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__77_ccff_tail[0])
  );


  cby_1__1_
  cby_7__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[273]),
    .prog_clk_0_W_in(prog_clk_0_wires[272]),
    .Reset_E_out(ResetWires[169]),
    .Reset_W_in(ResetWires[168]),
    .pReset_S_in(pResetWires[334]),
    .Test_en_E_out(Test_enWires[169]),
    .Test_en_W_in(Test_enWires[168]),
    .chany_bottom_in(sb_1__1__71_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__72_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_78_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__78_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__78_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__78_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__78_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__78_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__78_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__78_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__78_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__78_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__78_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__78_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__78_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__78_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__78_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__78_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__78_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__78_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__78_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__78_ccff_tail[0])
  );


  cby_1__1_
  cby_7__8_
  (
    .clk_2_S_out(clk_2_wires[98]),
    .clk_2_N_in(clk_2_wires[97]),
    .prog_clk_2_S_out(prog_clk_2_wires[98]),
    .prog_clk_2_N_in(prog_clk_2_wires[97]),
    .prog_clk_0_S_out(prog_clk_0_wires[276]),
    .prog_clk_0_W_in(prog_clk_0_wires[275]),
    .Reset_E_out(ResetWires[191]),
    .Reset_W_in(ResetWires[190]),
    .pReset_S_in(pResetWires[383]),
    .Test_en_E_out(Test_enWires[191]),
    .Test_en_W_in(Test_enWires[190]),
    .chany_bottom_in(sb_1__1__72_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__73_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_79_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__79_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__79_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__79_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__79_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__79_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__79_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__79_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__79_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__79_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__79_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__79_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__79_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__79_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__79_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__79_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__79_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__79_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__79_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__79_ccff_tail[0])
  );


  cby_1__1_
  cby_7__9_
  (
    .clk_2_N_out(clk_2_wires[96]),
    .clk_2_S_in(clk_2_wires[95]),
    .prog_clk_2_N_out(prog_clk_2_wires[96]),
    .prog_clk_2_S_in(prog_clk_2_wires[95]),
    .prog_clk_0_S_out(prog_clk_0_wires[279]),
    .prog_clk_0_W_in(prog_clk_0_wires[278]),
    .Reset_E_out(ResetWires[213]),
    .Reset_W_in(ResetWires[212]),
    .pReset_S_in(pResetWires[432]),
    .Test_en_E_out(Test_enWires[213]),
    .Test_en_W_in(Test_enWires[212]),
    .chany_bottom_in(sb_1__1__73_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__74_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_80_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__80_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__80_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__80_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__80_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__80_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__80_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__80_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__80_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__80_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__80_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__80_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__80_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__80_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__80_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__80_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__80_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__80_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__80_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__80_ccff_tail[0])
  );


  cby_1__1_
  cby_7__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[282]),
    .prog_clk_0_W_in(prog_clk_0_wires[281]),
    .Reset_E_out(ResetWires[235]),
    .Reset_W_in(ResetWires[234]),
    .pReset_S_in(pResetWires[481]),
    .Test_en_E_out(Test_enWires[235]),
    .Test_en_W_in(Test_enWires[234]),
    .chany_bottom_in(sb_1__1__74_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__75_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_81_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__81_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__81_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__81_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__81_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__81_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__81_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__81_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__81_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__81_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__81_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__81_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__81_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__81_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__81_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__81_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__81_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__81_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__81_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__81_ccff_tail[0])
  );


  cby_1__1_
  cby_7__11_
  (
    .clk_2_N_out(clk_2_wires[109]),
    .clk_2_S_in(clk_2_wires[108]),
    .prog_clk_2_N_out(prog_clk_2_wires[109]),
    .prog_clk_2_S_in(prog_clk_2_wires[108]),
    .prog_clk_0_S_out(prog_clk_0_wires[285]),
    .prog_clk_0_W_in(prog_clk_0_wires[284]),
    .Reset_E_out(ResetWires[257]),
    .Reset_W_in(ResetWires[256]),
    .pReset_S_in(pResetWires[530]),
    .Test_en_E_out(Test_enWires[257]),
    .Test_en_W_in(Test_enWires[256]),
    .chany_bottom_in(sb_1__1__75_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__76_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_82_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__82_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__82_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__82_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__82_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__82_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__82_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__82_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__82_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__82_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__82_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__82_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__82_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__82_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__82_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__82_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__82_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__82_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__82_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__82_ccff_tail[0])
  );


  cby_1__1_
  cby_7__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[290]),
    .prog_clk_0_S_out(prog_clk_0_wires[288]),
    .prog_clk_0_W_in(prog_clk_0_wires[287]),
    .Reset_E_out(ResetWires[279]),
    .Reset_W_in(ResetWires[278]),
    .pReset_S_in(pResetWires[579]),
    .Test_en_E_out(Test_enWires[279]),
    .Test_en_W_in(Test_enWires[278]),
    .chany_bottom_in(sb_1__1__76_chany_top_out[0:29]),
    .chany_top_in(sb_1__12__6_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_83_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__83_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__83_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__83_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__83_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__83_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__83_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__83_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__83_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__83_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__83_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__83_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__83_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__83_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__83_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__83_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__83_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__83_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__83_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__83_ccff_tail[0])
  );


  cby_1__1_
  cby_8__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[293]),
    .prog_clk_0_W_in(prog_clk_0_wires[292]),
    .Reset_E_out(ResetWires[39]),
    .Reset_W_in(ResetWires[38]),
    .pReset_S_in(pResetWires[48]),
    .Test_en_E_out(Test_enWires[39]),
    .Test_en_W_in(Test_enWires[38]),
    .chany_bottom_in(sb_1__0__7_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__77_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_84_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__84_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__84_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__84_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__84_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__84_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__84_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__84_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__84_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__84_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__84_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__84_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__84_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__84_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__84_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__84_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__84_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__84_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__84_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__84_ccff_tail[0])
  );


  cby_1__1_
  cby_8__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[296]),
    .prog_clk_0_W_in(prog_clk_0_wires[295]),
    .Reset_E_out(ResetWires[61]),
    .Reset_W_in(ResetWires[60]),
    .pReset_S_in(pResetWires[93]),
    .Test_en_E_out(Test_enWires[61]),
    .Test_en_W_in(Test_enWires[60]),
    .chany_bottom_in(sb_1__1__77_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__78_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_85_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__85_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__85_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__85_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__85_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__85_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__85_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__85_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__85_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__85_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__85_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__85_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__85_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__85_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__85_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__85_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__85_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__85_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__85_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__85_ccff_tail[0])
  );


  cby_1__1_
  cby_8__3_
  (
    .clk_3_S_out(clk_3_wires[43]),
    .clk_3_N_in(clk_3_wires[42]),
    .prog_clk_3_S_out(prog_clk_3_wires[43]),
    .prog_clk_3_N_in(prog_clk_3_wires[42]),
    .prog_clk_0_S_out(prog_clk_0_wires[299]),
    .prog_clk_0_W_in(prog_clk_0_wires[298]),
    .Reset_E_out(ResetWires[83]),
    .Reset_W_in(ResetWires[82]),
    .pReset_S_in(pResetWires[142]),
    .Test_en_E_out(Test_enWires[83]),
    .Test_en_W_in(Test_enWires[82]),
    .chany_bottom_in(sb_1__1__78_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__79_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_86_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__86_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__86_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__86_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__86_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__86_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__86_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__86_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__86_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__86_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__86_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__86_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__86_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__86_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__86_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__86_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__86_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__86_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__86_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__86_ccff_tail[0])
  );


  cby_1__1_
  cby_8__4_
  (
    .clk_3_S_out(clk_3_wires[39]),
    .clk_3_N_in(clk_3_wires[38]),
    .prog_clk_3_S_out(prog_clk_3_wires[39]),
    .prog_clk_3_N_in(prog_clk_3_wires[38]),
    .prog_clk_0_S_out(prog_clk_0_wires[302]),
    .prog_clk_0_W_in(prog_clk_0_wires[301]),
    .Reset_E_out(ResetWires[105]),
    .Reset_W_in(ResetWires[104]),
    .pReset_S_in(pResetWires[191]),
    .Test_en_E_out(Test_enWires[105]),
    .Test_en_W_in(Test_enWires[104]),
    .chany_bottom_in(sb_1__1__79_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__80_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_87_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__87_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__87_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__87_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__87_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__87_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__87_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__87_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__87_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__87_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__87_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__87_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__87_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__87_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__87_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__87_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__87_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__87_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__87_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__87_ccff_tail[0])
  );


  cby_1__1_
  cby_8__5_
  (
    .clk_3_S_out(clk_3_wires[33]),
    .clk_3_N_in(clk_3_wires[32]),
    .prog_clk_3_S_out(prog_clk_3_wires[33]),
    .prog_clk_3_N_in(prog_clk_3_wires[32]),
    .prog_clk_0_S_out(prog_clk_0_wires[305]),
    .prog_clk_0_W_in(prog_clk_0_wires[304]),
    .Reset_E_out(ResetWires[127]),
    .Reset_W_in(ResetWires[126]),
    .pReset_S_in(pResetWires[240]),
    .Test_en_E_out(Test_enWires[127]),
    .Test_en_W_in(Test_enWires[126]),
    .chany_bottom_in(sb_1__1__80_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__81_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_88_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__88_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__88_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__88_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__88_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__88_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__88_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__88_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__88_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__88_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__88_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__88_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__88_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__88_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__88_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__88_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__88_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__88_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__88_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__88_ccff_tail[0])
  );


  cby_1__1_
  cby_8__6_
  (
    .clk_3_S_out(clk_3_wires[29]),
    .clk_3_N_in(clk_3_wires[28]),
    .prog_clk_3_S_out(prog_clk_3_wires[29]),
    .prog_clk_3_N_in(prog_clk_3_wires[28]),
    .prog_clk_0_S_out(prog_clk_0_wires[308]),
    .prog_clk_0_W_in(prog_clk_0_wires[307]),
    .Reset_E_out(ResetWires[149]),
    .Reset_W_in(ResetWires[148]),
    .pReset_S_in(pResetWires[289]),
    .Test_en_E_out(Test_enWires[149]),
    .Test_en_W_in(Test_enWires[148]),
    .chany_bottom_in(sb_1__1__81_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__82_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_89_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__89_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__89_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__89_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__89_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__89_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__89_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__89_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__89_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__89_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__89_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__89_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__89_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__89_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__89_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__89_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__89_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__89_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__89_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__89_ccff_tail[0])
  );


  cby_1__1_
  cby_8__7_
  (
    .clk_3_N_out(clk_3_wires[27]),
    .clk_3_S_in(clk_3_wires[26]),
    .prog_clk_3_N_out(prog_clk_3_wires[27]),
    .prog_clk_3_S_in(prog_clk_3_wires[26]),
    .prog_clk_0_S_out(prog_clk_0_wires[311]),
    .prog_clk_0_W_in(prog_clk_0_wires[310]),
    .Reset_E_out(ResetWires[171]),
    .Reset_W_in(ResetWires[170]),
    .pReset_S_in(pResetWires[338]),
    .Test_en_E_out(Test_enWires[171]),
    .Test_en_W_in(Test_enWires[170]),
    .chany_bottom_in(sb_1__1__82_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__83_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_90_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__90_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__90_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__90_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__90_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__90_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__90_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__90_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__90_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__90_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__90_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__90_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__90_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__90_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__90_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__90_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__90_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__90_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__90_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__90_ccff_tail[0])
  );


  cby_1__1_
  cby_8__8_
  (
    .clk_3_N_out(clk_3_wires[31]),
    .clk_3_S_in(clk_3_wires[30]),
    .prog_clk_3_N_out(prog_clk_3_wires[31]),
    .prog_clk_3_S_in(prog_clk_3_wires[30]),
    .prog_clk_0_S_out(prog_clk_0_wires[314]),
    .prog_clk_0_W_in(prog_clk_0_wires[313]),
    .Reset_E_out(ResetWires[193]),
    .Reset_W_in(ResetWires[192]),
    .pReset_S_in(pResetWires[387]),
    .Test_en_E_out(Test_enWires[193]),
    .Test_en_W_in(Test_enWires[192]),
    .chany_bottom_in(sb_1__1__83_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__84_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_91_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__91_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__91_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__91_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__91_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__91_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__91_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__91_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__91_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__91_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__91_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__91_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__91_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__91_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__91_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__91_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__91_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__91_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__91_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__91_ccff_tail[0])
  );


  cby_1__1_
  cby_8__9_
  (
    .clk_3_N_out(clk_3_wires[37]),
    .clk_3_S_in(clk_3_wires[36]),
    .prog_clk_3_N_out(prog_clk_3_wires[37]),
    .prog_clk_3_S_in(prog_clk_3_wires[36]),
    .prog_clk_0_S_out(prog_clk_0_wires[317]),
    .prog_clk_0_W_in(prog_clk_0_wires[316]),
    .Reset_E_out(ResetWires[215]),
    .Reset_W_in(ResetWires[214]),
    .pReset_S_in(pResetWires[436]),
    .Test_en_E_out(Test_enWires[215]),
    .Test_en_W_in(Test_enWires[214]),
    .chany_bottom_in(sb_1__1__84_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__85_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_92_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__92_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__92_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__92_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__92_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__92_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__92_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__92_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__92_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__92_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__92_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__92_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__92_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__92_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__92_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__92_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__92_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__92_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__92_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__92_ccff_tail[0])
  );


  cby_1__1_
  cby_8__10_
  (
    .clk_3_N_out(clk_3_wires[41]),
    .clk_3_S_in(clk_3_wires[40]),
    .prog_clk_3_N_out(prog_clk_3_wires[41]),
    .prog_clk_3_S_in(prog_clk_3_wires[40]),
    .prog_clk_0_S_out(prog_clk_0_wires[320]),
    .prog_clk_0_W_in(prog_clk_0_wires[319]),
    .Reset_E_out(ResetWires[237]),
    .Reset_W_in(ResetWires[236]),
    .pReset_S_in(pResetWires[485]),
    .Test_en_E_out(Test_enWires[237]),
    .Test_en_W_in(Test_enWires[236]),
    .chany_bottom_in(sb_1__1__85_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__86_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_93_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__93_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__93_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__93_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__93_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__93_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__93_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__93_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__93_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__93_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__93_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__93_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__93_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__93_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__93_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__93_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__93_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__93_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__93_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__93_ccff_tail[0])
  );


  cby_1__1_
  cby_8__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[323]),
    .prog_clk_0_W_in(prog_clk_0_wires[322]),
    .Reset_E_out(ResetWires[259]),
    .Reset_W_in(ResetWires[258]),
    .pReset_S_in(pResetWires[534]),
    .Test_en_E_out(Test_enWires[259]),
    .Test_en_W_in(Test_enWires[258]),
    .chany_bottom_in(sb_1__1__86_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__87_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_94_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__94_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__94_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__94_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__94_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__94_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__94_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__94_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__94_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__94_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__94_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__94_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__94_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__94_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__94_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__94_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__94_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__94_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__94_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__94_ccff_tail[0])
  );


  cby_1__1_
  cby_8__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[328]),
    .prog_clk_0_S_out(prog_clk_0_wires[326]),
    .prog_clk_0_W_in(prog_clk_0_wires[325]),
    .Reset_E_out(ResetWires[281]),
    .Reset_W_in(ResetWires[280]),
    .pReset_S_in(pResetWires[583]),
    .Test_en_E_out(Test_enWires[281]),
    .Test_en_W_in(Test_enWires[280]),
    .chany_bottom_in(sb_1__1__87_chany_top_out[0:29]),
    .chany_top_in(sb_1__12__7_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_95_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__95_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__95_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__95_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__95_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__95_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__95_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__95_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__95_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__95_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__95_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__95_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__95_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__95_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__95_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__95_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__95_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__95_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__95_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__95_ccff_tail[0])
  );


  cby_1__1_
  cby_9__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[331]),
    .prog_clk_0_W_in(prog_clk_0_wires[330]),
    .Reset_E_out(ResetWires[41]),
    .Reset_W_in(ResetWires[40]),
    .pReset_S_in(pResetWires[51]),
    .Test_en_E_out(Test_enWires[41]),
    .Test_en_W_in(Test_enWires[40]),
    .chany_bottom_in(sb_1__0__8_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__88_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_96_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__96_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__96_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__96_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__96_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__96_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__96_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__96_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__96_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__96_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__96_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__96_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__96_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__96_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__96_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__96_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__96_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__96_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__96_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__96_ccff_tail[0])
  );


  cby_1__1_
  cby_9__2_
  (
    .clk_2_S_out(clk_2_wires[76]),
    .clk_2_N_in(clk_2_wires[75]),
    .prog_clk_2_S_out(prog_clk_2_wires[76]),
    .prog_clk_2_N_in(prog_clk_2_wires[75]),
    .prog_clk_0_S_out(prog_clk_0_wires[334]),
    .prog_clk_0_W_in(prog_clk_0_wires[333]),
    .Reset_E_out(ResetWires[63]),
    .Reset_W_in(ResetWires[62]),
    .pReset_S_in(pResetWires[97]),
    .Test_en_E_out(Test_enWires[63]),
    .Test_en_W_in(Test_enWires[62]),
    .chany_bottom_in(sb_1__1__88_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__89_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_97_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__97_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__97_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__97_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__97_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__97_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__97_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__97_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__97_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__97_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__97_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__97_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__97_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__97_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__97_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__97_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__97_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__97_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__97_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__97_ccff_tail[0])
  );


  cby_1__1_
  cby_9__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[337]),
    .prog_clk_0_W_in(prog_clk_0_wires[336]),
    .Reset_E_out(ResetWires[85]),
    .Reset_W_in(ResetWires[84]),
    .pReset_S_in(pResetWires[146]),
    .Test_en_E_out(Test_enWires[85]),
    .Test_en_W_in(Test_enWires[84]),
    .chany_bottom_in(sb_1__1__89_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__90_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_98_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__98_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__98_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__98_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__98_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__98_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__98_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__98_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__98_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__98_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__98_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__98_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__98_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__98_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__98_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__98_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__98_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__98_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__98_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__98_ccff_tail[0])
  );


  cby_1__1_
  cby_9__4_
  (
    .clk_2_S_out(clk_2_wires[89]),
    .clk_2_N_in(clk_2_wires[88]),
    .prog_clk_2_S_out(prog_clk_2_wires[89]),
    .prog_clk_2_N_in(prog_clk_2_wires[88]),
    .prog_clk_0_S_out(prog_clk_0_wires[340]),
    .prog_clk_0_W_in(prog_clk_0_wires[339]),
    .Reset_E_out(ResetWires[107]),
    .Reset_W_in(ResetWires[106]),
    .pReset_S_in(pResetWires[195]),
    .Test_en_E_out(Test_enWires[107]),
    .Test_en_W_in(Test_enWires[106]),
    .chany_bottom_in(sb_1__1__90_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__91_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_99_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__99_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__99_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__99_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__99_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__99_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__99_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__99_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__99_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__99_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__99_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__99_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__99_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__99_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__99_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__99_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__99_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__99_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__99_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__99_ccff_tail[0])
  );


  cby_1__1_
  cby_9__5_
  (
    .clk_2_N_out(clk_2_wires[87]),
    .clk_2_S_in(clk_2_wires[86]),
    .prog_clk_2_N_out(prog_clk_2_wires[87]),
    .prog_clk_2_S_in(prog_clk_2_wires[86]),
    .prog_clk_0_S_out(prog_clk_0_wires[343]),
    .prog_clk_0_W_in(prog_clk_0_wires[342]),
    .Reset_E_out(ResetWires[129]),
    .Reset_W_in(ResetWires[128]),
    .pReset_S_in(pResetWires[244]),
    .Test_en_E_out(Test_enWires[129]),
    .Test_en_W_in(Test_enWires[128]),
    .chany_bottom_in(sb_1__1__91_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__92_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_100_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__100_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__100_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__100_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__100_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__100_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__100_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__100_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__100_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__100_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__100_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__100_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__100_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__100_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__100_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__100_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__100_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__100_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__100_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__100_ccff_tail[0])
  );


  cby_1__1_
  cby_9__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[346]),
    .prog_clk_0_W_in(prog_clk_0_wires[345]),
    .Reset_E_out(ResetWires[151]),
    .Reset_W_in(ResetWires[150]),
    .pReset_S_in(pResetWires[293]),
    .Test_en_E_out(Test_enWires[151]),
    .Test_en_W_in(Test_enWires[150]),
    .chany_bottom_in(sb_1__1__92_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__93_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_101_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__101_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__101_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__101_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__101_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__101_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__101_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__101_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__101_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__101_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__101_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__101_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__101_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__101_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__101_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__101_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__101_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__101_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__101_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__101_ccff_tail[0])
  );


  cby_1__1_
  cby_9__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[349]),
    .prog_clk_0_W_in(prog_clk_0_wires[348]),
    .Reset_E_out(ResetWires[173]),
    .Reset_W_in(ResetWires[172]),
    .pReset_S_in(pResetWires[342]),
    .Test_en_E_out(Test_enWires[173]),
    .Test_en_W_in(Test_enWires[172]),
    .chany_bottom_in(sb_1__1__93_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__94_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_102_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__102_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__102_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__102_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__102_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__102_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__102_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__102_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__102_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__102_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__102_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__102_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__102_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__102_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__102_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__102_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__102_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__102_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__102_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__102_ccff_tail[0])
  );


  cby_1__1_
  cby_9__8_
  (
    .clk_2_S_out(clk_2_wires[102]),
    .clk_2_N_in(clk_2_wires[101]),
    .prog_clk_2_S_out(prog_clk_2_wires[102]),
    .prog_clk_2_N_in(prog_clk_2_wires[101]),
    .prog_clk_0_S_out(prog_clk_0_wires[352]),
    .prog_clk_0_W_in(prog_clk_0_wires[351]),
    .Reset_E_out(ResetWires[195]),
    .Reset_W_in(ResetWires[194]),
    .pReset_S_in(pResetWires[391]),
    .Test_en_E_out(Test_enWires[195]),
    .Test_en_W_in(Test_enWires[194]),
    .chany_bottom_in(sb_1__1__94_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__95_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_103_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__103_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__103_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__103_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__103_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__103_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__103_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__103_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__103_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__103_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__103_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__103_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__103_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__103_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__103_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__103_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__103_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__103_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__103_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__103_ccff_tail[0])
  );


  cby_1__1_
  cby_9__9_
  (
    .clk_2_N_out(clk_2_wires[100]),
    .clk_2_S_in(clk_2_wires[99]),
    .prog_clk_2_N_out(prog_clk_2_wires[100]),
    .prog_clk_2_S_in(prog_clk_2_wires[99]),
    .prog_clk_0_S_out(prog_clk_0_wires[355]),
    .prog_clk_0_W_in(prog_clk_0_wires[354]),
    .Reset_E_out(ResetWires[217]),
    .Reset_W_in(ResetWires[216]),
    .pReset_S_in(pResetWires[440]),
    .Test_en_E_out(Test_enWires[217]),
    .Test_en_W_in(Test_enWires[216]),
    .chany_bottom_in(sb_1__1__95_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__96_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_104_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__104_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__104_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__104_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__104_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__104_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__104_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__104_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__104_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__104_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__104_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__104_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__104_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__104_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__104_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__104_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__104_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__104_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__104_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__104_ccff_tail[0])
  );


  cby_1__1_
  cby_9__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[358]),
    .prog_clk_0_W_in(prog_clk_0_wires[357]),
    .Reset_E_out(ResetWires[239]),
    .Reset_W_in(ResetWires[238]),
    .pReset_S_in(pResetWires[489]),
    .Test_en_E_out(Test_enWires[239]),
    .Test_en_W_in(Test_enWires[238]),
    .chany_bottom_in(sb_1__1__96_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__97_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_105_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__105_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__105_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__105_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__105_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__105_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__105_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__105_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__105_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__105_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__105_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__105_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__105_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__105_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__105_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__105_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__105_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__105_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__105_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__105_ccff_tail[0])
  );


  cby_1__1_
  cby_9__11_
  (
    .clk_2_N_out(clk_2_wires[111]),
    .clk_2_S_in(clk_2_wires[110]),
    .prog_clk_2_N_out(prog_clk_2_wires[111]),
    .prog_clk_2_S_in(prog_clk_2_wires[110]),
    .prog_clk_0_S_out(prog_clk_0_wires[361]),
    .prog_clk_0_W_in(prog_clk_0_wires[360]),
    .Reset_E_out(ResetWires[261]),
    .Reset_W_in(ResetWires[260]),
    .pReset_S_in(pResetWires[538]),
    .Test_en_E_out(Test_enWires[261]),
    .Test_en_W_in(Test_enWires[260]),
    .chany_bottom_in(sb_1__1__97_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__98_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_106_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__106_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__106_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__106_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__106_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__106_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__106_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__106_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__106_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__106_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__106_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__106_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__106_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__106_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__106_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__106_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__106_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__106_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__106_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__106_ccff_tail[0])
  );


  cby_1__1_
  cby_9__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[366]),
    .prog_clk_0_S_out(prog_clk_0_wires[364]),
    .prog_clk_0_W_in(prog_clk_0_wires[363]),
    .Reset_E_out(ResetWires[283]),
    .Reset_W_in(ResetWires[282]),
    .pReset_S_in(pResetWires[587]),
    .Test_en_E_out(Test_enWires[283]),
    .Test_en_W_in(Test_enWires[282]),
    .chany_bottom_in(sb_1__1__98_chany_top_out[0:29]),
    .chany_top_in(sb_1__12__8_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_107_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__107_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__107_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__107_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__107_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__107_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__107_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__107_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__107_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__107_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__107_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__107_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__107_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__107_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__107_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__107_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__107_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__107_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__107_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__107_ccff_tail[0])
  );


  cby_1__1_
  cby_10__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[369]),
    .prog_clk_0_W_in(prog_clk_0_wires[368]),
    .Reset_E_out(ResetWires[43]),
    .Reset_W_in(ResetWires[42]),
    .pReset_S_in(pResetWires[54]),
    .Test_en_E_out(Test_enWires[43]),
    .Test_en_W_in(Test_enWires[42]),
    .chany_bottom_in(sb_1__0__9_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__99_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_108_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__108_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__108_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__108_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__108_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__108_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__108_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__108_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__108_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__108_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__108_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__108_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__108_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__108_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__108_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__108_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__108_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__108_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__108_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__108_ccff_tail[0])
  );


  cby_1__1_
  cby_10__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[372]),
    .prog_clk_0_W_in(prog_clk_0_wires[371]),
    .Reset_E_out(ResetWires[65]),
    .Reset_W_in(ResetWires[64]),
    .pReset_S_in(pResetWires[101]),
    .Test_en_E_out(Test_enWires[65]),
    .Test_en_W_in(Test_enWires[64]),
    .chany_bottom_in(sb_1__1__99_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__100_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_109_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__109_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__109_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__109_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__109_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__109_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__109_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__109_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__109_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__109_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__109_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__109_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__109_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__109_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__109_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__109_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__109_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__109_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__109_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__109_ccff_tail[0])
  );


  cby_1__1_
  cby_10__3_
  (
    .clk_3_S_out(clk_3_wires[87]),
    .clk_3_N_in(clk_3_wires[86]),
    .prog_clk_3_S_out(prog_clk_3_wires[87]),
    .prog_clk_3_N_in(prog_clk_3_wires[86]),
    .prog_clk_0_S_out(prog_clk_0_wires[375]),
    .prog_clk_0_W_in(prog_clk_0_wires[374]),
    .Reset_E_out(ResetWires[87]),
    .Reset_W_in(ResetWires[86]),
    .pReset_S_in(pResetWires[150]),
    .Test_en_E_out(Test_enWires[87]),
    .Test_en_W_in(Test_enWires[86]),
    .chany_bottom_in(sb_1__1__100_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__101_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_110_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__110_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__110_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__110_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__110_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__110_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__110_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__110_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__110_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__110_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__110_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__110_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__110_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__110_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__110_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__110_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__110_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__110_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__110_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__110_ccff_tail[0])
  );


  cby_1__1_
  cby_10__4_
  (
    .clk_3_S_out(clk_3_wires[83]),
    .clk_3_N_in(clk_3_wires[82]),
    .prog_clk_3_S_out(prog_clk_3_wires[83]),
    .prog_clk_3_N_in(prog_clk_3_wires[82]),
    .prog_clk_0_S_out(prog_clk_0_wires[378]),
    .prog_clk_0_W_in(prog_clk_0_wires[377]),
    .Reset_E_out(ResetWires[109]),
    .Reset_W_in(ResetWires[108]),
    .pReset_S_in(pResetWires[199]),
    .Test_en_E_out(Test_enWires[109]),
    .Test_en_W_in(Test_enWires[108]),
    .chany_bottom_in(sb_1__1__101_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__102_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_111_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__111_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__111_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__111_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__111_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__111_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__111_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__111_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__111_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__111_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__111_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__111_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__111_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__111_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__111_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__111_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__111_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__111_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__111_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__111_ccff_tail[0])
  );


  cby_1__1_
  cby_10__5_
  (
    .clk_3_S_out(clk_3_wires[77]),
    .clk_3_N_in(clk_3_wires[76]),
    .prog_clk_3_S_out(prog_clk_3_wires[77]),
    .prog_clk_3_N_in(prog_clk_3_wires[76]),
    .prog_clk_0_S_out(prog_clk_0_wires[381]),
    .prog_clk_0_W_in(prog_clk_0_wires[380]),
    .Reset_E_out(ResetWires[131]),
    .Reset_W_in(ResetWires[130]),
    .pReset_S_in(pResetWires[248]),
    .Test_en_E_out(Test_enWires[131]),
    .Test_en_W_in(Test_enWires[130]),
    .chany_bottom_in(sb_1__1__102_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__103_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_112_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__112_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__112_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__112_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__112_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__112_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__112_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__112_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__112_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__112_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__112_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__112_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__112_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__112_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__112_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__112_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__112_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__112_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__112_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__112_ccff_tail[0])
  );


  cby_1__1_
  cby_10__6_
  (
    .clk_3_S_out(clk_3_wires[73]),
    .clk_3_N_in(clk_3_wires[72]),
    .prog_clk_3_S_out(prog_clk_3_wires[73]),
    .prog_clk_3_N_in(prog_clk_3_wires[72]),
    .prog_clk_0_S_out(prog_clk_0_wires[384]),
    .prog_clk_0_W_in(prog_clk_0_wires[383]),
    .Reset_E_out(ResetWires[153]),
    .Reset_W_in(ResetWires[152]),
    .pReset_S_in(pResetWires[297]),
    .Test_en_E_out(Test_enWires[153]),
    .Test_en_W_in(Test_enWires[152]),
    .chany_bottom_in(sb_1__1__103_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__104_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_113_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__113_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__113_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__113_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__113_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__113_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__113_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__113_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__113_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__113_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__113_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__113_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__113_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__113_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__113_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__113_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__113_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__113_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__113_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__113_ccff_tail[0])
  );


  cby_1__1_
  cby_10__7_
  (
    .clk_3_N_out(clk_3_wires[71]),
    .clk_3_S_in(clk_3_wires[70]),
    .prog_clk_3_N_out(prog_clk_3_wires[71]),
    .prog_clk_3_S_in(prog_clk_3_wires[70]),
    .prog_clk_0_S_out(prog_clk_0_wires[387]),
    .prog_clk_0_W_in(prog_clk_0_wires[386]),
    .Reset_E_out(ResetWires[175]),
    .Reset_W_in(ResetWires[174]),
    .pReset_S_in(pResetWires[346]),
    .Test_en_E_out(Test_enWires[175]),
    .Test_en_W_in(Test_enWires[174]),
    .chany_bottom_in(sb_1__1__104_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__105_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_114_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__114_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__114_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__114_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__114_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__114_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__114_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__114_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__114_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__114_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__114_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__114_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__114_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__114_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__114_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__114_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__114_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__114_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__114_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__114_ccff_tail[0])
  );


  cby_1__1_
  cby_10__8_
  (
    .clk_3_N_out(clk_3_wires[75]),
    .clk_3_S_in(clk_3_wires[74]),
    .prog_clk_3_N_out(prog_clk_3_wires[75]),
    .prog_clk_3_S_in(prog_clk_3_wires[74]),
    .prog_clk_0_S_out(prog_clk_0_wires[390]),
    .prog_clk_0_W_in(prog_clk_0_wires[389]),
    .Reset_E_out(ResetWires[197]),
    .Reset_W_in(ResetWires[196]),
    .pReset_S_in(pResetWires[395]),
    .Test_en_E_out(Test_enWires[197]),
    .Test_en_W_in(Test_enWires[196]),
    .chany_bottom_in(sb_1__1__105_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__106_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_115_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__115_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__115_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__115_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__115_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__115_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__115_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__115_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__115_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__115_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__115_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__115_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__115_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__115_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__115_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__115_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__115_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__115_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__115_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__115_ccff_tail[0])
  );


  cby_1__1_
  cby_10__9_
  (
    .clk_3_N_out(clk_3_wires[81]),
    .clk_3_S_in(clk_3_wires[80]),
    .prog_clk_3_N_out(prog_clk_3_wires[81]),
    .prog_clk_3_S_in(prog_clk_3_wires[80]),
    .prog_clk_0_S_out(prog_clk_0_wires[393]),
    .prog_clk_0_W_in(prog_clk_0_wires[392]),
    .Reset_E_out(ResetWires[219]),
    .Reset_W_in(ResetWires[218]),
    .pReset_S_in(pResetWires[444]),
    .Test_en_E_out(Test_enWires[219]),
    .Test_en_W_in(Test_enWires[218]),
    .chany_bottom_in(sb_1__1__106_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__107_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_116_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__116_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__116_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__116_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__116_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__116_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__116_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__116_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__116_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__116_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__116_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__116_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__116_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__116_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__116_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__116_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__116_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__116_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__116_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__116_ccff_tail[0])
  );


  cby_1__1_
  cby_10__10_
  (
    .clk_3_N_out(clk_3_wires[85]),
    .clk_3_S_in(clk_3_wires[84]),
    .prog_clk_3_N_out(prog_clk_3_wires[85]),
    .prog_clk_3_S_in(prog_clk_3_wires[84]),
    .prog_clk_0_S_out(prog_clk_0_wires[396]),
    .prog_clk_0_W_in(prog_clk_0_wires[395]),
    .Reset_E_out(ResetWires[241]),
    .Reset_W_in(ResetWires[240]),
    .pReset_S_in(pResetWires[493]),
    .Test_en_E_out(Test_enWires[241]),
    .Test_en_W_in(Test_enWires[240]),
    .chany_bottom_in(sb_1__1__107_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__108_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_117_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__117_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__117_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__117_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__117_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__117_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__117_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__117_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__117_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__117_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__117_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__117_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__117_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__117_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__117_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__117_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__117_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__117_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__117_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__117_ccff_tail[0])
  );


  cby_1__1_
  cby_10__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[399]),
    .prog_clk_0_W_in(prog_clk_0_wires[398]),
    .Reset_E_out(ResetWires[263]),
    .Reset_W_in(ResetWires[262]),
    .pReset_S_in(pResetWires[542]),
    .Test_en_E_out(Test_enWires[263]),
    .Test_en_W_in(Test_enWires[262]),
    .chany_bottom_in(sb_1__1__108_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__109_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_118_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__118_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__118_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__118_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__118_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__118_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__118_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__118_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__118_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__118_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__118_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__118_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__118_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__118_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__118_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__118_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__118_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__118_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__118_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__118_ccff_tail[0])
  );


  cby_1__1_
  cby_10__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[404]),
    .prog_clk_0_S_out(prog_clk_0_wires[402]),
    .prog_clk_0_W_in(prog_clk_0_wires[401]),
    .Reset_E_out(ResetWires[285]),
    .Reset_W_in(ResetWires[284]),
    .pReset_S_in(pResetWires[591]),
    .Test_en_E_out(Test_enWires[285]),
    .Test_en_W_in(Test_enWires[284]),
    .chany_bottom_in(sb_1__1__109_chany_top_out[0:29]),
    .chany_top_in(sb_1__12__9_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_119_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__119_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__119_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__119_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__119_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__119_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__119_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__119_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__119_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__119_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__119_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__119_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__119_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__119_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__119_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__119_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__119_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__119_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__119_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__119_ccff_tail[0])
  );


  cby_1__1_
  cby_11__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[407]),
    .prog_clk_0_W_in(prog_clk_0_wires[406]),
    .Reset_E_out(ResetWires[45]),
    .Reset_W_in(ResetWires[44]),
    .pReset_S_in(pResetWires[57]),
    .Test_en_E_out(Test_enWires[45]),
    .Test_en_W_in(Test_enWires[44]),
    .chany_bottom_in(sb_1__0__10_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__110_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_120_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__120_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__120_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__120_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__120_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__120_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__120_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__120_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__120_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__120_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__120_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__120_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__120_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__120_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__120_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__120_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__120_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__120_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__120_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__120_ccff_tail[0])
  );


  cby_1__1_
  cby_11__2_
  (
    .clk_2_S_out(clk_2_wires[116]),
    .clk_2_N_in(clk_2_wires[115]),
    .prog_clk_2_S_out(prog_clk_2_wires[116]),
    .prog_clk_2_N_in(prog_clk_2_wires[115]),
    .prog_clk_0_S_out(prog_clk_0_wires[410]),
    .prog_clk_0_W_in(prog_clk_0_wires[409]),
    .Reset_E_out(ResetWires[67]),
    .Reset_W_in(ResetWires[66]),
    .pReset_S_in(pResetWires[105]),
    .Test_en_E_out(Test_enWires[67]),
    .Test_en_W_in(Test_enWires[66]),
    .chany_bottom_in(sb_1__1__110_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__111_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_121_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__121_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__121_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__121_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__121_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__121_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__121_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__121_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__121_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__121_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__121_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__121_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__121_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__121_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__121_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__121_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__121_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__121_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__121_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__121_ccff_tail[0])
  );


  cby_1__1_
  cby_11__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[413]),
    .prog_clk_0_W_in(prog_clk_0_wires[412]),
    .Reset_E_out(ResetWires[89]),
    .Reset_W_in(ResetWires[88]),
    .pReset_S_in(pResetWires[154]),
    .Test_en_E_out(Test_enWires[89]),
    .Test_en_W_in(Test_enWires[88]),
    .chany_bottom_in(sb_1__1__111_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__112_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_122_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__122_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__122_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__122_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__122_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__122_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__122_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__122_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__122_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__122_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__122_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__122_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__122_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__122_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__122_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__122_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__122_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__122_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__122_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__122_ccff_tail[0])
  );


  cby_1__1_
  cby_11__4_
  (
    .clk_2_S_out(clk_2_wires[123]),
    .clk_2_N_in(clk_2_wires[122]),
    .prog_clk_2_S_out(prog_clk_2_wires[123]),
    .prog_clk_2_N_in(prog_clk_2_wires[122]),
    .prog_clk_0_S_out(prog_clk_0_wires[416]),
    .prog_clk_0_W_in(prog_clk_0_wires[415]),
    .Reset_E_out(ResetWires[111]),
    .Reset_W_in(ResetWires[110]),
    .pReset_S_in(pResetWires[203]),
    .Test_en_E_out(Test_enWires[111]),
    .Test_en_W_in(Test_enWires[110]),
    .chany_bottom_in(sb_1__1__112_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__113_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_123_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__123_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__123_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__123_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__123_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__123_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__123_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__123_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__123_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__123_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__123_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__123_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__123_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__123_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__123_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__123_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__123_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__123_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__123_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__123_ccff_tail[0])
  );


  cby_1__1_
  cby_11__5_
  (
    .clk_2_N_out(clk_2_wires[121]),
    .clk_2_S_in(clk_2_wires[120]),
    .prog_clk_2_N_out(prog_clk_2_wires[121]),
    .prog_clk_2_S_in(prog_clk_2_wires[120]),
    .prog_clk_0_S_out(prog_clk_0_wires[419]),
    .prog_clk_0_W_in(prog_clk_0_wires[418]),
    .Reset_E_out(ResetWires[133]),
    .Reset_W_in(ResetWires[132]),
    .pReset_S_in(pResetWires[252]),
    .Test_en_E_out(Test_enWires[133]),
    .Test_en_W_in(Test_enWires[132]),
    .chany_bottom_in(sb_1__1__113_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__114_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_124_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__124_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__124_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__124_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__124_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__124_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__124_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__124_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__124_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__124_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__124_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__124_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__124_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__124_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__124_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__124_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__124_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__124_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__124_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__124_ccff_tail[0])
  );


  cby_1__1_
  cby_11__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[422]),
    .prog_clk_0_W_in(prog_clk_0_wires[421]),
    .Reset_E_out(ResetWires[155]),
    .Reset_W_in(ResetWires[154]),
    .pReset_S_in(pResetWires[301]),
    .Test_en_E_out(Test_enWires[155]),
    .Test_en_W_in(Test_enWires[154]),
    .chany_bottom_in(sb_1__1__114_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__115_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_125_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__125_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__125_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__125_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__125_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__125_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__125_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__125_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__125_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__125_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__125_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__125_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__125_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__125_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__125_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__125_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__125_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__125_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__125_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__125_ccff_tail[0])
  );


  cby_1__1_
  cby_11__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[425]),
    .prog_clk_0_W_in(prog_clk_0_wires[424]),
    .Reset_E_out(ResetWires[177]),
    .Reset_W_in(ResetWires[176]),
    .pReset_S_in(pResetWires[350]),
    .Test_en_E_out(Test_enWires[177]),
    .Test_en_W_in(Test_enWires[176]),
    .chany_bottom_in(sb_1__1__115_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__116_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_126_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__126_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__126_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__126_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__126_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__126_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__126_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__126_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__126_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__126_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__126_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__126_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__126_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__126_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__126_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__126_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__126_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__126_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__126_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__126_ccff_tail[0])
  );


  cby_1__1_
  cby_11__8_
  (
    .clk_2_S_out(clk_2_wires[130]),
    .clk_2_N_in(clk_2_wires[129]),
    .prog_clk_2_S_out(prog_clk_2_wires[130]),
    .prog_clk_2_N_in(prog_clk_2_wires[129]),
    .prog_clk_0_S_out(prog_clk_0_wires[428]),
    .prog_clk_0_W_in(prog_clk_0_wires[427]),
    .Reset_E_out(ResetWires[199]),
    .Reset_W_in(ResetWires[198]),
    .pReset_S_in(pResetWires[399]),
    .Test_en_E_out(Test_enWires[199]),
    .Test_en_W_in(Test_enWires[198]),
    .chany_bottom_in(sb_1__1__116_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__117_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_127_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__127_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__127_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__127_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__127_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__127_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__127_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__127_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__127_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__127_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__127_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__127_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__127_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__127_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__127_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__127_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__127_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__127_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__127_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__127_ccff_tail[0])
  );


  cby_1__1_
  cby_11__9_
  (
    .clk_2_N_out(clk_2_wires[128]),
    .clk_2_S_in(clk_2_wires[127]),
    .prog_clk_2_N_out(prog_clk_2_wires[128]),
    .prog_clk_2_S_in(prog_clk_2_wires[127]),
    .prog_clk_0_S_out(prog_clk_0_wires[431]),
    .prog_clk_0_W_in(prog_clk_0_wires[430]),
    .Reset_E_out(ResetWires[221]),
    .Reset_W_in(ResetWires[220]),
    .pReset_S_in(pResetWires[448]),
    .Test_en_E_out(Test_enWires[221]),
    .Test_en_W_in(Test_enWires[220]),
    .chany_bottom_in(sb_1__1__117_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__118_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_128_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__128_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__128_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__128_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__128_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__128_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__128_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__128_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__128_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__128_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__128_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__128_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__128_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__128_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__128_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__128_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__128_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__128_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__128_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__128_ccff_tail[0])
  );


  cby_1__1_
  cby_11__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[434]),
    .prog_clk_0_W_in(prog_clk_0_wires[433]),
    .Reset_E_out(ResetWires[243]),
    .Reset_W_in(ResetWires[242]),
    .pReset_S_in(pResetWires[497]),
    .Test_en_E_out(Test_enWires[243]),
    .Test_en_W_in(Test_enWires[242]),
    .chany_bottom_in(sb_1__1__118_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__119_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_129_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__129_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__129_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__129_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__129_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__129_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__129_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__129_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__129_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__129_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__129_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__129_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__129_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__129_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__129_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__129_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__129_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__129_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__129_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__129_ccff_tail[0])
  );


  cby_1__1_
  cby_11__11_
  (
    .clk_2_N_out(clk_2_wires[135]),
    .clk_2_S_in(clk_2_wires[134]),
    .prog_clk_2_N_out(prog_clk_2_wires[135]),
    .prog_clk_2_S_in(prog_clk_2_wires[134]),
    .prog_clk_0_S_out(prog_clk_0_wires[437]),
    .prog_clk_0_W_in(prog_clk_0_wires[436]),
    .Reset_E_out(ResetWires[265]),
    .Reset_W_in(ResetWires[264]),
    .pReset_S_in(pResetWires[546]),
    .Test_en_E_out(Test_enWires[265]),
    .Test_en_W_in(Test_enWires[264]),
    .chany_bottom_in(sb_1__1__119_chany_top_out[0:29]),
    .chany_top_in(sb_1__1__120_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_130_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__130_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__130_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__130_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__130_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__130_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__130_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__130_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__130_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__130_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__130_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__130_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__130_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__130_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__130_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__130_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__130_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__130_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__130_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__130_ccff_tail[0])
  );


  cby_1__1_
  cby_11__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[442]),
    .prog_clk_0_S_out(prog_clk_0_wires[440]),
    .prog_clk_0_W_in(prog_clk_0_wires[439]),
    .Reset_E_out(ResetWires[287]),
    .Reset_W_in(ResetWires[286]),
    .pReset_S_in(pResetWires[595]),
    .Test_en_E_out(Test_enWires[287]),
    .Test_en_W_in(Test_enWires[286]),
    .chany_bottom_in(sb_1__1__120_chany_top_out[0:29]),
    .chany_top_in(sb_1__12__10_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_131_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__131_chany_bottom_out[0:29]),
    .chany_top_out(cby_1__1__131_chany_top_out[0:29]),
    .left_grid_pin_16_(cby_1__1__131_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__131_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__131_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__131_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__131_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__131_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__131_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__131_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__131_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__131_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__131_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__131_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__131_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__131_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__131_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__131_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__131_ccff_tail[0])
  );


  cby_2__1_
  cby_12__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[445]),
    .prog_clk_0_W_in(prog_clk_0_wires[444]),
    .pReset_S_in(pResetWires[60]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_11_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_11_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__0_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__0__0_chany_top_out[0:29]),
    .chany_top_in(sb_12__1__0_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_132_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__0_chany_bottom_out[0:29]),
    .chany_top_out(cby_12__1__0_chany_top_out[0:29]),
    .right_grid_pin_0_(cby_12__1__0_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__0_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__0_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__0_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__0_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__0_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__0_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__0_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__0_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__0_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__0_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__0_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__0_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__0_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__0_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__0_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__0_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_11_ccff_tail[0])
  );


  cby_2__1_
  cby_12__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[448]),
    .prog_clk_0_W_in(prog_clk_0_wires[447]),
    .pReset_S_in(pResetWires[109]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_10_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_10_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__1_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__0_chany_top_out[0:29]),
    .chany_top_in(sb_12__1__1_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_133_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__1_chany_bottom_out[0:29]),
    .chany_top_out(cby_12__1__1_chany_top_out[0:29]),
    .right_grid_pin_0_(cby_12__1__1_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__1_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__1_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__1_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__1_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__1_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__1_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__1_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__1_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__1_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__1_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__1_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__1_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__1_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__1_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__1_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__1_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_10_ccff_tail[0])
  );


  cby_2__1_
  cby_12__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[451]),
    .prog_clk_0_W_in(prog_clk_0_wires[450]),
    .pReset_S_in(pResetWires[158]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_9_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_9_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__2_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__1_chany_top_out[0:29]),
    .chany_top_in(sb_12__1__2_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_134_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__2_chany_bottom_out[0:29]),
    .chany_top_out(cby_12__1__2_chany_top_out[0:29]),
    .right_grid_pin_0_(cby_12__1__2_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__2_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__2_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__2_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__2_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__2_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__2_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__2_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__2_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__2_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__2_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__2_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__2_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__2_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__2_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__2_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__2_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_9_ccff_tail[0])
  );


  cby_2__1_
  cby_12__4_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[454]),
    .prog_clk_0_W_in(prog_clk_0_wires[453]),
    .pReset_S_in(pResetWires[207]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_8_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_8_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__3_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__2_chany_top_out[0:29]),
    .chany_top_in(sb_12__1__3_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_135_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__3_chany_bottom_out[0:29]),
    .chany_top_out(cby_12__1__3_chany_top_out[0:29]),
    .right_grid_pin_0_(cby_12__1__3_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__3_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__3_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__3_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__3_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__3_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__3_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__3_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__3_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__3_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__3_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__3_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__3_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__3_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__3_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__3_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__3_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_8_ccff_tail[0])
  );


  cby_2__1_
  cby_12__5_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[457]),
    .prog_clk_0_W_in(prog_clk_0_wires[456]),
    .pReset_S_in(pResetWires[256]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_7_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_7_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__4_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__3_chany_top_out[0:29]),
    .chany_top_in(sb_12__1__4_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_136_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__4_chany_bottom_out[0:29]),
    .chany_top_out(cby_12__1__4_chany_top_out[0:29]),
    .right_grid_pin_0_(cby_12__1__4_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__4_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__4_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__4_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__4_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__4_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__4_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__4_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__4_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__4_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__4_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__4_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__4_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__4_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__4_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__4_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__4_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_7_ccff_tail[0])
  );


  cby_2__1_
  cby_12__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[460]),
    .prog_clk_0_W_in(prog_clk_0_wires[459]),
    .pReset_S_in(pResetWires[305]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_6_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_6_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__5_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__4_chany_top_out[0:29]),
    .chany_top_in(sb_12__1__5_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_137_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__5_chany_bottom_out[0:29]),
    .chany_top_out(cby_12__1__5_chany_top_out[0:29]),
    .right_grid_pin_0_(cby_12__1__5_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__5_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__5_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__5_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__5_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__5_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__5_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__5_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__5_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__5_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__5_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__5_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__5_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__5_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__5_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__5_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__5_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_6_ccff_tail[0])
  );


  cby_2__1_
  cby_12__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[463]),
    .prog_clk_0_W_in(prog_clk_0_wires[462]),
    .pReset_S_in(pResetWires[354]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_5_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_5_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__6_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__5_chany_top_out[0:29]),
    .chany_top_in(sb_12__1__6_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_138_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__6_chany_bottom_out[0:29]),
    .chany_top_out(cby_12__1__6_chany_top_out[0:29]),
    .right_grid_pin_0_(cby_12__1__6_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__6_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__6_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__6_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__6_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__6_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__6_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__6_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__6_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__6_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__6_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__6_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__6_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__6_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__6_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__6_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__6_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_5_ccff_tail[0])
  );


  cby_2__1_
  cby_12__8_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[466]),
    .prog_clk_0_W_in(prog_clk_0_wires[465]),
    .pReset_S_in(pResetWires[403]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_4_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_4_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__7_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__6_chany_top_out[0:29]),
    .chany_top_in(sb_12__1__7_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_139_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__7_chany_bottom_out[0:29]),
    .chany_top_out(cby_12__1__7_chany_top_out[0:29]),
    .right_grid_pin_0_(cby_12__1__7_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__7_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__7_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__7_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__7_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__7_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__7_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__7_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__7_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__7_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__7_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__7_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__7_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__7_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__7_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__7_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__7_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_4_ccff_tail[0])
  );


  cby_2__1_
  cby_12__9_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[469]),
    .prog_clk_0_W_in(prog_clk_0_wires[468]),
    .pReset_S_in(pResetWires[452]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_3_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_3_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__8_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__7_chany_top_out[0:29]),
    .chany_top_in(sb_12__1__8_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_140_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__8_chany_bottom_out[0:29]),
    .chany_top_out(cby_12__1__8_chany_top_out[0:29]),
    .right_grid_pin_0_(cby_12__1__8_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__8_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__8_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__8_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__8_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__8_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__8_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__8_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__8_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__8_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__8_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__8_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__8_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__8_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__8_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__8_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__8_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_3_ccff_tail[0])
  );


  cby_2__1_
  cby_12__10_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[472]),
    .prog_clk_0_W_in(prog_clk_0_wires[471]),
    .pReset_S_in(pResetWires[501]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_2_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_2_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__9_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__8_chany_top_out[0:29]),
    .chany_top_in(sb_12__1__9_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_141_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__9_chany_bottom_out[0:29]),
    .chany_top_out(cby_12__1__9_chany_top_out[0:29]),
    .right_grid_pin_0_(cby_12__1__9_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__9_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__9_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__9_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__9_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__9_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__9_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__9_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__9_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__9_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__9_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__9_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__9_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__9_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__9_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__9_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__9_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_2_ccff_tail[0])
  );


  cby_2__1_
  cby_12__11_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[475]),
    .prog_clk_0_W_in(prog_clk_0_wires[474]),
    .pReset_S_in(pResetWires[550]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_1_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_1_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__10_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__9_chany_top_out[0:29]),
    .chany_top_in(sb_12__1__10_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_142_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__10_chany_bottom_out[0:29]),
    .chany_top_out(cby_12__1__10_chany_top_out[0:29]),
    .right_grid_pin_0_(cby_12__1__10_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__10_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__10_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__10_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__10_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__10_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__10_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__10_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__10_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__10_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__10_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__10_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__10_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__10_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__10_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__10_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__10_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_1_ccff_tail[0])
  );


  cby_2__1_
  cby_12__12_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[480]),
    .prog_clk_0_S_out(prog_clk_0_wires[478]),
    .prog_clk_0_W_in(prog_clk_0_wires[477]),
    .pReset_S_in(pResetWires[599]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_0_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_0_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_12__1__11_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_12__1__10_chany_top_out[0:29]),
    .chany_top_in(sb_12__12__0_chany_bottom_out[0:29]),
    .ccff_head(grid_clb_143_ccff_tail[0]),
    .chany_bottom_out(cby_12__1__11_chany_bottom_out[0:29]),
    .chany_top_out(cby_12__1__11_chany_top_out[0:29]),
    .right_grid_pin_0_(cby_12__1__11_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_12__1__11_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_12__1__11_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_12__1__11_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_12__1__11_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_12__1__11_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_12__1__11_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_12__1__11_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_12__1__11_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_12__1__11_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_12__1__11_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_12__1__11_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_12__1__11_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_12__1__11_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_12__1__11_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_12__1__11_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_12__1__11_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_0_ccff_tail[0])
  );


  direct_interc
  direct_interc_0_
  (
    .in(grid_clb_1_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_0_out[0])
  );


  direct_interc
  direct_interc_1_
  (
    .in(grid_clb_2_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_1_out[0])
  );


  direct_interc
  direct_interc_2_
  (
    .in(grid_clb_3_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_2_out[0])
  );


  direct_interc
  direct_interc_3_
  (
    .in(grid_clb_4_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_3_out[0])
  );


  direct_interc
  direct_interc_4_
  (
    .in(grid_clb_5_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_4_out[0])
  );


  direct_interc
  direct_interc_5_
  (
    .in(grid_clb_6_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_5_out[0])
  );


  direct_interc
  direct_interc_6_
  (
    .in(grid_clb_7_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_6_out[0])
  );


  direct_interc
  direct_interc_7_
  (
    .in(grid_clb_8_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_7_out[0])
  );


  direct_interc
  direct_interc_8_
  (
    .in(grid_clb_9_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_8_out[0])
  );


  direct_interc
  direct_interc_9_
  (
    .in(grid_clb_10_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_9_out[0])
  );


  direct_interc
  direct_interc_10_
  (
    .in(grid_clb_11_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_10_out[0])
  );


  direct_interc
  direct_interc_11_
  (
    .in(grid_clb_13_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_11_out[0])
  );


  direct_interc
  direct_interc_12_
  (
    .in(grid_clb_14_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_12_out[0])
  );


  direct_interc
  direct_interc_13_
  (
    .in(grid_clb_15_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_13_out[0])
  );


  direct_interc
  direct_interc_14_
  (
    .in(grid_clb_16_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_14_out[0])
  );


  direct_interc
  direct_interc_15_
  (
    .in(grid_clb_17_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_15_out[0])
  );


  direct_interc
  direct_interc_16_
  (
    .in(grid_clb_18_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_16_out[0])
  );


  direct_interc
  direct_interc_17_
  (
    .in(grid_clb_19_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_17_out[0])
  );


  direct_interc
  direct_interc_18_
  (
    .in(grid_clb_20_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_18_out[0])
  );


  direct_interc
  direct_interc_19_
  (
    .in(grid_clb_21_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_19_out[0])
  );


  direct_interc
  direct_interc_20_
  (
    .in(grid_clb_22_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_20_out[0])
  );


  direct_interc
  direct_interc_21_
  (
    .in(grid_clb_23_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_21_out[0])
  );


  direct_interc
  direct_interc_22_
  (
    .in(grid_clb_25_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_22_out[0])
  );


  direct_interc
  direct_interc_23_
  (
    .in(grid_clb_26_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_23_out[0])
  );


  direct_interc
  direct_interc_24_
  (
    .in(grid_clb_27_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_24_out[0])
  );


  direct_interc
  direct_interc_25_
  (
    .in(grid_clb_28_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_25_out[0])
  );


  direct_interc
  direct_interc_26_
  (
    .in(grid_clb_29_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_26_out[0])
  );


  direct_interc
  direct_interc_27_
  (
    .in(grid_clb_30_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_27_out[0])
  );


  direct_interc
  direct_interc_28_
  (
    .in(grid_clb_31_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_28_out[0])
  );


  direct_interc
  direct_interc_29_
  (
    .in(grid_clb_32_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_29_out[0])
  );


  direct_interc
  direct_interc_30_
  (
    .in(grid_clb_33_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_30_out[0])
  );


  direct_interc
  direct_interc_31_
  (
    .in(grid_clb_34_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_31_out[0])
  );


  direct_interc
  direct_interc_32_
  (
    .in(grid_clb_35_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_32_out[0])
  );


  direct_interc
  direct_interc_33_
  (
    .in(grid_clb_37_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_33_out[0])
  );


  direct_interc
  direct_interc_34_
  (
    .in(grid_clb_38_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_34_out[0])
  );


  direct_interc
  direct_interc_35_
  (
    .in(grid_clb_39_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_35_out[0])
  );


  direct_interc
  direct_interc_36_
  (
    .in(grid_clb_40_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_36_out[0])
  );


  direct_interc
  direct_interc_37_
  (
    .in(grid_clb_41_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_37_out[0])
  );


  direct_interc
  direct_interc_38_
  (
    .in(grid_clb_42_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_38_out[0])
  );


  direct_interc
  direct_interc_39_
  (
    .in(grid_clb_43_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_39_out[0])
  );


  direct_interc
  direct_interc_40_
  (
    .in(grid_clb_44_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_40_out[0])
  );


  direct_interc
  direct_interc_41_
  (
    .in(grid_clb_45_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_41_out[0])
  );


  direct_interc
  direct_interc_42_
  (
    .in(grid_clb_46_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_42_out[0])
  );


  direct_interc
  direct_interc_43_
  (
    .in(grid_clb_47_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_43_out[0])
  );


  direct_interc
  direct_interc_44_
  (
    .in(grid_clb_49_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_44_out[0])
  );


  direct_interc
  direct_interc_45_
  (
    .in(grid_clb_50_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_45_out[0])
  );


  direct_interc
  direct_interc_46_
  (
    .in(grid_clb_51_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_46_out[0])
  );


  direct_interc
  direct_interc_47_
  (
    .in(grid_clb_52_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_47_out[0])
  );


  direct_interc
  direct_interc_48_
  (
    .in(grid_clb_53_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_48_out[0])
  );


  direct_interc
  direct_interc_49_
  (
    .in(grid_clb_54_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_49_out[0])
  );


  direct_interc
  direct_interc_50_
  (
    .in(grid_clb_55_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_50_out[0])
  );


  direct_interc
  direct_interc_51_
  (
    .in(grid_clb_56_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_51_out[0])
  );


  direct_interc
  direct_interc_52_
  (
    .in(grid_clb_57_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_52_out[0])
  );


  direct_interc
  direct_interc_53_
  (
    .in(grid_clb_58_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_53_out[0])
  );


  direct_interc
  direct_interc_54_
  (
    .in(grid_clb_59_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_54_out[0])
  );


  direct_interc
  direct_interc_55_
  (
    .in(grid_clb_61_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_55_out[0])
  );


  direct_interc
  direct_interc_56_
  (
    .in(grid_clb_62_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_56_out[0])
  );


  direct_interc
  direct_interc_57_
  (
    .in(grid_clb_63_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_57_out[0])
  );


  direct_interc
  direct_interc_58_
  (
    .in(grid_clb_64_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_58_out[0])
  );


  direct_interc
  direct_interc_59_
  (
    .in(grid_clb_65_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_59_out[0])
  );


  direct_interc
  direct_interc_60_
  (
    .in(grid_clb_66_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_60_out[0])
  );


  direct_interc
  direct_interc_61_
  (
    .in(grid_clb_67_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_61_out[0])
  );


  direct_interc
  direct_interc_62_
  (
    .in(grid_clb_68_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_62_out[0])
  );


  direct_interc
  direct_interc_63_
  (
    .in(grid_clb_69_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_63_out[0])
  );


  direct_interc
  direct_interc_64_
  (
    .in(grid_clb_70_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_64_out[0])
  );


  direct_interc
  direct_interc_65_
  (
    .in(grid_clb_71_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_65_out[0])
  );


  direct_interc
  direct_interc_66_
  (
    .in(grid_clb_73_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_66_out[0])
  );


  direct_interc
  direct_interc_67_
  (
    .in(grid_clb_74_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_67_out[0])
  );


  direct_interc
  direct_interc_68_
  (
    .in(grid_clb_75_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_68_out[0])
  );


  direct_interc
  direct_interc_69_
  (
    .in(grid_clb_76_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_69_out[0])
  );


  direct_interc
  direct_interc_70_
  (
    .in(grid_clb_77_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_70_out[0])
  );


  direct_interc
  direct_interc_71_
  (
    .in(grid_clb_78_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_71_out[0])
  );


  direct_interc
  direct_interc_72_
  (
    .in(grid_clb_79_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_72_out[0])
  );


  direct_interc
  direct_interc_73_
  (
    .in(grid_clb_80_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_73_out[0])
  );


  direct_interc
  direct_interc_74_
  (
    .in(grid_clb_81_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_74_out[0])
  );


  direct_interc
  direct_interc_75_
  (
    .in(grid_clb_82_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_75_out[0])
  );


  direct_interc
  direct_interc_76_
  (
    .in(grid_clb_83_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_76_out[0])
  );


  direct_interc
  direct_interc_77_
  (
    .in(grid_clb_85_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_77_out[0])
  );


  direct_interc
  direct_interc_78_
  (
    .in(grid_clb_86_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_78_out[0])
  );


  direct_interc
  direct_interc_79_
  (
    .in(grid_clb_87_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_79_out[0])
  );


  direct_interc
  direct_interc_80_
  (
    .in(grid_clb_88_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_80_out[0])
  );


  direct_interc
  direct_interc_81_
  (
    .in(grid_clb_89_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_81_out[0])
  );


  direct_interc
  direct_interc_82_
  (
    .in(grid_clb_90_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_82_out[0])
  );


  direct_interc
  direct_interc_83_
  (
    .in(grid_clb_91_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_83_out[0])
  );


  direct_interc
  direct_interc_84_
  (
    .in(grid_clb_92_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_84_out[0])
  );


  direct_interc
  direct_interc_85_
  (
    .in(grid_clb_93_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_85_out[0])
  );


  direct_interc
  direct_interc_86_
  (
    .in(grid_clb_94_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_86_out[0])
  );


  direct_interc
  direct_interc_87_
  (
    .in(grid_clb_95_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_87_out[0])
  );


  direct_interc
  direct_interc_88_
  (
    .in(grid_clb_97_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_88_out[0])
  );


  direct_interc
  direct_interc_89_
  (
    .in(grid_clb_98_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_89_out[0])
  );


  direct_interc
  direct_interc_90_
  (
    .in(grid_clb_99_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_90_out[0])
  );


  direct_interc
  direct_interc_91_
  (
    .in(grid_clb_100_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_91_out[0])
  );


  direct_interc
  direct_interc_92_
  (
    .in(grid_clb_101_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_92_out[0])
  );


  direct_interc
  direct_interc_93_
  (
    .in(grid_clb_102_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_93_out[0])
  );


  direct_interc
  direct_interc_94_
  (
    .in(grid_clb_103_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_94_out[0])
  );


  direct_interc
  direct_interc_95_
  (
    .in(grid_clb_104_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_95_out[0])
  );


  direct_interc
  direct_interc_96_
  (
    .in(grid_clb_105_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_96_out[0])
  );


  direct_interc
  direct_interc_97_
  (
    .in(grid_clb_106_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_97_out[0])
  );


  direct_interc
  direct_interc_98_
  (
    .in(grid_clb_107_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_98_out[0])
  );


  direct_interc
  direct_interc_99_
  (
    .in(grid_clb_109_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_99_out[0])
  );


  direct_interc
  direct_interc_100_
  (
    .in(grid_clb_110_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_100_out[0])
  );


  direct_interc
  direct_interc_101_
  (
    .in(grid_clb_111_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_101_out[0])
  );


  direct_interc
  direct_interc_102_
  (
    .in(grid_clb_112_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_102_out[0])
  );


  direct_interc
  direct_interc_103_
  (
    .in(grid_clb_113_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_103_out[0])
  );


  direct_interc
  direct_interc_104_
  (
    .in(grid_clb_114_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_104_out[0])
  );


  direct_interc
  direct_interc_105_
  (
    .in(grid_clb_115_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_105_out[0])
  );


  direct_interc
  direct_interc_106_
  (
    .in(grid_clb_116_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_106_out[0])
  );


  direct_interc
  direct_interc_107_
  (
    .in(grid_clb_117_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_107_out[0])
  );


  direct_interc
  direct_interc_108_
  (
    .in(grid_clb_118_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_108_out[0])
  );


  direct_interc
  direct_interc_109_
  (
    .in(grid_clb_119_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_109_out[0])
  );


  direct_interc
  direct_interc_110_
  (
    .in(grid_clb_121_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_110_out[0])
  );


  direct_interc
  direct_interc_111_
  (
    .in(grid_clb_122_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_111_out[0])
  );


  direct_interc
  direct_interc_112_
  (
    .in(grid_clb_123_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_112_out[0])
  );


  direct_interc
  direct_interc_113_
  (
    .in(grid_clb_124_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_113_out[0])
  );


  direct_interc
  direct_interc_114_
  (
    .in(grid_clb_125_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_114_out[0])
  );


  direct_interc
  direct_interc_115_
  (
    .in(grid_clb_126_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_115_out[0])
  );


  direct_interc
  direct_interc_116_
  (
    .in(grid_clb_127_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_116_out[0])
  );


  direct_interc
  direct_interc_117_
  (
    .in(grid_clb_128_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_117_out[0])
  );


  direct_interc
  direct_interc_118_
  (
    .in(grid_clb_129_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_118_out[0])
  );


  direct_interc
  direct_interc_119_
  (
    .in(grid_clb_130_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_119_out[0])
  );


  direct_interc
  direct_interc_120_
  (
    .in(grid_clb_131_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_120_out[0])
  );


  direct_interc
  direct_interc_121_
  (
    .in(grid_clb_133_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_121_out[0])
  );


  direct_interc
  direct_interc_122_
  (
    .in(grid_clb_134_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_122_out[0])
  );


  direct_interc
  direct_interc_123_
  (
    .in(grid_clb_135_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_123_out[0])
  );


  direct_interc
  direct_interc_124_
  (
    .in(grid_clb_136_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_124_out[0])
  );


  direct_interc
  direct_interc_125_
  (
    .in(grid_clb_137_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_125_out[0])
  );


  direct_interc
  direct_interc_126_
  (
    .in(grid_clb_138_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_126_out[0])
  );


  direct_interc
  direct_interc_127_
  (
    .in(grid_clb_139_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_127_out[0])
  );


  direct_interc
  direct_interc_128_
  (
    .in(grid_clb_140_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_128_out[0])
  );


  direct_interc
  direct_interc_129_
  (
    .in(grid_clb_141_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_129_out[0])
  );


  direct_interc
  direct_interc_130_
  (
    .in(grid_clb_142_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_130_out[0])
  );


  direct_interc
  direct_interc_131_
  (
    .in(grid_clb_143_bottom_width_0_height_0__pin_54_[0]),
    .out(direct_interc_131_out[0])
  );


  direct_interc
  direct_interc_132_
  (
    .in(grid_clb_1_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_132_out[0])
  );


  direct_interc
  direct_interc_133_
  (
    .in(grid_clb_2_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_133_out[0])
  );


  direct_interc
  direct_interc_134_
  (
    .in(grid_clb_3_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_134_out[0])
  );


  direct_interc
  direct_interc_135_
  (
    .in(grid_clb_4_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_135_out[0])
  );


  direct_interc
  direct_interc_136_
  (
    .in(grid_clb_5_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_136_out[0])
  );


  direct_interc
  direct_interc_137_
  (
    .in(grid_clb_6_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_137_out[0])
  );


  direct_interc
  direct_interc_138_
  (
    .in(grid_clb_7_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_138_out[0])
  );


  direct_interc
  direct_interc_139_
  (
    .in(grid_clb_8_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_139_out[0])
  );


  direct_interc
  direct_interc_140_
  (
    .in(grid_clb_9_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_140_out[0])
  );


  direct_interc
  direct_interc_141_
  (
    .in(grid_clb_10_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_141_out[0])
  );


  direct_interc
  direct_interc_142_
  (
    .in(grid_clb_11_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_142_out[0])
  );


  direct_interc
  direct_interc_143_
  (
    .in(grid_clb_13_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_143_out[0])
  );


  direct_interc
  direct_interc_144_
  (
    .in(grid_clb_14_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_144_out[0])
  );


  direct_interc
  direct_interc_145_
  (
    .in(grid_clb_15_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_145_out[0])
  );


  direct_interc
  direct_interc_146_
  (
    .in(grid_clb_16_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_146_out[0])
  );


  direct_interc
  direct_interc_147_
  (
    .in(grid_clb_17_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_147_out[0])
  );


  direct_interc
  direct_interc_148_
  (
    .in(grid_clb_18_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_148_out[0])
  );


  direct_interc
  direct_interc_149_
  (
    .in(grid_clb_19_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_149_out[0])
  );


  direct_interc
  direct_interc_150_
  (
    .in(grid_clb_20_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_150_out[0])
  );


  direct_interc
  direct_interc_151_
  (
    .in(grid_clb_21_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_151_out[0])
  );


  direct_interc
  direct_interc_152_
  (
    .in(grid_clb_22_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_152_out[0])
  );


  direct_interc
  direct_interc_153_
  (
    .in(grid_clb_23_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_153_out[0])
  );


  direct_interc
  direct_interc_154_
  (
    .in(grid_clb_25_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_154_out[0])
  );


  direct_interc
  direct_interc_155_
  (
    .in(grid_clb_26_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_155_out[0])
  );


  direct_interc
  direct_interc_156_
  (
    .in(grid_clb_27_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_156_out[0])
  );


  direct_interc
  direct_interc_157_
  (
    .in(grid_clb_28_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_157_out[0])
  );


  direct_interc
  direct_interc_158_
  (
    .in(grid_clb_29_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_158_out[0])
  );


  direct_interc
  direct_interc_159_
  (
    .in(grid_clb_30_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_159_out[0])
  );


  direct_interc
  direct_interc_160_
  (
    .in(grid_clb_31_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_160_out[0])
  );


  direct_interc
  direct_interc_161_
  (
    .in(grid_clb_32_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_161_out[0])
  );


  direct_interc
  direct_interc_162_
  (
    .in(grid_clb_33_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_162_out[0])
  );


  direct_interc
  direct_interc_163_
  (
    .in(grid_clb_34_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_163_out[0])
  );


  direct_interc
  direct_interc_164_
  (
    .in(grid_clb_35_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_164_out[0])
  );


  direct_interc
  direct_interc_165_
  (
    .in(grid_clb_37_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_165_out[0])
  );


  direct_interc
  direct_interc_166_
  (
    .in(grid_clb_38_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_166_out[0])
  );


  direct_interc
  direct_interc_167_
  (
    .in(grid_clb_39_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_167_out[0])
  );


  direct_interc
  direct_interc_168_
  (
    .in(grid_clb_40_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_168_out[0])
  );


  direct_interc
  direct_interc_169_
  (
    .in(grid_clb_41_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_169_out[0])
  );


  direct_interc
  direct_interc_170_
  (
    .in(grid_clb_42_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_170_out[0])
  );


  direct_interc
  direct_interc_171_
  (
    .in(grid_clb_43_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_171_out[0])
  );


  direct_interc
  direct_interc_172_
  (
    .in(grid_clb_44_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_172_out[0])
  );


  direct_interc
  direct_interc_173_
  (
    .in(grid_clb_45_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_173_out[0])
  );


  direct_interc
  direct_interc_174_
  (
    .in(grid_clb_46_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_174_out[0])
  );


  direct_interc
  direct_interc_175_
  (
    .in(grid_clb_47_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_175_out[0])
  );


  direct_interc
  direct_interc_176_
  (
    .in(grid_clb_49_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_176_out[0])
  );


  direct_interc
  direct_interc_177_
  (
    .in(grid_clb_50_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_177_out[0])
  );


  direct_interc
  direct_interc_178_
  (
    .in(grid_clb_51_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_178_out[0])
  );


  direct_interc
  direct_interc_179_
  (
    .in(grid_clb_52_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_179_out[0])
  );


  direct_interc
  direct_interc_180_
  (
    .in(grid_clb_53_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_180_out[0])
  );


  direct_interc
  direct_interc_181_
  (
    .in(grid_clb_54_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_181_out[0])
  );


  direct_interc
  direct_interc_182_
  (
    .in(grid_clb_55_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_182_out[0])
  );


  direct_interc
  direct_interc_183_
  (
    .in(grid_clb_56_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_183_out[0])
  );


  direct_interc
  direct_interc_184_
  (
    .in(grid_clb_57_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_184_out[0])
  );


  direct_interc
  direct_interc_185_
  (
    .in(grid_clb_58_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_185_out[0])
  );


  direct_interc
  direct_interc_186_
  (
    .in(grid_clb_59_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_186_out[0])
  );


  direct_interc
  direct_interc_187_
  (
    .in(grid_clb_61_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_187_out[0])
  );


  direct_interc
  direct_interc_188_
  (
    .in(grid_clb_62_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_188_out[0])
  );


  direct_interc
  direct_interc_189_
  (
    .in(grid_clb_63_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_189_out[0])
  );


  direct_interc
  direct_interc_190_
  (
    .in(grid_clb_64_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_190_out[0])
  );


  direct_interc
  direct_interc_191_
  (
    .in(grid_clb_65_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_191_out[0])
  );


  direct_interc
  direct_interc_192_
  (
    .in(grid_clb_66_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_192_out[0])
  );


  direct_interc
  direct_interc_193_
  (
    .in(grid_clb_67_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_193_out[0])
  );


  direct_interc
  direct_interc_194_
  (
    .in(grid_clb_68_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_194_out[0])
  );


  direct_interc
  direct_interc_195_
  (
    .in(grid_clb_69_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_195_out[0])
  );


  direct_interc
  direct_interc_196_
  (
    .in(grid_clb_70_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_196_out[0])
  );


  direct_interc
  direct_interc_197_
  (
    .in(grid_clb_71_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_197_out[0])
  );


  direct_interc
  direct_interc_198_
  (
    .in(grid_clb_73_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_198_out[0])
  );


  direct_interc
  direct_interc_199_
  (
    .in(grid_clb_74_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_199_out[0])
  );


  direct_interc
  direct_interc_200_
  (
    .in(grid_clb_75_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_200_out[0])
  );


  direct_interc
  direct_interc_201_
  (
    .in(grid_clb_76_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_201_out[0])
  );


  direct_interc
  direct_interc_202_
  (
    .in(grid_clb_77_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_202_out[0])
  );


  direct_interc
  direct_interc_203_
  (
    .in(grid_clb_78_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_203_out[0])
  );


  direct_interc
  direct_interc_204_
  (
    .in(grid_clb_79_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_204_out[0])
  );


  direct_interc
  direct_interc_205_
  (
    .in(grid_clb_80_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_205_out[0])
  );


  direct_interc
  direct_interc_206_
  (
    .in(grid_clb_81_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_206_out[0])
  );


  direct_interc
  direct_interc_207_
  (
    .in(grid_clb_82_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_207_out[0])
  );


  direct_interc
  direct_interc_208_
  (
    .in(grid_clb_83_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_208_out[0])
  );


  direct_interc
  direct_interc_209_
  (
    .in(grid_clb_85_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_209_out[0])
  );


  direct_interc
  direct_interc_210_
  (
    .in(grid_clb_86_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_210_out[0])
  );


  direct_interc
  direct_interc_211_
  (
    .in(grid_clb_87_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_211_out[0])
  );


  direct_interc
  direct_interc_212_
  (
    .in(grid_clb_88_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_212_out[0])
  );


  direct_interc
  direct_interc_213_
  (
    .in(grid_clb_89_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_213_out[0])
  );


  direct_interc
  direct_interc_214_
  (
    .in(grid_clb_90_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_214_out[0])
  );


  direct_interc
  direct_interc_215_
  (
    .in(grid_clb_91_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_215_out[0])
  );


  direct_interc
  direct_interc_216_
  (
    .in(grid_clb_92_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_216_out[0])
  );


  direct_interc
  direct_interc_217_
  (
    .in(grid_clb_93_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_217_out[0])
  );


  direct_interc
  direct_interc_218_
  (
    .in(grid_clb_94_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_218_out[0])
  );


  direct_interc
  direct_interc_219_
  (
    .in(grid_clb_95_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_219_out[0])
  );


  direct_interc
  direct_interc_220_
  (
    .in(grid_clb_97_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_220_out[0])
  );


  direct_interc
  direct_interc_221_
  (
    .in(grid_clb_98_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_221_out[0])
  );


  direct_interc
  direct_interc_222_
  (
    .in(grid_clb_99_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_222_out[0])
  );


  direct_interc
  direct_interc_223_
  (
    .in(grid_clb_100_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_223_out[0])
  );


  direct_interc
  direct_interc_224_
  (
    .in(grid_clb_101_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_224_out[0])
  );


  direct_interc
  direct_interc_225_
  (
    .in(grid_clb_102_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_225_out[0])
  );


  direct_interc
  direct_interc_226_
  (
    .in(grid_clb_103_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_226_out[0])
  );


  direct_interc
  direct_interc_227_
  (
    .in(grid_clb_104_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_227_out[0])
  );


  direct_interc
  direct_interc_228_
  (
    .in(grid_clb_105_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_228_out[0])
  );


  direct_interc
  direct_interc_229_
  (
    .in(grid_clb_106_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_229_out[0])
  );


  direct_interc
  direct_interc_230_
  (
    .in(grid_clb_107_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_230_out[0])
  );


  direct_interc
  direct_interc_231_
  (
    .in(grid_clb_109_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_231_out[0])
  );


  direct_interc
  direct_interc_232_
  (
    .in(grid_clb_110_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_232_out[0])
  );


  direct_interc
  direct_interc_233_
  (
    .in(grid_clb_111_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_233_out[0])
  );


  direct_interc
  direct_interc_234_
  (
    .in(grid_clb_112_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_234_out[0])
  );


  direct_interc
  direct_interc_235_
  (
    .in(grid_clb_113_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_235_out[0])
  );


  direct_interc
  direct_interc_236_
  (
    .in(grid_clb_114_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_236_out[0])
  );


  direct_interc
  direct_interc_237_
  (
    .in(grid_clb_115_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_237_out[0])
  );


  direct_interc
  direct_interc_238_
  (
    .in(grid_clb_116_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_238_out[0])
  );


  direct_interc
  direct_interc_239_
  (
    .in(grid_clb_117_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_239_out[0])
  );


  direct_interc
  direct_interc_240_
  (
    .in(grid_clb_118_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_240_out[0])
  );


  direct_interc
  direct_interc_241_
  (
    .in(grid_clb_119_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_241_out[0])
  );


  direct_interc
  direct_interc_242_
  (
    .in(grid_clb_121_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_242_out[0])
  );


  direct_interc
  direct_interc_243_
  (
    .in(grid_clb_122_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_243_out[0])
  );


  direct_interc
  direct_interc_244_
  (
    .in(grid_clb_123_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_244_out[0])
  );


  direct_interc
  direct_interc_245_
  (
    .in(grid_clb_124_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_245_out[0])
  );


  direct_interc
  direct_interc_246_
  (
    .in(grid_clb_125_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_246_out[0])
  );


  direct_interc
  direct_interc_247_
  (
    .in(grid_clb_126_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_247_out[0])
  );


  direct_interc
  direct_interc_248_
  (
    .in(grid_clb_127_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_248_out[0])
  );


  direct_interc
  direct_interc_249_
  (
    .in(grid_clb_128_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_249_out[0])
  );


  direct_interc
  direct_interc_250_
  (
    .in(grid_clb_129_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_250_out[0])
  );


  direct_interc
  direct_interc_251_
  (
    .in(grid_clb_130_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_251_out[0])
  );


  direct_interc
  direct_interc_252_
  (
    .in(grid_clb_131_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_252_out[0])
  );


  direct_interc
  direct_interc_253_
  (
    .in(grid_clb_133_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_253_out[0])
  );


  direct_interc
  direct_interc_254_
  (
    .in(grid_clb_134_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_254_out[0])
  );


  direct_interc
  direct_interc_255_
  (
    .in(grid_clb_135_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_255_out[0])
  );


  direct_interc
  direct_interc_256_
  (
    .in(grid_clb_136_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_256_out[0])
  );


  direct_interc
  direct_interc_257_
  (
    .in(grid_clb_137_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_257_out[0])
  );


  direct_interc
  direct_interc_258_
  (
    .in(grid_clb_138_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_258_out[0])
  );


  direct_interc
  direct_interc_259_
  (
    .in(grid_clb_139_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_259_out[0])
  );


  direct_interc
  direct_interc_260_
  (
    .in(grid_clb_140_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_260_out[0])
  );


  direct_interc
  direct_interc_261_
  (
    .in(grid_clb_141_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_261_out[0])
  );


  direct_interc
  direct_interc_262_
  (
    .in(grid_clb_142_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_262_out[0])
  );


  direct_interc
  direct_interc_263_
  (
    .in(grid_clb_143_bottom_width_0_height_0__pin_52_[0]),
    .out(direct_interc_263_out[0])
  );


  direct_interc
  direct_interc_264_
  (
    .in(grid_clb_1_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_264_out[0])
  );


  direct_interc
  direct_interc_265_
  (
    .in(grid_clb_2_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_265_out[0])
  );


  direct_interc
  direct_interc_266_
  (
    .in(grid_clb_3_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_266_out[0])
  );


  direct_interc
  direct_interc_267_
  (
    .in(grid_clb_4_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_267_out[0])
  );


  direct_interc
  direct_interc_268_
  (
    .in(grid_clb_5_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_268_out[0])
  );


  direct_interc
  direct_interc_269_
  (
    .in(grid_clb_6_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_269_out[0])
  );


  direct_interc
  direct_interc_270_
  (
    .in(grid_clb_7_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_270_out[0])
  );


  direct_interc
  direct_interc_271_
  (
    .in(grid_clb_8_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_271_out[0])
  );


  direct_interc
  direct_interc_272_
  (
    .in(grid_clb_9_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_272_out[0])
  );


  direct_interc
  direct_interc_273_
  (
    .in(grid_clb_10_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_273_out[0])
  );


  direct_interc
  direct_interc_274_
  (
    .in(grid_clb_11_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_274_out[0])
  );


  direct_interc
  direct_interc_275_
  (
    .in(grid_clb_13_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_275_out[0])
  );


  direct_interc
  direct_interc_276_
  (
    .in(grid_clb_14_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_276_out[0])
  );


  direct_interc
  direct_interc_277_
  (
    .in(grid_clb_15_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_277_out[0])
  );


  direct_interc
  direct_interc_278_
  (
    .in(grid_clb_16_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_278_out[0])
  );


  direct_interc
  direct_interc_279_
  (
    .in(grid_clb_17_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_279_out[0])
  );


  direct_interc
  direct_interc_280_
  (
    .in(grid_clb_18_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_280_out[0])
  );


  direct_interc
  direct_interc_281_
  (
    .in(grid_clb_19_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_281_out[0])
  );


  direct_interc
  direct_interc_282_
  (
    .in(grid_clb_20_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_282_out[0])
  );


  direct_interc
  direct_interc_283_
  (
    .in(grid_clb_21_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_283_out[0])
  );


  direct_interc
  direct_interc_284_
  (
    .in(grid_clb_22_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_284_out[0])
  );


  direct_interc
  direct_interc_285_
  (
    .in(grid_clb_23_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_285_out[0])
  );


  direct_interc
  direct_interc_286_
  (
    .in(grid_clb_25_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_286_out[0])
  );


  direct_interc
  direct_interc_287_
  (
    .in(grid_clb_26_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_287_out[0])
  );


  direct_interc
  direct_interc_288_
  (
    .in(grid_clb_27_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_288_out[0])
  );


  direct_interc
  direct_interc_289_
  (
    .in(grid_clb_28_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_289_out[0])
  );


  direct_interc
  direct_interc_290_
  (
    .in(grid_clb_29_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_290_out[0])
  );


  direct_interc
  direct_interc_291_
  (
    .in(grid_clb_30_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_291_out[0])
  );


  direct_interc
  direct_interc_292_
  (
    .in(grid_clb_31_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_292_out[0])
  );


  direct_interc
  direct_interc_293_
  (
    .in(grid_clb_32_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_293_out[0])
  );


  direct_interc
  direct_interc_294_
  (
    .in(grid_clb_33_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_294_out[0])
  );


  direct_interc
  direct_interc_295_
  (
    .in(grid_clb_34_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_295_out[0])
  );


  direct_interc
  direct_interc_296_
  (
    .in(grid_clb_35_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_296_out[0])
  );


  direct_interc
  direct_interc_297_
  (
    .in(grid_clb_37_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_297_out[0])
  );


  direct_interc
  direct_interc_298_
  (
    .in(grid_clb_38_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_298_out[0])
  );


  direct_interc
  direct_interc_299_
  (
    .in(grid_clb_39_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_299_out[0])
  );


  direct_interc
  direct_interc_300_
  (
    .in(grid_clb_40_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_300_out[0])
  );


  direct_interc
  direct_interc_301_
  (
    .in(grid_clb_41_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_301_out[0])
  );


  direct_interc
  direct_interc_302_
  (
    .in(grid_clb_42_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_302_out[0])
  );


  direct_interc
  direct_interc_303_
  (
    .in(grid_clb_43_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_303_out[0])
  );


  direct_interc
  direct_interc_304_
  (
    .in(grid_clb_44_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_304_out[0])
  );


  direct_interc
  direct_interc_305_
  (
    .in(grid_clb_45_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_305_out[0])
  );


  direct_interc
  direct_interc_306_
  (
    .in(grid_clb_46_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_306_out[0])
  );


  direct_interc
  direct_interc_307_
  (
    .in(grid_clb_47_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_307_out[0])
  );


  direct_interc
  direct_interc_308_
  (
    .in(grid_clb_49_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_308_out[0])
  );


  direct_interc
  direct_interc_309_
  (
    .in(grid_clb_50_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_309_out[0])
  );


  direct_interc
  direct_interc_310_
  (
    .in(grid_clb_51_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_310_out[0])
  );


  direct_interc
  direct_interc_311_
  (
    .in(grid_clb_52_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_311_out[0])
  );


  direct_interc
  direct_interc_312_
  (
    .in(grid_clb_53_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_312_out[0])
  );


  direct_interc
  direct_interc_313_
  (
    .in(grid_clb_54_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_313_out[0])
  );


  direct_interc
  direct_interc_314_
  (
    .in(grid_clb_55_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_314_out[0])
  );


  direct_interc
  direct_interc_315_
  (
    .in(grid_clb_56_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_315_out[0])
  );


  direct_interc
  direct_interc_316_
  (
    .in(grid_clb_57_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_316_out[0])
  );


  direct_interc
  direct_interc_317_
  (
    .in(grid_clb_58_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_317_out[0])
  );


  direct_interc
  direct_interc_318_
  (
    .in(grid_clb_59_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_318_out[0])
  );


  direct_interc
  direct_interc_319_
  (
    .in(grid_clb_61_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_319_out[0])
  );


  direct_interc
  direct_interc_320_
  (
    .in(grid_clb_62_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_320_out[0])
  );


  direct_interc
  direct_interc_321_
  (
    .in(grid_clb_63_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_321_out[0])
  );


  direct_interc
  direct_interc_322_
  (
    .in(grid_clb_64_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_322_out[0])
  );


  direct_interc
  direct_interc_323_
  (
    .in(grid_clb_65_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_323_out[0])
  );


  direct_interc
  direct_interc_324_
  (
    .in(grid_clb_66_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_324_out[0])
  );


  direct_interc
  direct_interc_325_
  (
    .in(grid_clb_67_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_325_out[0])
  );


  direct_interc
  direct_interc_326_
  (
    .in(grid_clb_68_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_326_out[0])
  );


  direct_interc
  direct_interc_327_
  (
    .in(grid_clb_69_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_327_out[0])
  );


  direct_interc
  direct_interc_328_
  (
    .in(grid_clb_70_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_328_out[0])
  );


  direct_interc
  direct_interc_329_
  (
    .in(grid_clb_71_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_329_out[0])
  );


  direct_interc
  direct_interc_330_
  (
    .in(grid_clb_73_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_330_out[0])
  );


  direct_interc
  direct_interc_331_
  (
    .in(grid_clb_74_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_331_out[0])
  );


  direct_interc
  direct_interc_332_
  (
    .in(grid_clb_75_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_332_out[0])
  );


  direct_interc
  direct_interc_333_
  (
    .in(grid_clb_76_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_333_out[0])
  );


  direct_interc
  direct_interc_334_
  (
    .in(grid_clb_77_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_334_out[0])
  );


  direct_interc
  direct_interc_335_
  (
    .in(grid_clb_78_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_335_out[0])
  );


  direct_interc
  direct_interc_336_
  (
    .in(grid_clb_79_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_336_out[0])
  );


  direct_interc
  direct_interc_337_
  (
    .in(grid_clb_80_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_337_out[0])
  );


  direct_interc
  direct_interc_338_
  (
    .in(grid_clb_81_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_338_out[0])
  );


  direct_interc
  direct_interc_339_
  (
    .in(grid_clb_82_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_339_out[0])
  );


  direct_interc
  direct_interc_340_
  (
    .in(grid_clb_83_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_340_out[0])
  );


  direct_interc
  direct_interc_341_
  (
    .in(grid_clb_85_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_341_out[0])
  );


  direct_interc
  direct_interc_342_
  (
    .in(grid_clb_86_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_342_out[0])
  );


  direct_interc
  direct_interc_343_
  (
    .in(grid_clb_87_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_343_out[0])
  );


  direct_interc
  direct_interc_344_
  (
    .in(grid_clb_88_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_344_out[0])
  );


  direct_interc
  direct_interc_345_
  (
    .in(grid_clb_89_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_345_out[0])
  );


  direct_interc
  direct_interc_346_
  (
    .in(grid_clb_90_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_346_out[0])
  );


  direct_interc
  direct_interc_347_
  (
    .in(grid_clb_91_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_347_out[0])
  );


  direct_interc
  direct_interc_348_
  (
    .in(grid_clb_92_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_348_out[0])
  );


  direct_interc
  direct_interc_349_
  (
    .in(grid_clb_93_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_349_out[0])
  );


  direct_interc
  direct_interc_350_
  (
    .in(grid_clb_94_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_350_out[0])
  );


  direct_interc
  direct_interc_351_
  (
    .in(grid_clb_95_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_351_out[0])
  );


  direct_interc
  direct_interc_352_
  (
    .in(grid_clb_97_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_352_out[0])
  );


  direct_interc
  direct_interc_353_
  (
    .in(grid_clb_98_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_353_out[0])
  );


  direct_interc
  direct_interc_354_
  (
    .in(grid_clb_99_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_354_out[0])
  );


  direct_interc
  direct_interc_355_
  (
    .in(grid_clb_100_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_355_out[0])
  );


  direct_interc
  direct_interc_356_
  (
    .in(grid_clb_101_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_356_out[0])
  );


  direct_interc
  direct_interc_357_
  (
    .in(grid_clb_102_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_357_out[0])
  );


  direct_interc
  direct_interc_358_
  (
    .in(grid_clb_103_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_358_out[0])
  );


  direct_interc
  direct_interc_359_
  (
    .in(grid_clb_104_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_359_out[0])
  );


  direct_interc
  direct_interc_360_
  (
    .in(grid_clb_105_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_360_out[0])
  );


  direct_interc
  direct_interc_361_
  (
    .in(grid_clb_106_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_361_out[0])
  );


  direct_interc
  direct_interc_362_
  (
    .in(grid_clb_107_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_362_out[0])
  );


  direct_interc
  direct_interc_363_
  (
    .in(grid_clb_109_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_363_out[0])
  );


  direct_interc
  direct_interc_364_
  (
    .in(grid_clb_110_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_364_out[0])
  );


  direct_interc
  direct_interc_365_
  (
    .in(grid_clb_111_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_365_out[0])
  );


  direct_interc
  direct_interc_366_
  (
    .in(grid_clb_112_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_366_out[0])
  );


  direct_interc
  direct_interc_367_
  (
    .in(grid_clb_113_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_367_out[0])
  );


  direct_interc
  direct_interc_368_
  (
    .in(grid_clb_114_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_368_out[0])
  );


  direct_interc
  direct_interc_369_
  (
    .in(grid_clb_115_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_369_out[0])
  );


  direct_interc
  direct_interc_370_
  (
    .in(grid_clb_116_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_370_out[0])
  );


  direct_interc
  direct_interc_371_
  (
    .in(grid_clb_117_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_371_out[0])
  );


  direct_interc
  direct_interc_372_
  (
    .in(grid_clb_118_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_372_out[0])
  );


  direct_interc
  direct_interc_373_
  (
    .in(grid_clb_119_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_373_out[0])
  );


  direct_interc
  direct_interc_374_
  (
    .in(grid_clb_121_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_374_out[0])
  );


  direct_interc
  direct_interc_375_
  (
    .in(grid_clb_122_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_375_out[0])
  );


  direct_interc
  direct_interc_376_
  (
    .in(grid_clb_123_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_376_out[0])
  );


  direct_interc
  direct_interc_377_
  (
    .in(grid_clb_124_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_377_out[0])
  );


  direct_interc
  direct_interc_378_
  (
    .in(grid_clb_125_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_378_out[0])
  );


  direct_interc
  direct_interc_379_
  (
    .in(grid_clb_126_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_379_out[0])
  );


  direct_interc
  direct_interc_380_
  (
    .in(grid_clb_127_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_380_out[0])
  );


  direct_interc
  direct_interc_381_
  (
    .in(grid_clb_128_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_381_out[0])
  );


  direct_interc
  direct_interc_382_
  (
    .in(grid_clb_129_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_382_out[0])
  );


  direct_interc
  direct_interc_383_
  (
    .in(grid_clb_130_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_383_out[0])
  );


  direct_interc
  direct_interc_384_
  (
    .in(grid_clb_131_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_384_out[0])
  );


  direct_interc
  direct_interc_385_
  (
    .in(grid_clb_133_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_385_out[0])
  );


  direct_interc
  direct_interc_386_
  (
    .in(grid_clb_134_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_386_out[0])
  );


  direct_interc
  direct_interc_387_
  (
    .in(grid_clb_135_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_387_out[0])
  );


  direct_interc
  direct_interc_388_
  (
    .in(grid_clb_136_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_388_out[0])
  );


  direct_interc
  direct_interc_389_
  (
    .in(grid_clb_137_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_389_out[0])
  );


  direct_interc
  direct_interc_390_
  (
    .in(grid_clb_138_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_390_out[0])
  );


  direct_interc
  direct_interc_391_
  (
    .in(grid_clb_139_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_391_out[0])
  );


  direct_interc
  direct_interc_392_
  (
    .in(grid_clb_140_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_392_out[0])
  );


  direct_interc
  direct_interc_393_
  (
    .in(grid_clb_141_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_393_out[0])
  );


  direct_interc
  direct_interc_394_
  (
    .in(grid_clb_142_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_394_out[0])
  );


  direct_interc
  direct_interc_395_
  (
    .in(grid_clb_143_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_395_out[0])
  );


  direct_interc
  direct_interc_396_
  (
    .in(grid_clb_0_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_396_out[0])
  );


  direct_interc
  direct_interc_397_
  (
    .in(grid_clb_12_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_397_out[0])
  );


  direct_interc
  direct_interc_398_
  (
    .in(grid_clb_24_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_398_out[0])
  );


  direct_interc
  direct_interc_399_
  (
    .in(grid_clb_36_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_399_out[0])
  );


  direct_interc
  direct_interc_400_
  (
    .in(grid_clb_48_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_400_out[0])
  );


  direct_interc
  direct_interc_401_
  (
    .in(grid_clb_60_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_401_out[0])
  );


  direct_interc
  direct_interc_402_
  (
    .in(grid_clb_72_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_402_out[0])
  );


  direct_interc
  direct_interc_403_
  (
    .in(grid_clb_84_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_403_out[0])
  );


  direct_interc
  direct_interc_404_
  (
    .in(grid_clb_96_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_404_out[0])
  );


  direct_interc
  direct_interc_405_
  (
    .in(grid_clb_108_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_405_out[0])
  );


  direct_interc
  direct_interc_406_
  (
    .in(grid_clb_120_bottom_width_0_height_0__pin_53_[0]),
    .out(direct_interc_406_out[0])
  );


endmodule

