VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO cby_2__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 73.6 BY 87.04 ;
  SYMMETRY X Y ;
  PIN pReset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 44.3 0.595 44.44 ;
    END
  END pReset[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5 0 59.64 0.485 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.98 0 54.12 0.485 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.14 0 52.28 0.485 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.66 0 57.8 0.485 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.4 0 20.54 0.485 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.98 0 31.12 0.485 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.74 0 56.88 0.485 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.46 0 25.6 0.485 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.54 0 24.68 0.485 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.76 0 27.9 0.485 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.16 0 23.3 0.485 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.94 0 43.08 0.485 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.66 0 34.8 0.485 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.4 0 66.54 0.485 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.38 0 49.52 0.485 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.62 0 46.76 0.485 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.24 0 22.38 0.485 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.86 0 44 0.485 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.9 0 32.04 0.485 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.96 0 37.1 0.485 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.72 0 39.86 0.485 ;
    END
  END chany_bottom_in[20]
  PIN chany_bottom_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.68 0 28.82 0.485 ;
    END
  END chany_bottom_in[21]
  PIN chany_bottom_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.5 0 13.64 0.485 ;
    END
  END chany_bottom_in[22]
  PIN chany_bottom_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.02 0 42.16 0.485 ;
    END
  END chany_bottom_in[23]
  PIN chany_bottom_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.64 0 40.78 0.485 ;
    END
  END chany_bottom_in[24]
  PIN chany_bottom_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.06 0 30.2 0.485 ;
    END
  END chany_bottom_in[25]
  PIN chany_bottom_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.7 0 45.84 0.485 ;
    END
  END chany_bottom_in[26]
  PIN chany_bottom_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.32 0 21.46 0.485 ;
    END
  END chany_bottom_in[27]
  PIN chany_bottom_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.78 0 44.92 0.485 ;
    END
  END chany_bottom_in[28]
  PIN chany_bottom_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.64 0 63.78 0.485 ;
    END
  END chany_bottom_in[29]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.6 86.555 6.74 87.04 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.68 86.555 5.82 87.04 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.76 86.555 4.9 87.04 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.74 86.555 10.88 87.04 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.32 86.555 21.46 87.04 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.82 86.555 9.96 87.04 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.98 86.555 54.12 87.04 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.4 86.555 20.54 87.04 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.9 86.555 55.04 87.04 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.42 86.555 37.56 87.04 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.46 86.555 48.6 87.04 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.62 86.555 46.76 87.04 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.48 86.555 19.62 87.04 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.3 86.555 50.44 87.04 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.14 86.555 52.28 87.04 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.86 86.555 44 87.04 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.24 86.555 22.38 87.04 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.7 86.555 45.84 87.04 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.16 86.555 23.3 87.04 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.06 86.555 53.2 87.04 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 86.555 35.72 87.04 ;
    END
  END chany_top_in[20]
  PIN chany_top_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5 86.555 59.64 87.04 ;
    END
  END chany_top_in[21]
  PIN chany_top_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.5 86.555 36.64 87.04 ;
    END
  END chany_top_in[22]
  PIN chany_top_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.2 86.555 34.34 87.04 ;
    END
  END chany_top_in[23]
  PIN chany_top_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.28 86.555 33.42 87.04 ;
    END
  END chany_top_in[24]
  PIN chany_top_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.64 86.555 17.78 87.04 ;
    END
  END chany_top_in[25]
  PIN chany_top_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.38 86.555 49.52 87.04 ;
    END
  END chany_top_in[26]
  PIN chany_top_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.08 86.555 24.22 87.04 ;
    END
  END chany_top_in[27]
  PIN chany_top_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.78 86.555 44.92 87.04 ;
    END
  END chany_top_in[28]
  PIN chany_top_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 86.555 64.24 87.04 ;
    END
  END chany_top_in[29]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 75.24 0.595 75.38 ;
    END
  END ccff_head[0]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.56 0 64.7 0.485 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.67 0 30.97 0.8 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.28 0 10.42 0.485 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.48 0 65.62 0.485 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.56 0 18.7 0.485 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 32.51 0 32.81 0.8 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.24 0 68.38 0.485 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.74 0 33.88 0.485 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.8 0 38.94 0.485 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 0 62.4 0.485 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.48 0 19.62 0.485 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.82 0 32.96 0.485 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.46 0 48.6 0.485 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.06 0 53.2 0.485 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.88 0 38.02 0.485 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.54 0 47.68 0.485 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.3 0 50.44 0.485 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.16 0 69.3 0.485 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.9 0 55.04 0.485 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.04 0 36.18 0.485 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.64 0 17.78 0.485 ;
    END
  END chany_bottom_out[20]
  PIN chany_bottom_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.38 0 26.52 0.485 ;
    END
  END chany_bottom_out[21]
  PIN chany_bottom_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.52 0 7.66 0.485 ;
    END
  END chany_bottom_out[22]
  PIN chany_bottom_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.2 0 11.34 0.485 ;
    END
  END chany_bottom_out[23]
  PIN chany_bottom_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.32 0 67.46 0.485 ;
    END
  END chany_bottom_out[24]
  PIN chany_bottom_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.22 0 51.36 0.485 ;
    END
  END chany_bottom_out[25]
  PIN chany_bottom_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71 0 71.14 0.485 ;
    END
  END chany_bottom_out[26]
  PIN chany_bottom_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.71 0 42.01 0.8 ;
    END
  END chany_bottom_out[27]
  PIN chany_bottom_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 0 61.48 0.485 ;
    END
  END chany_bottom_out[28]
  PIN chany_bottom_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.08 0 70.22 0.485 ;
    END
  END chany_bottom_out[29]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 32.51 86.24 32.81 87.04 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.67 86.24 30.97 87.04 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 34.35 86.24 34.65 87.04 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.88 86.555 15.02 87.04 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 86.555 39.4 87.04 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.94 86.555 66.08 87.04 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.56 86.555 18.7 87.04 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.66 86.555 57.8 87.04 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 86.555 41.24 87.04 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.02 86.555 42.16 87.04 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.3 86.555 27.44 87.04 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.8 86.555 15.94 87.04 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.92 86.555 26.06 87.04 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.54 86.555 47.68 87.04 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.22 86.555 28.36 87.04 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 86.555 62.4 87.04 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 86.555 61.48 87.04 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 86.555 65.16 87.04 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.06 86.555 30.2 87.04 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.72 86.555 16.86 87.04 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.94 86.555 43.08 87.04 ;
    END
  END chany_top_out[20]
  PIN chany_top_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.22 86.555 51.36 87.04 ;
    END
  END chany_top_out[21]
  PIN chany_top_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.82 86.555 55.96 87.04 ;
    END
  END chany_top_out[22]
  PIN chany_top_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.18 86.555 40.32 87.04 ;
    END
  END chany_top_out[23]
  PIN chany_top_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.36 86.555 32.5 87.04 ;
    END
  END chany_top_out[24]
  PIN chany_top_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.18 86.555 63.32 87.04 ;
    END
  END chany_top_out[25]
  PIN chany_top_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.98 86.555 31.12 87.04 ;
    END
  END chany_top_out[26]
  PIN chany_top_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25 86.555 25.14 87.04 ;
    END
  END chany_top_out[27]
  PIN chany_top_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.42 86.555 60.56 87.04 ;
    END
  END chany_top_out[28]
  PIN chany_top_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.74 86.555 56.88 87.04 ;
    END
  END chany_top_out[29]
  PIN right_grid_pin_0_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 57.35 86.24 57.65 87.04 ;
    END
  END right_grid_pin_0_[0]
  PIN left_grid_pin_16_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 22.54 0.595 22.68 ;
    END
  END left_grid_pin_16_[0]
  PIN left_grid_pin_17_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 14.72 0.595 14.86 ;
    END
  END left_grid_pin_17_[0]
  PIN left_grid_pin_18_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 15.4 0.595 15.54 ;
    END
  END left_grid_pin_18_[0]
  PIN left_grid_pin_19_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 23.22 0.595 23.36 ;
    END
  END left_grid_pin_19_[0]
  PIN left_grid_pin_20_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 6.22 0.595 6.36 ;
    END
  END left_grid_pin_20_[0]
  PIN left_grid_pin_21_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 6.9 0.595 7.04 ;
    END
  END left_grid_pin_21_[0]
  PIN left_grid_pin_22_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 1.8 0.595 1.94 ;
    END
  END left_grid_pin_22_[0]
  PIN left_grid_pin_23_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 4.52 0.595 4.66 ;
    END
  END left_grid_pin_23_[0]
  PIN left_grid_pin_24_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 18.12 0.595 18.26 ;
    END
  END left_grid_pin_24_[0]
  PIN left_grid_pin_25_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 17.44 0.595 17.58 ;
    END
  END left_grid_pin_25_[0]
  PIN left_grid_pin_26_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 20.5 0.595 20.64 ;
    END
  END left_grid_pin_26_[0]
  PIN left_grid_pin_27_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 19.82 0.595 19.96 ;
    END
  END left_grid_pin_27_[0]
  PIN left_grid_pin_28_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 60.96 0.595 61.1 ;
    END
  END left_grid_pin_28_[0]
  PIN left_grid_pin_29_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 64.02 0.595 64.16 ;
    END
  END left_grid_pin_29_[0]
  PIN left_grid_pin_30_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 61.64 0.595 61.78 ;
    END
  END left_grid_pin_30_[0]
  PIN left_grid_pin_31_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 63.34 0.595 63.48 ;
    END
  END left_grid_pin_31_[0]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.82 0 55.96 0.485 ;
    END
  END ccff_tail[0]
  PIN IO_ISOL_N[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 8.94 0.595 9.08 ;
    END
  END IO_ISOL_N[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 73.005 82.72 73.6 82.86 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 73.005 83.4 73.6 83.54 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 73.005 85.1 73.6 85.24 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN left_width_0_height_0__pin_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 60.11 86.24 60.41 87.04 ;
    END
  END left_width_0_height_0__pin_0_[0]
  PIN left_width_0_height_0__pin_1_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 86.555 38.48 87.04 ;
    END
  END left_width_0_height_0__pin_1_upper[0]
  PIN left_width_0_height_0__pin_1_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.42 0 60.56 0.485 ;
    END
  END left_width_0_height_0__pin_1_lower[0]
  PIN pReset_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.6 0 6.74 0.485 ;
    END
  END pReset_S_in
  PIN prog_clk_0_W_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 0 3.84 0.595 3.98 ;
    END
  END prog_clk_0_W_in
  PIN prog_clk_0_S_out
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 2.46 0 2.6 0.485 ;
    END
  END prog_clk_0_S_out
  PIN prog_clk_0_N_out
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 11.66 86.555 11.8 87.04 ;
    END
  END prog_clk_0_N_out
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 1.12 3.2 4.32 ;
        RECT 70.4 1.12 73.6 4.32 ;
        RECT 0 41.92 3.2 45.12 ;
        RECT 70.4 41.92 73.6 45.12 ;
        RECT 0 82.72 3.2 85.92 ;
        RECT 70.4 82.72 73.6 85.92 ;
      LAYER met4 ;
        RECT 14.42 0 15.02 0.6 ;
        RECT 43.86 0 44.46 0.6 ;
        RECT 14.42 86.44 15.02 87.04 ;
        RECT 43.86 86.44 44.46 87.04 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 73.12 2.48 73.6 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 73.12 7.92 73.6 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 73.12 13.36 73.6 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 73.12 18.8 73.6 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 73.12 24.24 73.6 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 73.12 29.68 73.6 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 73.12 35.12 73.6 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 73.12 40.56 73.6 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 73.12 46 73.6 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 73.12 51.44 73.6 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 73.12 56.88 73.6 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 73.12 62.32 73.6 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 73.12 67.76 73.6 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 73.12 73.2 73.6 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 73.12 78.64 73.6 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 73.12 84.08 73.6 84.56 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 21.52 3.2 24.72 ;
        RECT 70.4 21.52 73.6 24.72 ;
        RECT 0 62.32 3.2 65.52 ;
        RECT 70.4 62.32 73.6 65.52 ;
      LAYER met4 ;
        RECT 29.14 0 29.74 0.6 ;
        RECT 58.58 0 59.18 0.6 ;
        RECT 29.14 86.44 29.74 87.04 ;
        RECT 58.58 86.44 59.18 87.04 ;
      LAYER met1 ;
        RECT 0 -0.24 0.48 0.24 ;
        RECT 73.12 -0.24 73.6 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 73.12 5.2 73.6 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 73.12 10.64 73.6 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 73.12 16.08 73.6 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 73.12 21.52 73.6 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 73.12 26.96 73.6 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 73.12 32.4 73.6 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 73.12 37.84 73.6 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 73.12 43.28 73.6 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 73.12 48.72 73.6 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 73.12 54.16 73.6 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 73.12 59.6 73.6 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 73.12 65.04 73.6 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 73.12 70.48 73.6 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 73.12 75.92 73.6 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 73.12 81.36 73.6 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 73.12 86.8 73.6 87.28 ;
    END
  END VSS
  OBS
    LAYER met1 ;
      POLYGON 72.84 87.28 72.84 86.8 59.04 86.8 59.04 86.79 58.72 86.79 58.72 86.8 29.6 86.8 29.6 86.79 29.28 86.79 29.28 86.8 0.76 86.8 0.76 87.28 ;
      POLYGON 59.04 0.25 59.04 0.24 72.84 0.24 72.84 -0.24 0.76 -0.24 0.76 0.24 29.28 0.24 29.28 0.25 29.6 0.25 29.6 0.24 58.72 0.24 58.72 0.25 ;
      POLYGON 72.84 86.76 72.84 86.52 73.32 86.52 73.32 85.52 72.725 85.52 72.725 84.82 72.84 84.82 72.84 83.82 72.725 83.82 72.725 82.44 73.32 82.44 73.32 82.12 72.84 82.12 72.84 81.08 73.32 81.08 73.32 79.4 72.84 79.4 72.84 78.36 73.32 78.36 73.32 76.68 72.84 76.68 72.84 75.64 73.32 75.64 73.32 73.96 72.84 73.96 72.84 72.92 73.32 72.92 73.32 71.24 72.84 71.24 72.84 70.2 73.32 70.2 73.32 68.52 72.84 68.52 72.84 67.48 73.32 67.48 73.32 65.8 72.84 65.8 72.84 64.76 73.32 64.76 73.32 63.08 72.84 63.08 72.84 62.04 73.32 62.04 73.32 60.36 72.84 60.36 72.84 59.32 73.32 59.32 73.32 57.64 72.84 57.64 72.84 56.6 73.32 56.6 73.32 54.92 72.84 54.92 72.84 53.88 73.32 53.88 73.32 52.2 72.84 52.2 72.84 51.16 73.32 51.16 73.32 49.48 72.84 49.48 72.84 48.44 73.32 48.44 73.32 46.76 72.84 46.76 72.84 45.72 73.32 45.72 73.32 44.04 72.84 44.04 72.84 43 73.32 43 73.32 41.32 72.84 41.32 72.84 40.28 73.32 40.28 73.32 38.6 72.84 38.6 72.84 37.56 73.32 37.56 73.32 35.88 72.84 35.88 72.84 34.84 73.32 34.84 73.32 33.16 72.84 33.16 72.84 32.12 73.32 32.12 73.32 30.44 72.84 30.44 72.84 29.4 73.32 29.4 73.32 27.72 72.84 27.72 72.84 26.68 73.32 26.68 73.32 25 72.84 25 72.84 23.96 73.32 23.96 73.32 22.28 72.84 22.28 72.84 21.24 73.32 21.24 73.32 19.56 72.84 19.56 72.84 18.52 73.32 18.52 73.32 16.84 72.84 16.84 72.84 15.8 73.32 15.8 73.32 14.12 72.84 14.12 72.84 13.08 73.32 13.08 73.32 11.4 72.84 11.4 72.84 10.36 73.32 10.36 73.32 8.68 72.84 8.68 72.84 7.64 73.32 7.64 73.32 5.96 72.84 5.96 72.84 4.92 73.32 4.92 73.32 3.24 72.84 3.24 72.84 2.2 73.32 2.2 73.32 0.52 72.84 0.52 72.84 0.28 0.76 0.28 0.76 0.52 0.28 0.52 0.28 1.52 0.875 1.52 0.875 2.22 0.76 2.22 0.76 3.24 0.28 3.24 0.28 3.56 0.875 3.56 0.875 4.94 0.76 4.94 0.76 5.94 0.875 5.94 0.875 7.32 0.28 7.32 0.28 7.64 0.76 7.64 0.76 8.66 0.875 8.66 0.875 9.36 0.28 9.36 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 14.44 0.875 14.44 0.875 15.82 0.76 15.82 0.76 16.84 0.28 16.84 0.28 17.16 0.875 17.16 0.875 18.54 0.76 18.54 0.76 19.54 0.875 19.54 0.875 20.92 0.28 20.92 0.28 21.24 0.76 21.24 0.76 22.26 0.875 22.26 0.875 23.64 0.28 23.64 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.02 0.875 44.02 0.875 44.72 0.28 44.72 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 60.68 0.875 60.68 0.875 62.06 0.76 62.06 0.76 63.06 0.875 63.06 0.875 64.44 0.28 64.44 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 74.96 0.875 74.96 0.875 75.66 0.76 75.66 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 86.76 ;
    LAYER met2 ;
      RECT 58.74 86.735 59.02 87.105 ;
      RECT 29.3 86.735 29.58 87.105 ;
      POLYGON 31.58 86.94 31.58 82.04 31.44 82.04 31.44 86.8 31.4 86.8 31.4 86.94 ;
      RECT 18.96 86.37 19.22 86.69 ;
      RECT 57.14 86.03 57.4 86.35 ;
      POLYGON 9.5 5.85 9.5 0.24 10 0.24 10 0.1 9.36 0.1 9.36 5.85 ;
      RECT 30.46 0.69 30.72 1.01 ;
      RECT 40.12 0.35 40.38 0.67 ;
      RECT 26.78 0.35 27.04 0.67 ;
      RECT 20.8 0.35 21.06 0.67 ;
      RECT 17.12 0.35 17.38 0.67 ;
      RECT 58.74 -0.065 59.02 0.305 ;
      RECT 29.3 -0.065 29.58 0.305 ;
      POLYGON 73.32 86.76 73.32 0.28 71.42 0.28 71.42 0.765 70.72 0.765 70.72 0.28 70.5 0.28 70.5 0.765 69.8 0.765 69.8 0.28 69.58 0.28 69.58 0.765 68.88 0.765 68.88 0.28 68.66 0.28 68.66 0.765 67.96 0.765 67.96 0.28 67.74 0.28 67.74 0.765 67.04 0.765 67.04 0.28 66.82 0.28 66.82 0.765 66.12 0.765 66.12 0.28 65.9 0.28 65.9 0.765 65.2 0.765 65.2 0.28 64.98 0.28 64.98 0.765 64.28 0.765 64.28 0.28 64.06 0.28 64.06 0.765 63.36 0.765 63.36 0.28 62.68 0.28 62.68 0.765 61.98 0.765 61.98 0.28 61.76 0.28 61.76 0.765 61.06 0.765 61.06 0.28 60.84 0.28 60.84 0.765 60.14 0.765 60.14 0.28 59.92 0.28 59.92 0.765 59.22 0.765 59.22 0.28 58.08 0.28 58.08 0.765 57.38 0.765 57.38 0.28 57.16 0.28 57.16 0.765 56.46 0.765 56.46 0.28 56.24 0.28 56.24 0.765 55.54 0.765 55.54 0.28 55.32 0.28 55.32 0.765 54.62 0.765 54.62 0.28 54.4 0.28 54.4 0.765 53.7 0.765 53.7 0.28 53.48 0.28 53.48 0.765 52.78 0.765 52.78 0.28 52.56 0.28 52.56 0.765 51.86 0.765 51.86 0.28 51.64 0.28 51.64 0.765 50.94 0.765 50.94 0.28 50.72 0.28 50.72 0.765 50.02 0.765 50.02 0.28 49.8 0.28 49.8 0.765 49.1 0.765 49.1 0.28 48.88 0.28 48.88 0.765 48.18 0.765 48.18 0.28 47.96 0.28 47.96 0.765 47.26 0.765 47.26 0.28 47.04 0.28 47.04 0.765 46.34 0.765 46.34 0.28 46.12 0.28 46.12 0.765 45.42 0.765 45.42 0.28 45.2 0.28 45.2 0.765 44.5 0.765 44.5 0.28 44.28 0.28 44.28 0.765 43.58 0.765 43.58 0.28 43.36 0.28 43.36 0.765 42.66 0.765 42.66 0.28 42.44 0.28 42.44 0.765 41.74 0.765 41.74 0.28 41.06 0.28 41.06 0.765 40.36 0.765 40.36 0.28 40.14 0.28 40.14 0.765 39.44 0.765 39.44 0.28 39.22 0.28 39.22 0.765 38.52 0.765 38.52 0.28 38.3 0.28 38.3 0.765 37.6 0.765 37.6 0.28 37.38 0.28 37.38 0.765 36.68 0.765 36.68 0.28 36.46 0.28 36.46 0.765 35.76 0.765 35.76 0.28 35.08 0.28 35.08 0.765 34.38 0.765 34.38 0.28 34.16 0.28 34.16 0.765 33.46 0.765 33.46 0.28 33.24 0.28 33.24 0.765 32.54 0.765 32.54 0.28 32.32 0.28 32.32 0.765 31.62 0.765 31.62 0.28 31.4 0.28 31.4 0.765 30.7 0.765 30.7 0.28 30.48 0.28 30.48 0.765 29.78 0.765 29.78 0.28 29.1 0.28 29.1 0.765 28.4 0.765 28.4 0.28 28.18 0.28 28.18 0.765 27.48 0.765 27.48 0.28 26.8 0.28 26.8 0.765 26.1 0.765 26.1 0.28 25.88 0.28 25.88 0.765 25.18 0.765 25.18 0.28 24.96 0.28 24.96 0.765 24.26 0.765 24.26 0.28 23.58 0.28 23.58 0.765 22.88 0.765 22.88 0.28 22.66 0.28 22.66 0.765 21.96 0.765 21.96 0.28 21.74 0.28 21.74 0.765 21.04 0.765 21.04 0.28 20.82 0.28 20.82 0.765 20.12 0.765 20.12 0.28 19.9 0.28 19.9 0.765 19.2 0.765 19.2 0.28 18.98 0.28 18.98 0.765 18.28 0.765 18.28 0.28 18.06 0.28 18.06 0.765 17.36 0.765 17.36 0.28 13.92 0.28 13.92 0.765 13.22 0.765 13.22 0.28 11.62 0.28 11.62 0.765 10.92 0.765 10.92 0.28 10.7 0.28 10.7 0.765 10 0.765 10 0.28 7.94 0.28 7.94 0.765 7.24 0.765 7.24 0.28 7.02 0.28 7.02 0.765 6.32 0.765 6.32 0.28 2.88 0.28 2.88 0.765 2.18 0.765 2.18 0.28 0.28 0.28 0.28 86.76 4.48 86.76 4.48 86.275 5.18 86.275 5.18 86.76 5.4 86.76 5.4 86.275 6.1 86.275 6.1 86.76 6.32 86.76 6.32 86.275 7.02 86.275 7.02 86.76 9.54 86.76 9.54 86.275 10.24 86.275 10.24 86.76 10.46 86.76 10.46 86.275 11.16 86.275 11.16 86.76 11.38 86.76 11.38 86.275 12.08 86.275 12.08 86.76 14.6 86.76 14.6 86.275 15.3 86.275 15.3 86.76 15.52 86.76 15.52 86.275 16.22 86.275 16.22 86.76 16.44 86.76 16.44 86.275 17.14 86.275 17.14 86.76 17.36 86.76 17.36 86.275 18.06 86.275 18.06 86.76 18.28 86.76 18.28 86.275 18.98 86.275 18.98 86.76 19.2 86.76 19.2 86.275 19.9 86.275 19.9 86.76 20.12 86.76 20.12 86.275 20.82 86.275 20.82 86.76 21.04 86.76 21.04 86.275 21.74 86.275 21.74 86.76 21.96 86.76 21.96 86.275 22.66 86.275 22.66 86.76 22.88 86.76 22.88 86.275 23.58 86.275 23.58 86.76 23.8 86.76 23.8 86.275 24.5 86.275 24.5 86.76 24.72 86.76 24.72 86.275 25.42 86.275 25.42 86.76 25.64 86.76 25.64 86.275 26.34 86.275 26.34 86.76 27.02 86.76 27.02 86.275 27.72 86.275 27.72 86.76 27.94 86.76 27.94 86.275 28.64 86.275 28.64 86.76 29.78 86.76 29.78 86.275 30.48 86.275 30.48 86.76 30.7 86.76 30.7 86.275 31.4 86.275 31.4 86.76 32.08 86.76 32.08 86.275 32.78 86.275 32.78 86.76 33 86.76 33 86.275 33.7 86.275 33.7 86.76 33.92 86.76 33.92 86.275 34.62 86.275 34.62 86.76 35.3 86.76 35.3 86.275 36 86.275 36 86.76 36.22 86.76 36.22 86.275 36.92 86.275 36.92 86.76 37.14 86.76 37.14 86.275 37.84 86.275 37.84 86.76 38.06 86.76 38.06 86.275 38.76 86.275 38.76 86.76 38.98 86.76 38.98 86.275 39.68 86.275 39.68 86.76 39.9 86.76 39.9 86.275 40.6 86.275 40.6 86.76 40.82 86.76 40.82 86.275 41.52 86.275 41.52 86.76 41.74 86.76 41.74 86.275 42.44 86.275 42.44 86.76 42.66 86.76 42.66 86.275 43.36 86.275 43.36 86.76 43.58 86.76 43.58 86.275 44.28 86.275 44.28 86.76 44.5 86.76 44.5 86.275 45.2 86.275 45.2 86.76 45.42 86.76 45.42 86.275 46.12 86.275 46.12 86.76 46.34 86.76 46.34 86.275 47.04 86.275 47.04 86.76 47.26 86.76 47.26 86.275 47.96 86.275 47.96 86.76 48.18 86.76 48.18 86.275 48.88 86.275 48.88 86.76 49.1 86.76 49.1 86.275 49.8 86.275 49.8 86.76 50.02 86.76 50.02 86.275 50.72 86.275 50.72 86.76 50.94 86.76 50.94 86.275 51.64 86.275 51.64 86.76 51.86 86.76 51.86 86.275 52.56 86.275 52.56 86.76 52.78 86.76 52.78 86.275 53.48 86.275 53.48 86.76 53.7 86.76 53.7 86.275 54.4 86.275 54.4 86.76 54.62 86.76 54.62 86.275 55.32 86.275 55.32 86.76 55.54 86.76 55.54 86.275 56.24 86.275 56.24 86.76 56.46 86.76 56.46 86.275 57.16 86.275 57.16 86.76 57.38 86.76 57.38 86.275 58.08 86.275 58.08 86.76 59.22 86.76 59.22 86.275 59.92 86.275 59.92 86.76 60.14 86.76 60.14 86.275 60.84 86.275 60.84 86.76 61.06 86.76 61.06 86.275 61.76 86.275 61.76 86.76 61.98 86.76 61.98 86.275 62.68 86.275 62.68 86.76 62.9 86.76 62.9 86.275 63.6 86.275 63.6 86.76 63.82 86.76 63.82 86.275 64.52 86.275 64.52 86.76 64.74 86.76 64.74 86.275 65.44 86.275 65.44 86.76 65.66 86.76 65.66 86.275 66.36 86.275 66.36 86.76 ;
    LAYER met4 ;
      POLYGON 26.385 86.865 26.385 86.535 26.37 86.535 26.37 41.67 26.07 41.67 26.07 86.535 26.055 86.535 26.055 86.865 ;
      POLYGON 73.2 86.64 73.2 0.4 59.58 0.4 59.58 1 58.18 1 58.18 0.4 44.86 0.4 44.86 1 43.46 1 43.46 0.4 42.41 0.4 42.41 1.2 41.31 1.2 41.31 0.4 33.21 0.4 33.21 1.2 32.11 1.2 32.11 0.4 31.37 0.4 31.37 1.2 30.27 1.2 30.27 0.4 30.14 0.4 30.14 1 28.74 1 28.74 0.4 15.42 0.4 15.42 1 14.02 1 14.02 0.4 0.4 0.4 0.4 86.64 14.02 86.64 14.02 86.04 15.42 86.04 15.42 86.64 28.74 86.64 28.74 86.04 30.14 86.04 30.14 86.64 30.27 86.64 30.27 85.84 31.37 85.84 31.37 86.64 32.11 86.64 32.11 85.84 33.21 85.84 33.21 86.64 33.95 86.64 33.95 85.84 35.05 85.84 35.05 86.64 43.46 86.64 43.46 86.04 44.86 86.04 44.86 86.64 56.95 86.64 56.95 85.84 58.05 85.84 58.05 86.64 58.18 86.64 58.18 86.04 59.58 86.04 59.58 86.64 59.71 86.64 59.71 85.84 60.81 85.84 60.81 86.64 ;
    LAYER met5 ;
      RECT 4.8 82.72 68.8 85.92 ;
      RECT 4.8 1.12 68.8 4.32 ;
      POLYGON 68.8 85.44 68.8 81.12 72 81.12 72 67.12 68.8 67.12 68.8 60.72 72 60.72 72 46.72 68.8 46.72 68.8 40.32 72 40.32 72 26.32 68.8 26.32 68.8 19.92 72 19.92 72 5.92 68.8 5.92 68.8 1.6 4.8 1.6 4.8 5.92 1.6 5.92 1.6 19.92 4.8 19.92 4.8 26.32 1.6 26.32 1.6 40.32 4.8 40.32 4.8 46.72 1.6 46.72 1.6 60.72 4.8 60.72 4.8 67.12 1.6 67.12 1.6 81.12 4.8 81.12 4.8 85.44 ;
    LAYER li1 ;
      POLYGON 73.6 87.125 73.6 86.955 67.535 86.955 67.535 86.23 67.245 86.23 67.245 86.955 64.695 86.955 64.695 86.555 64.365 86.555 64.365 86.955 63.855 86.955 63.855 86.555 63.525 86.555 63.525 86.955 62.11 86.955 62.11 86.445 61.695 86.445 61.695 86.955 57.485 86.955 57.485 86.155 57.155 86.155 57.155 86.955 56.645 86.955 56.645 86.475 56.315 86.475 56.315 86.955 55.805 86.955 55.805 86.475 55.475 86.475 55.475 86.955 54.965 86.955 54.965 86.475 54.635 86.475 54.635 86.955 54.125 86.955 54.125 86.475 53.795 86.475 53.795 86.955 53.285 86.955 53.285 86.475 52.955 86.475 52.955 86.955 52.355 86.955 52.355 86.23 52.065 86.23 52.065 86.955 49.205 86.955 49.205 86.155 48.875 86.155 48.875 86.955 48.365 86.955 48.365 86.475 48.035 86.475 48.035 86.955 47.525 86.955 47.525 86.475 47.195 86.475 47.195 86.955 46.685 86.955 46.685 86.475 46.355 86.475 46.355 86.955 45.845 86.955 45.845 86.475 45.515 86.475 45.515 86.955 45.005 86.955 45.005 86.475 44.675 86.475 44.675 86.955 43.645 86.955 43.645 86.475 43.315 86.475 43.315 86.955 42.805 86.955 42.805 86.475 42.475 86.475 42.475 86.955 41.965 86.955 41.965 86.475 41.635 86.475 41.635 86.955 41.125 86.955 41.125 86.475 40.795 86.475 40.795 86.955 40.285 86.955 40.285 86.475 39.955 86.475 39.955 86.955 39.445 86.955 39.445 86.155 39.115 86.155 39.115 86.955 37.635 86.955 37.635 86.23 37.345 86.23 37.345 86.955 36.785 86.955 36.785 86.155 36.455 86.155 36.455 86.955 35.945 86.955 35.945 86.475 35.615 86.475 35.615 86.955 35.105 86.955 35.105 86.475 34.775 86.475 34.775 86.955 34.265 86.955 34.265 86.475 33.935 86.475 33.935 86.955 33.425 86.955 33.425 86.475 33.095 86.475 33.095 86.955 32.585 86.955 32.585 86.475 32.255 86.475 32.255 86.955 31.1 86.955 31.1 86.495 30.775 86.495 30.775 86.955 28.985 86.955 28.985 86.495 28.715 86.495 28.715 86.955 27.545 86.955 27.545 86.475 27.215 86.475 27.215 86.955 26.705 86.955 26.705 86.475 26.375 86.475 26.375 86.955 25.865 86.955 25.865 86.475 25.535 86.475 25.535 86.955 25.025 86.955 25.025 86.475 24.695 86.475 24.695 86.955 24.185 86.955 24.185 86.475 23.855 86.475 23.855 86.955 23.345 86.955 23.345 86.155 23.015 86.155 23.015 86.955 22.455 86.955 22.455 86.23 22.165 86.23 22.165 86.955 21.605 86.955 21.605 86.155 21.275 86.155 21.275 86.955 20.765 86.955 20.765 86.475 20.435 86.475 20.435 86.955 19.925 86.955 19.925 86.475 19.595 86.475 19.595 86.955 19.085 86.955 19.085 86.475 18.755 86.475 18.755 86.955 18.245 86.955 18.245 86.475 17.915 86.475 17.915 86.955 17.405 86.955 17.405 86.475 17.075 86.475 17.075 86.955 12.865 86.955 12.865 86.155 12.535 86.155 12.535 86.955 12.025 86.955 12.025 86.475 11.695 86.475 11.695 86.955 11.185 86.955 11.185 86.475 10.855 86.475 10.855 86.955 10.345 86.955 10.345 86.475 10.015 86.475 10.015 86.955 9.505 86.955 9.505 86.475 9.175 86.475 9.175 86.955 8.665 86.955 8.665 86.475 8.335 86.475 8.335 86.955 7.735 86.955 7.735 86.23 7.445 86.23 7.445 86.955 6.535 86.955 6.535 86.42 6.025 86.42 6.025 86.955 4.065 86.955 4.065 86.555 3.735 86.555 3.735 86.955 0 86.955 0 87.125 ;
      RECT 69.92 84.235 73.6 84.405 ;
      RECT 0 84.235 1.84 84.405 ;
      RECT 69.92 81.515 73.6 81.685 ;
      RECT 0 81.515 1.84 81.685 ;
      RECT 72.68 78.795 73.6 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 72.68 76.075 73.6 76.245 ;
      RECT 0 76.075 1.84 76.245 ;
      RECT 69.92 73.355 73.6 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 69.92 70.635 73.6 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 72.68 67.915 73.6 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 72.68 65.195 73.6 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 72.68 62.475 73.6 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 72.68 59.755 73.6 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 72.68 57.035 73.6 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 72.68 54.315 73.6 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 72.68 51.595 73.6 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 72.68 48.875 73.6 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 72.68 46.155 73.6 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 72.68 43.435 73.6 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 72.68 40.715 73.6 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 72.68 37.995 73.6 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 72.68 35.275 73.6 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 72.68 32.555 73.6 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 72.68 29.835 73.6 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 72.68 27.115 73.6 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 72.68 24.395 73.6 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 72.68 21.675 73.6 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 72.68 18.955 73.6 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 72.68 16.235 73.6 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 72.68 13.515 73.6 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 72.68 10.795 73.6 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 72.68 8.075 73.6 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 72.68 5.355 73.6 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 72.68 2.635 73.6 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      POLYGON 63.925 0.885 63.925 0.085 67.245 0.085 67.245 0.81 67.535 0.81 67.535 0.085 73.6 0.085 73.6 -0.085 0 -0.085 0 0.085 3.735 0.085 3.735 0.485 4.065 0.485 4.065 0.085 6.025 0.085 6.025 0.62 6.535 0.62 6.535 0.085 7.445 0.085 7.445 0.81 7.735 0.81 7.735 0.085 8.255 0.085 8.255 0.565 8.425 0.565 8.425 0.085 9.095 0.085 9.095 0.565 9.265 0.565 9.265 0.085 9.855 0.085 9.855 0.565 10.185 0.565 10.185 0.085 10.695 0.085 10.695 0.565 11.025 0.565 11.025 0.085 11.535 0.085 11.535 0.885 11.865 0.885 11.865 0.085 13.435 0.085 13.435 0.885 13.765 0.885 13.765 0.085 14.275 0.085 14.275 0.565 14.605 0.565 14.605 0.085 15.115 0.085 15.115 0.565 15.445 0.565 15.445 0.085 16.035 0.085 16.035 0.565 16.205 0.565 16.205 0.085 16.875 0.085 16.875 0.565 17.045 0.565 17.045 0.085 18.455 0.085 18.455 0.485 18.785 0.485 18.785 0.085 20.745 0.085 20.745 0.62 21.255 0.62 21.255 0.085 22.165 0.085 22.165 0.81 22.455 0.81 22.455 0.085 23.015 0.085 23.015 0.885 23.345 0.885 23.345 0.085 23.855 0.085 23.855 0.565 24.185 0.565 24.185 0.085 24.695 0.085 24.695 0.565 25.025 0.565 25.025 0.085 25.535 0.085 25.535 0.565 25.865 0.565 25.865 0.085 26.375 0.085 26.375 0.565 26.705 0.565 26.705 0.085 27.215 0.085 27.215 0.565 27.545 0.565 27.545 0.085 29.495 0.085 29.495 0.565 29.825 0.565 29.825 0.085 30.335 0.085 30.335 0.565 30.665 0.565 30.665 0.085 31.175 0.085 31.175 0.565 31.505 0.565 31.505 0.085 32.015 0.085 32.015 0.565 32.345 0.565 32.345 0.085 32.855 0.085 32.855 0.565 33.185 0.565 33.185 0.085 33.695 0.085 33.695 0.885 34.025 0.885 34.025 0.085 37.345 0.085 37.345 0.81 37.635 0.81 37.635 0.085 40.535 0.085 40.535 0.565 40.865 0.565 40.865 0.085 41.375 0.085 41.375 0.565 41.705 0.565 41.705 0.085 42.215 0.085 42.215 0.565 42.545 0.565 42.545 0.085 43.055 0.085 43.055 0.565 43.385 0.565 43.385 0.085 43.895 0.085 43.895 0.565 44.225 0.565 44.225 0.085 44.735 0.085 44.735 0.885 45.065 0.885 45.065 0.085 46.975 0.085 46.975 0.565 47.305 0.565 47.305 0.085 47.815 0.085 47.815 0.565 48.145 0.565 48.145 0.085 48.655 0.085 48.655 0.565 48.985 0.565 48.985 0.085 49.495 0.085 49.495 0.565 49.825 0.565 49.825 0.085 50.335 0.085 50.335 0.565 50.665 0.565 50.665 0.085 51.175 0.085 51.175 0.885 51.505 0.885 51.505 0.085 52.065 0.085 52.065 0.81 52.355 0.81 52.355 0.085 52.955 0.085 52.955 0.565 53.285 0.565 53.285 0.085 53.795 0.085 53.795 0.565 54.125 0.565 54.125 0.085 54.635 0.085 54.635 0.565 54.965 0.565 54.965 0.085 55.475 0.085 55.475 0.565 55.805 0.565 55.805 0.085 56.315 0.085 56.315 0.565 56.645 0.565 56.645 0.085 57.155 0.085 57.155 0.885 57.485 0.885 57.485 0.085 59.395 0.085 59.395 0.565 59.725 0.565 59.725 0.085 60.235 0.085 60.235 0.565 60.565 0.565 60.565 0.085 61.075 0.085 61.075 0.565 61.405 0.565 61.405 0.085 61.915 0.085 61.915 0.565 62.245 0.565 62.245 0.085 62.755 0.085 62.755 0.565 63.085 0.565 63.085 0.085 63.595 0.085 63.595 0.885 ;
      RECT 0.17 0.17 73.43 86.87 ;
    LAYER met3 ;
      POLYGON 59.045 87.085 59.045 87.08 59.26 87.08 59.26 86.76 59.045 86.76 59.045 86.755 58.715 86.755 58.715 86.76 58.5 86.76 58.5 87.08 58.715 87.08 58.715 87.085 ;
      POLYGON 29.605 87.085 29.605 87.08 29.82 87.08 29.82 86.76 29.605 86.76 29.605 86.755 29.275 86.755 29.275 86.76 29.06 86.76 29.06 87.08 29.275 87.08 29.275 87.085 ;
      POLYGON 16.035 86.865 16.035 86.85 26.03 86.85 26.03 86.86 26.41 86.86 26.41 86.54 26.03 86.54 26.03 86.55 16.035 86.55 16.035 86.535 15.705 86.535 15.705 86.865 ;
      POLYGON 59.045 0.285 59.045 0.28 59.26 0.28 59.26 -0.04 59.045 -0.04 59.045 -0.045 58.715 -0.045 58.715 -0.04 58.5 -0.04 58.5 0.28 58.715 0.28 58.715 0.285 ;
      POLYGON 29.605 0.285 29.605 0.28 29.82 0.28 29.82 -0.04 29.605 -0.04 29.605 -0.045 29.275 -0.045 29.275 -0.04 29.06 -0.04 29.06 0.28 29.275 0.28 29.275 0.285 ;
      RECT 0.4 0.4 73.2 86.64 ;
    LAYER via ;
      RECT 58.805 86.845 58.955 86.995 ;
      RECT 29.365 86.845 29.515 86.995 ;
      RECT 48.455 86.455 48.605 86.605 ;
      RECT 33.275 86.455 33.425 86.605 ;
      RECT 14.875 86.455 15.025 86.605 ;
      RECT 37.875 0.435 38.025 0.585 ;
      RECT 22.235 0.435 22.385 0.585 ;
      RECT 58.805 0.045 58.955 0.195 ;
      RECT 29.365 0.045 29.515 0.195 ;
    LAYER via2 ;
      RECT 58.78 86.82 58.98 87.02 ;
      RECT 29.34 86.82 29.54 87.02 ;
      RECT 15.77 86.6 15.97 86.8 ;
      RECT 58.78 0.02 58.98 0.22 ;
      RECT 29.34 0.02 29.54 0.22 ;
    LAYER via3 ;
      RECT 58.78 86.82 58.98 87.02 ;
      RECT 29.34 86.82 29.54 87.02 ;
      RECT 26.12 86.6 26.32 86.8 ;
      RECT 60.16 85.92 60.36 86.12 ;
      RECT 58.78 0.02 58.98 0.22 ;
      RECT 29.34 0.02 29.54 0.22 ;
    LAYER via4 ;
      RECT 43.76 84.72 44.56 85.52 ;
      RECT 14.32 84.72 15.12 85.52 ;
      RECT 43.76 1.52 44.56 2.32 ;
      RECT 14.32 1.52 15.12 2.32 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 87.04 73.6 87.04 73.6 0 ;
  END
END cby_2__1_

END LIBRARY
