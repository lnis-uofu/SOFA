//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module sky130_fd_sc_hd__or2_1
(
    A,
    B,
    X
);

    input A;
    input B;
    output X;

    wire A;
    wire B;
    wire X;

endmodule

