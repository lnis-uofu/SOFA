VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO cby_2__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 66.24 BY 76.16 ;
  SYMMETRY X Y ;
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.76 0 50.9 0.485 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.1 0 18.24 0.485 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.84 0 49.98 0.485 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.68 0 51.82 0.485 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.2 0 34.34 0.485 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.86 0 21 0.485 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.14 0 29.28 0.485 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.6 0 52.74 0.485 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 0 41.24 0.485 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.06 0 30.2 0.485 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.78 0 21.92 0.485 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 0 35.72 0.485 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.58 0 12.72 0.485 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.52 0 53.66 0.485 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25 0 25.14 0.485 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.08 0 24.22 0.485 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.6 0 6.74 0.485 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.16 0 46.3 0.485 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.52 0 7.66 0.485 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.24 0 45.38 0.485 ;
    END
  END chany_bottom_in[19]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.58 75.675 12.72 76.16 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.92 75.675 49.06 76.16 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.68 75.675 5.82 76.16 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.5 75.675 36.64 76.16 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.72 75.675 39.86 76.16 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.62 75.675 23.76 76.16 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.56 75.675 41.7 76.16 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.48 75.675 42.62 76.16 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.28 75.675 33.42 76.16 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.54 75.675 24.68 76.16 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.36 75.675 9.5 76.16 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 75.675 35.72 76.16 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.2 75.675 34.34 76.16 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.74 75.675 56.88 76.16 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.52 75.675 30.66 76.16 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.36 75.675 32.5 76.16 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.24 75.675 22.38 76.16 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.08 75.675 47.22 76.16 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.98 75.675 8.12 76.16 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.16 75.675 46.3 76.16 ;
    END
  END chany_top_in[19]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 6.31 0.8 6.61 ;
    END
  END ccff_head[0]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.98 0 31.12 0.485 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.28 0 33.42 0.485 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 0 39.4 0.485 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.32 0 44.46 0.485 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.42 0 37.56 0.485 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.02 0 42.16 0.485 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.38 0 26.52 0.485 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.3 0 27.44 0.485 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.94 0 20.08 0.485 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.18 0 40.32 0.485 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 0 38.48 0.485 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.92 0 49.06 0.485 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.5 0 36.64 0.485 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.08 0 47.22 0.485 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.22 0 28.36 0.485 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.36 0 32.5 0.485 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.7 0 22.84 0.485 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48 0 48.14 0.485 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.02 0 19.16 0.485 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.4 0 43.54 0.485 ;
    END
  END chany_bottom_out[19]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.32 75.675 44.46 76.16 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.82 75.675 55.96 76.16 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.44 75.675 31.58 76.16 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.44 75.675 54.58 76.16 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.8 75.675 38.94 76.16 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.76 75.675 50.9 76.16 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.6 75.675 29.74 76.16 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48 75.675 48.14 76.16 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.88 75.675 38.02 76.16 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.4 75.675 43.54 76.16 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.38 75.675 26.52 76.16 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.24 75.675 45.38 76.16 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.84 75.675 49.98 76.16 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.6 75.675 52.74 76.16 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.68 75.675 28.82 76.16 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.64 75.675 40.78 76.16 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.32 75.675 21.46 76.16 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.68 75.675 51.82 76.16 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.3 75.675 27.44 76.16 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.52 75.675 53.66 76.16 ;
    END
  END chany_top_out[19]
  PIN right_grid_pin_0_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 14.47 0.8 14.77 ;
    END
  END right_grid_pin_0_[0]
  PIN left_grid_pin_16_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 26.03 0.8 26.33 ;
    END
  END left_grid_pin_16_[0]
  PIN left_grid_pin_17_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 21.95 0.8 22.25 ;
    END
  END left_grid_pin_17_[0]
  PIN left_grid_pin_18_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 23.31 0.8 23.61 ;
    END
  END left_grid_pin_18_[0]
  PIN left_grid_pin_19_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.03 0.8 43.33 ;
    END
  END left_grid_pin_19_[0]
  PIN left_grid_pin_20_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 45.75 0.8 46.05 ;
    END
  END left_grid_pin_20_[0]
  PIN left_grid_pin_21_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 47.11 0.8 47.41 ;
    END
  END left_grid_pin_21_[0]
  PIN left_grid_pin_22_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.39 0.8 44.69 ;
    END
  END left_grid_pin_22_[0]
  PIN left_grid_pin_23_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 24.67 0.8 24.97 ;
    END
  END left_grid_pin_23_[0]
  PIN left_grid_pin_24_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 49.83 0.8 50.13 ;
    END
  END left_grid_pin_24_[0]
  PIN left_grid_pin_25_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 19.23 0.8 19.53 ;
    END
  END left_grid_pin_25_[0]
  PIN left_grid_pin_26_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 4.95 0.8 5.25 ;
    END
  END left_grid_pin_26_[0]
  PIN left_grid_pin_27_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 7.67 0.8 7.97 ;
    END
  END left_grid_pin_27_[0]
  PIN left_grid_pin_28_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 10.39 0.8 10.69 ;
    END
  END left_grid_pin_28_[0]
  PIN left_grid_pin_29_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 9.03 0.8 9.33 ;
    END
  END left_grid_pin_29_[0]
  PIN left_grid_pin_30_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.47 0.8 48.77 ;
    END
  END left_grid_pin_30_[0]
  PIN left_grid_pin_31_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 20.59 0.8 20.89 ;
    END
  END left_grid_pin_31_[0]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.76 0 4.9 0.485 ;
    END
  END ccff_tail[0]
  PIN IO_ISOL_N[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 11.75 0.8 12.05 ;
    END
  END IO_ISOL_N[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65.44 10.39 66.24 10.69 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65.44 6.31 66.24 6.61 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65.44 4.95 66.24 5.25 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN left_width_0_height_0__pin_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 13.11 0.8 13.41 ;
    END
  END left_width_0_height_0__pin_0_[0]
  PIN left_width_0_height_0__pin_1_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.6 75.675 6.74 76.16 ;
    END
  END left_width_0_height_0__pin_1_upper[0]
  PIN left_width_0_height_0__pin_1_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.68 0 5.82 0.485 ;
    END
  END left_width_0_height_0__pin_1_lower[0]
  PIN prog_clk_0_W_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met3 ;
        RECT 0 3.59 0.8 3.89 ;
    END
  END prog_clk_0_W_in
  PIN prog_clk_0_S_out
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 11.66 0 11.8 0.485 ;
    END
  END prog_clk_0_S_out
  PIN prog_clk_0_N_out
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 13.5 75.675 13.64 76.16 ;
    END
  END prog_clk_0_N_out
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 65.76 2.48 66.24 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 65.76 7.92 66.24 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 65.76 13.36 66.24 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 65.76 18.8 66.24 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 65.76 24.24 66.24 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 65.76 29.68 66.24 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 65.76 35.12 66.24 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 65.76 40.56 66.24 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 65.76 46 66.24 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 65.76 51.44 66.24 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 65.76 56.88 66.24 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 65.76 62.32 66.24 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 65.76 67.76 66.24 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 65.76 73.2 66.24 73.68 ;
      LAYER met4 ;
        RECT 10.74 0 11.34 0.6 ;
        RECT 40.18 0 40.78 0.6 ;
        RECT 10.74 75.56 11.34 76.16 ;
        RECT 40.18 75.56 40.78 76.16 ;
      LAYER met5 ;
        RECT 0 5.88 3.2 9.08 ;
        RECT 63.04 5.88 66.24 9.08 ;
        RECT 0 46.68 3.2 49.88 ;
        RECT 63.04 46.68 66.24 49.88 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 0 45.4 0.24 ;
        RECT 46.6 0 66.24 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 65.76 5.2 66.24 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 65.76 10.64 66.24 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 65.76 16.08 66.24 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 65.76 21.52 66.24 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 65.76 26.96 66.24 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 65.76 32.4 66.24 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 65.76 37.84 66.24 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 65.76 43.28 66.24 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 65.76 48.72 66.24 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 65.76 54.16 66.24 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 65.76 59.6 66.24 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 65.76 65.04 66.24 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 65.76 70.48 66.24 70.96 ;
        RECT 0 75.92 45.4 76.16 ;
        RECT 46.6 75.92 66.24 76.16 ;
      LAYER met4 ;
        RECT 25.46 0 26.06 0.6 ;
        RECT 54.9 0 55.5 0.6 ;
        RECT 25.46 75.56 26.06 76.16 ;
        RECT 54.9 75.56 55.5 76.16 ;
      LAYER met5 ;
        RECT 0 26.28 3.2 29.48 ;
        RECT 63.04 26.28 66.24 29.48 ;
        RECT 0 67.08 3.2 70.28 ;
        RECT 63.04 67.08 66.24 70.28 ;
    END
  END VSS
  OBS
    LAYER met2 ;
      RECT 55.06 75.975 55.34 76.345 ;
      RECT 25.62 75.975 25.9 76.345 ;
      RECT 55.06 -0.185 55.34 0.185 ;
      RECT 25.62 -0.185 25.9 0.185 ;
      POLYGON 65.96 75.88 65.96 0.28 53.94 0.28 53.94 0.765 53.24 0.765 53.24 0.28 53.02 0.28 53.02 0.765 52.32 0.765 52.32 0.28 52.1 0.28 52.1 0.765 51.4 0.765 51.4 0.28 51.18 0.28 51.18 0.765 50.48 0.765 50.48 0.28 50.26 0.28 50.26 0.765 49.56 0.765 49.56 0.28 49.34 0.28 49.34 0.765 48.64 0.765 48.64 0.28 48.42 0.28 48.42 0.765 47.72 0.765 47.72 0.28 47.5 0.28 47.5 0.765 46.8 0.765 46.8 0.28 46.58 0.28 46.58 0.765 45.88 0.765 45.88 0.28 45.66 0.28 45.66 0.765 44.96 0.765 44.96 0.28 44.74 0.28 44.74 0.765 44.04 0.765 44.04 0.28 43.82 0.28 43.82 0.765 43.12 0.765 43.12 0.28 42.44 0.28 42.44 0.765 41.74 0.765 41.74 0.28 41.52 0.28 41.52 0.765 40.82 0.765 40.82 0.28 40.6 0.28 40.6 0.765 39.9 0.765 39.9 0.28 39.68 0.28 39.68 0.765 38.98 0.765 38.98 0.28 38.76 0.28 38.76 0.765 38.06 0.765 38.06 0.28 37.84 0.28 37.84 0.765 37.14 0.765 37.14 0.28 36.92 0.28 36.92 0.765 36.22 0.765 36.22 0.28 36 0.28 36 0.765 35.3 0.765 35.3 0.28 34.62 0.28 34.62 0.765 33.92 0.765 33.92 0.28 33.7 0.28 33.7 0.765 33 0.765 33 0.28 32.78 0.28 32.78 0.765 32.08 0.765 32.08 0.28 31.4 0.28 31.4 0.765 30.7 0.765 30.7 0.28 30.48 0.28 30.48 0.765 29.78 0.765 29.78 0.28 29.56 0.28 29.56 0.765 28.86 0.765 28.86 0.28 28.64 0.28 28.64 0.765 27.94 0.765 27.94 0.28 27.72 0.28 27.72 0.765 27.02 0.765 27.02 0.28 26.8 0.28 26.8 0.765 26.1 0.765 26.1 0.28 25.42 0.28 25.42 0.765 24.72 0.765 24.72 0.28 24.5 0.28 24.5 0.765 23.8 0.765 23.8 0.28 23.12 0.28 23.12 0.765 22.42 0.765 22.42 0.28 22.2 0.28 22.2 0.765 21.5 0.765 21.5 0.28 21.28 0.28 21.28 0.765 20.58 0.765 20.58 0.28 20.36 0.28 20.36 0.765 19.66 0.765 19.66 0.28 19.44 0.28 19.44 0.765 18.74 0.765 18.74 0.28 18.52 0.28 18.52 0.765 17.82 0.765 17.82 0.28 13 0.28 13 0.765 12.3 0.765 12.3 0.28 12.08 0.28 12.08 0.765 11.38 0.765 11.38 0.28 7.94 0.28 7.94 0.765 7.24 0.765 7.24 0.28 7.02 0.28 7.02 0.765 6.32 0.765 6.32 0.28 6.1 0.28 6.1 0.765 5.4 0.765 5.4 0.28 5.18 0.28 5.18 0.765 4.48 0.765 4.48 0.28 0.28 0.28 0.28 75.88 5.4 75.88 5.4 75.395 6.1 75.395 6.1 75.88 6.32 75.88 6.32 75.395 7.02 75.395 7.02 75.88 7.7 75.88 7.7 75.395 8.4 75.395 8.4 75.88 9.08 75.88 9.08 75.395 9.78 75.395 9.78 75.88 12.3 75.88 12.3 75.395 13 75.395 13 75.88 13.22 75.88 13.22 75.395 13.92 75.395 13.92 75.88 21.04 75.88 21.04 75.395 21.74 75.395 21.74 75.88 21.96 75.88 21.96 75.395 22.66 75.395 22.66 75.88 23.34 75.88 23.34 75.395 24.04 75.395 24.04 75.88 24.26 75.88 24.26 75.395 24.96 75.395 24.96 75.88 26.1 75.88 26.1 75.395 26.8 75.395 26.8 75.88 27.02 75.88 27.02 75.395 27.72 75.395 27.72 75.88 28.4 75.88 28.4 75.395 29.1 75.395 29.1 75.88 29.32 75.88 29.32 75.395 30.02 75.395 30.02 75.88 30.24 75.88 30.24 75.395 30.94 75.395 30.94 75.88 31.16 75.88 31.16 75.395 31.86 75.395 31.86 75.88 32.08 75.88 32.08 75.395 32.78 75.395 32.78 75.88 33 75.88 33 75.395 33.7 75.395 33.7 75.88 33.92 75.88 33.92 75.395 34.62 75.395 34.62 75.88 35.3 75.88 35.3 75.395 36 75.395 36 75.88 36.22 75.88 36.22 75.395 36.92 75.395 36.92 75.88 37.6 75.88 37.6 75.395 38.3 75.395 38.3 75.88 38.52 75.88 38.52 75.395 39.22 75.395 39.22 75.88 39.44 75.88 39.44 75.395 40.14 75.395 40.14 75.88 40.36 75.88 40.36 75.395 41.06 75.395 41.06 75.88 41.28 75.88 41.28 75.395 41.98 75.395 41.98 75.88 42.2 75.88 42.2 75.395 42.9 75.395 42.9 75.88 43.12 75.88 43.12 75.395 43.82 75.395 43.82 75.88 44.04 75.88 44.04 75.395 44.74 75.395 44.74 75.88 44.96 75.88 44.96 75.395 45.66 75.395 45.66 75.88 45.88 75.88 45.88 75.395 46.58 75.395 46.58 75.88 46.8 75.88 46.8 75.395 47.5 75.395 47.5 75.88 47.72 75.88 47.72 75.395 48.42 75.395 48.42 75.88 48.64 75.88 48.64 75.395 49.34 75.395 49.34 75.88 49.56 75.88 49.56 75.395 50.26 75.395 50.26 75.88 50.48 75.88 50.48 75.395 51.18 75.395 51.18 75.88 51.4 75.88 51.4 75.395 52.1 75.395 52.1 75.88 52.32 75.88 52.32 75.395 53.02 75.395 53.02 75.88 53.24 75.88 53.24 75.395 53.94 75.395 53.94 75.88 54.16 75.88 54.16 75.395 54.86 75.395 54.86 75.88 55.54 75.88 55.54 75.395 56.24 75.395 56.24 75.88 56.46 75.88 56.46 75.395 57.16 75.395 57.16 75.88 ;
    LAYER met3 ;
      POLYGON 55.365 76.325 55.365 76.32 55.58 76.32 55.58 76 55.365 76 55.365 75.995 55.035 75.995 55.035 76 54.82 76 54.82 76.32 55.035 76.32 55.035 76.325 ;
      POLYGON 25.925 76.325 25.925 76.32 26.14 76.32 26.14 76 25.925 76 25.925 75.995 25.595 75.995 25.595 76 25.38 76 25.38 76.32 25.595 76.32 25.595 76.325 ;
      POLYGON 7.74 12.73 7.74 12.43 0.65 12.43 0.65 12.71 1.2 12.71 1.2 12.73 ;
      POLYGON 55.365 0.165 55.365 0.16 55.58 0.16 55.58 -0.16 55.365 -0.16 55.365 -0.165 55.035 -0.165 55.035 -0.16 54.82 -0.16 54.82 0.16 55.035 0.16 55.035 0.165 ;
      POLYGON 25.925 0.165 25.925 0.16 26.14 0.16 26.14 -0.16 25.925 -0.16 25.925 -0.165 25.595 -0.165 25.595 -0.16 25.38 -0.16 25.38 0.16 25.595 0.16 25.595 0.165 ;
      POLYGON 65.84 75.76 65.84 11.09 65.04 11.09 65.04 9.99 65.84 9.99 65.84 7.01 65.04 7.01 65.04 5.91 65.84 5.91 65.84 5.65 65.04 5.65 65.04 4.55 65.84 4.55 65.84 0.4 0.4 0.4 0.4 3.19 1.2 3.19 1.2 4.29 0.4 4.29 0.4 4.55 1.2 4.55 1.2 5.65 0.4 5.65 0.4 5.91 1.2 5.91 1.2 7.01 0.4 7.01 0.4 7.27 1.2 7.27 1.2 8.37 0.4 8.37 0.4 8.63 1.2 8.63 1.2 9.73 0.4 9.73 0.4 9.99 1.2 9.99 1.2 11.09 0.4 11.09 0.4 11.35 1.2 11.35 1.2 12.45 0.4 12.45 0.4 12.71 1.2 12.71 1.2 13.81 0.4 13.81 0.4 14.07 1.2 14.07 1.2 15.17 0.4 15.17 0.4 18.83 1.2 18.83 1.2 19.93 0.4 19.93 0.4 20.19 1.2 20.19 1.2 21.29 0.4 21.29 0.4 21.55 1.2 21.55 1.2 22.65 0.4 22.65 0.4 22.91 1.2 22.91 1.2 24.01 0.4 24.01 0.4 24.27 1.2 24.27 1.2 25.37 0.4 25.37 0.4 25.63 1.2 25.63 1.2 26.73 0.4 26.73 0.4 42.63 1.2 42.63 1.2 43.73 0.4 43.73 0.4 43.99 1.2 43.99 1.2 45.09 0.4 45.09 0.4 45.35 1.2 45.35 1.2 46.45 0.4 46.45 0.4 46.71 1.2 46.71 1.2 47.81 0.4 47.81 0.4 48.07 1.2 48.07 1.2 49.17 0.4 49.17 0.4 49.43 1.2 49.43 1.2 50.53 0.4 50.53 0.4 75.76 ;
    LAYER met5 ;
      POLYGON 64.64 74.56 64.64 71.88 61.44 71.88 61.44 65.48 64.64 65.48 64.64 51.48 61.44 51.48 61.44 45.08 64.64 45.08 64.64 31.08 61.44 31.08 61.44 24.68 64.64 24.68 64.64 10.68 61.44 10.68 61.44 4.28 64.64 4.28 64.64 1.6 1.6 1.6 1.6 4.28 4.8 4.28 4.8 10.68 1.6 10.68 1.6 24.68 4.8 24.68 4.8 31.08 1.6 31.08 1.6 45.08 4.8 45.08 4.8 51.48 1.6 51.48 1.6 65.48 4.8 65.48 4.8 71.88 1.6 71.88 1.6 74.56 ;
    LAYER met4 ;
      POLYGON 65.84 75.76 65.84 0.4 55.9 0.4 55.9 1 54.5 1 54.5 0.4 41.18 0.4 41.18 1 39.78 1 39.78 0.4 26.46 0.4 26.46 1 25.06 1 25.06 0.4 11.74 0.4 11.74 1 10.34 1 10.34 0.4 0.4 0.4 0.4 75.76 10.34 75.76 10.34 75.16 11.74 75.16 11.74 75.76 25.06 75.76 25.06 75.16 26.46 75.16 26.46 75.76 39.78 75.76 39.78 75.16 41.18 75.16 41.18 75.76 54.5 75.76 54.5 75.16 55.9 75.16 55.9 75.76 ;
    LAYER met1 ;
      RECT 45.68 75.92 46.32 76.4 ;
      RECT 45.68 -0.24 46.32 0.24 ;
      POLYGON 46.32 75.88 46.32 75.64 65.96 75.64 65.96 73.96 65.48 73.96 65.48 72.92 65.96 72.92 65.96 71.24 65.48 71.24 65.48 70.2 65.96 70.2 65.96 68.52 65.48 68.52 65.48 67.48 65.96 67.48 65.96 65.8 65.48 65.8 65.48 64.76 65.96 64.76 65.96 63.08 65.48 63.08 65.48 62.04 65.96 62.04 65.96 60.36 65.48 60.36 65.48 59.32 65.96 59.32 65.96 57.64 65.48 57.64 65.48 56.6 65.96 56.6 65.96 54.92 65.48 54.92 65.48 53.88 65.96 53.88 65.96 52.2 65.48 52.2 65.48 51.16 65.96 51.16 65.96 49.48 65.48 49.48 65.48 48.44 65.96 48.44 65.96 46.76 65.48 46.76 65.48 45.72 65.96 45.72 65.96 44.04 65.48 44.04 65.48 43 65.96 43 65.96 41.32 65.48 41.32 65.48 40.28 65.96 40.28 65.96 38.6 65.48 38.6 65.48 37.56 65.96 37.56 65.96 35.88 65.48 35.88 65.48 34.84 65.96 34.84 65.96 33.16 65.48 33.16 65.48 32.12 65.96 32.12 65.96 30.44 65.48 30.44 65.48 29.4 65.96 29.4 65.96 27.72 65.48 27.72 65.48 26.68 65.96 26.68 65.96 25 65.48 25 65.48 23.96 65.96 23.96 65.96 22.28 65.48 22.28 65.48 21.24 65.96 21.24 65.96 19.56 65.48 19.56 65.48 18.52 65.96 18.52 65.96 16.84 65.48 16.84 65.48 15.8 65.96 15.8 65.96 14.12 65.48 14.12 65.48 13.08 65.96 13.08 65.96 11.4 65.48 11.4 65.48 10.36 65.96 10.36 65.96 8.68 65.48 8.68 65.48 7.64 65.96 7.64 65.96 5.96 65.48 5.96 65.48 4.92 65.96 4.92 65.96 3.24 65.48 3.24 65.48 2.2 65.96 2.2 65.96 0.52 46.32 0.52 46.32 0.28 45.68 0.28 45.68 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 45.68 75.64 45.68 75.88 ;
    LAYER li1 ;
      RECT 0 76.075 66.24 76.245 ;
      RECT 62.56 73.355 66.24 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 65.32 70.635 66.24 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 65.32 67.915 66.24 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 65.32 65.195 66.24 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 65.32 62.475 66.24 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 65.32 59.755 66.24 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 65.32 57.035 66.24 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 65.32 54.315 66.24 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 65.32 51.595 66.24 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 65.32 48.875 66.24 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 65.32 46.155 66.24 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 65.32 43.435 66.24 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 65.32 40.715 66.24 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 65.32 37.995 66.24 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 65.32 35.275 66.24 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 65.32 32.555 66.24 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 65.32 29.835 66.24 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 65.32 27.115 66.24 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 65.32 24.395 66.24 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 65.32 21.675 66.24 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 65.32 18.955 66.24 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 65.32 16.235 66.24 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 65.32 13.515 66.24 13.685 ;
      RECT 0 13.515 1.84 13.685 ;
      RECT 65.32 10.795 66.24 10.965 ;
      RECT 0 10.795 1.84 10.965 ;
      RECT 65.32 8.075 66.24 8.245 ;
      RECT 0 8.075 1.84 8.245 ;
      RECT 65.32 5.355 66.24 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 62.56 2.635 66.24 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 66.24 0.085 ;
      RECT 0.17 0.17 66.07 75.99 ;
    LAYER via ;
      RECT 55.125 76.085 55.275 76.235 ;
      RECT 25.685 76.085 25.835 76.235 ;
      RECT 55.125 -0.075 55.275 0.075 ;
      RECT 25.685 -0.075 25.835 0.075 ;
    LAYER via2 ;
      RECT 55.1 76.06 55.3 76.26 ;
      RECT 25.66 76.06 25.86 76.26 ;
      RECT 1.05 45.8 1.25 46 ;
      RECT 64.99 6.36 65.19 6.56 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER via3 ;
      RECT 55.1 76.06 55.3 76.26 ;
      RECT 25.66 76.06 25.86 76.26 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 76.16 66.24 76.16 66.24 0 ;
  END
END cby_2__1_

END LIBRARY
