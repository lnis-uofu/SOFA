//
//
//
//
//
//
//
//
`timescale 1ns / 1ps

//
module const0(const0);
//
output [0:0] const0;

//
//


//
//

	assign const0[0] = 1'b0;
endmodule
//

//
module const1(const1);
//
output [0:0] const1;

//
//


//
//

	assign const1[0] = 1'b1;
endmodule
//


