VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_1__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 117.76 BY 108.8 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 52.83 0 52.97 1.36 ;
    END
  END prog_clk[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.87 107.44 64.01 108.8 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.27 107.44 59.41 108.8 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 67.93 107.44 68.23 108.8 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.13 107.44 78.27 108.8 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.35 107.44 58.49 108.8 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.93 107.44 69.07 108.8 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 107.44 46.53 108.8 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.53 107.44 73.67 108.8 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.51 107.44 56.65 108.8 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.21 107.44 77.35 108.8 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.17 107.44 66.31 108.8 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.63 107.44 43.77 108.8 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.33 107.44 63.63 108.8 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.61 107.44 49.75 108.8 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.19 107.44 83.33 108.8 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 107.44 45.61 108.8 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.05 107.44 79.19 108.8 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.09 107.44 67.23 108.8 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.55 107.44 44.69 108.8 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.65 107.44 60.79 108.8 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.13 96.56 9.27 97.92 ;
    END
  END top_left_grid_pin_42_[0]
  PIN top_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.83 96.56 6.97 97.92 ;
    END
  END top_left_grid_pin_43_[0]
  PIN top_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.81 96.56 12.95 97.92 ;
    END
  END top_left_grid_pin_44_[0]
  PIN top_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.99 107.44 28.13 108.8 ;
    END
  END top_left_grid_pin_45_[0]
  PIN top_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.19 96.56 14.33 97.92 ;
    END
  END top_left_grid_pin_46_[0]
  PIN top_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.75 96.56 7.89 97.92 ;
    END
  END top_left_grid_pin_47_[0]
  PIN top_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.03 96.56 16.17 97.92 ;
    END
  END top_left_grid_pin_48_[0]
  PIN top_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.91 107.44 29.05 108.8 ;
    END
  END top_left_grid_pin_49_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 66.49 117.76 66.79 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 82.81 117.76 83.11 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 92.33 117.76 92.63 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 36.57 117.76 36.87 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 74.65 117.76 74.95 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 77.37 117.76 77.67 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 33.85 117.76 34.15 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 46.09 117.76 46.39 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 56.97 117.76 57.27 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 73.29 117.76 73.59 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 84.17 117.76 84.47 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 90.97 117.76 91.27 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 81.45 117.76 81.75 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 44.73 117.76 45.03 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 31.81 117.76 32.11 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 61.73 117.76 62.03 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 65.13 117.76 65.43 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 48.81 117.76 49.11 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 69.21 117.76 69.51 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 89.61 117.76 89.91 ;
    END
  END chanx_right_in[19]
  PIN right_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.41 10.88 109.55 12.24 ;
    END
  END right_bottom_grid_pin_34_[0]
  PIN right_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.71 10.88 111.85 12.24 ;
    END
  END right_bottom_grid_pin_35_[0]
  PIN right_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.01 10.88 114.15 12.24 ;
    END
  END right_bottom_grid_pin_36_[0]
  PIN right_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.49 10.88 108.63 12.24 ;
    END
  END right_bottom_grid_pin_37_[0]
  PIN right_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.79 10.88 110.93 12.24 ;
    END
  END right_bottom_grid_pin_38_[0]
  PIN right_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.09 10.88 113.23 12.24 ;
    END
  END right_bottom_grid_pin_39_[0]
  PIN right_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.59 10.88 101.73 12.24 ;
    END
  END right_bottom_grid_pin_40_[0]
  PIN right_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.19 10.88 106.33 12.24 ;
    END
  END right_bottom_grid_pin_41_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.21 0 77.35 1.36 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.93 0 69.07 1.36 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.05 0 79.19 1.36 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.85 0 69.99 1.36 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.25 0 65.39 1.36 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.27 0 59.41 1.36 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.85 0 46.99 1.36 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.19 0 60.33 1.36 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.77 0 47.91 1.36 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.09 0 67.23 1.36 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.01 0 68.15 1.36 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.77 0 70.91 1.36 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.49 0 62.63 1.36 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.11 0 61.25 1.36 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.69 0 48.83 1.36 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.97 0 57.11 1.36 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.13 0 78.27 1.36 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.93 0 46.07 1.36 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.61 0 49.75 1.36 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.61 0 72.75 1.36 ;
    END
  END chany_bottom_in[19]
  PIN bottom_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 12.73 10.88 13.03 12.24 ;
    END
  END bottom_left_grid_pin_42_[0]
  PIN bottom_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 9.05 10.88 9.35 12.24 ;
    END
  END bottom_left_grid_pin_43_[0]
  PIN bottom_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.99 0 28.13 1.36 ;
    END
  END bottom_left_grid_pin_44_[0]
  PIN bottom_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.29 10.88 7.43 12.24 ;
    END
  END bottom_left_grid_pin_45_[0]
  PIN bottom_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.13 10.88 9.27 12.24 ;
    END
  END bottom_left_grid_pin_46_[0]
  PIN bottom_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.11 10.88 15.25 12.24 ;
    END
  END bottom_left_grid_pin_47_[0]
  PIN bottom_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.21 10.88 8.35 12.24 ;
    END
  END bottom_left_grid_pin_48_[0]
  PIN bottom_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.05 10.88 10.19 12.24 ;
    END
  END bottom_left_grid_pin_49_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 66.49 1.38 66.79 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 84.17 1.38 84.47 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 85.53 1.38 85.83 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.25 1.38 37.55 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.05 1.38 44.35 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.81 1.38 32.11 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 89.61 1.38 89.91 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 65.13 1.38 65.43 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.97 1.38 57.27 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 81.45 1.38 81.75 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 49.49 1.38 49.79 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 75.33 1.38 75.63 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 92.33 1.38 92.63 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 45.41 1.38 45.71 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 86.89 1.38 87.19 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 71.25 1.38 71.55 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 41.33 1.38 41.63 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 38.61 1.38 38.91 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 73.97 1.38 74.27 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 72.61 1.38 72.91 ;
    END
  END chanx_left_in[19]
  PIN left_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.91 0 29.05 1.36 ;
    END
  END left_bottom_grid_pin_34_[0]
  PIN left_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.81 10.88 12.95 12.24 ;
    END
  END left_bottom_grid_pin_35_[0]
  PIN left_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.99 10.88 5.13 12.24 ;
    END
  END left_bottom_grid_pin_36_[0]
  PIN left_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.07 10.88 4.21 12.24 ;
    END
  END left_bottom_grid_pin_37_[0]
  PIN left_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.37 10.88 6.51 12.24 ;
    END
  END left_bottom_grid_pin_38_[0]
  PIN left_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 4.45 10.88 4.75 12.24 ;
    END
  END left_bottom_grid_pin_39_[0]
  PIN left_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.89 10.88 12.03 12.24 ;
    END
  END left_bottom_grid_pin_40_[0]
  PIN left_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.03 10.88 16.17 12.24 ;
    END
  END left_bottom_grid_pin_41_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 43.37 117.76 43.67 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.97 107.44 80.11 108.8 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.49 107.44 62.63 108.8 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 107.44 47.45 108.8 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.37 107.44 75.51 108.8 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.37 107.44 52.51 108.8 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.29 107.44 76.43 108.8 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 107.44 57.57 108.8 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.85 107.44 69.99 108.8 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 107.44 48.37 108.8 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.23 107.44 71.37 108.8 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.57 107.44 61.71 108.8 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.79 107.44 64.93 108.8 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.11 107.44 84.25 108.8 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.01 107.44 68.15 108.8 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.43 107.44 34.57 108.8 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.61 107.44 72.75 108.8 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.53 107.44 50.67 108.8 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.45 107.44 74.59 108.8 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.29 107.44 53.43 108.8 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.27 107.44 82.41 108.8 ;
    END
  END chany_top_out[19]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 70.57 117.76 70.87 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 55.61 117.76 55.91 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 71.93 117.76 72.23 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 54.25 117.76 54.55 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 37.93 117.76 38.23 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 80.09 117.76 80.39 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 50.17 117.76 50.47 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 63.77 117.76 64.07 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 42.01 117.76 42.31 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 51.53 117.76 51.83 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 52.89 117.76 53.19 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 39.29 117.76 39.59 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 78.73 117.76 79.03 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 67.85 117.76 68.15 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 35.21 117.76 35.51 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 40.65 117.76 40.95 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 58.33 117.76 58.63 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 47.45 117.76 47.75 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 59.69 117.76 59.99 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 76.01 117.76 76.31 ;
    END
  END chanx_right_out[19]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.87 0 64.01 1.36 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.01 0 45.15 1.36 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.13 0 55.27 1.36 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.17 0 66.31 1.36 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.35 0 58.49 1.36 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.37 0 75.51 1.36 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.53 0 50.67 1.36 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.53 0 73.67 1.36 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.73 0 82.87 1.36 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.45 0 74.59 1.36 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.05 0 56.19 1.36 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.69 0 71.83 1.36 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.97 0 80.11 1.36 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.29 0 76.43 1.36 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.43 0 34.57 1.36 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.25 0 88.39 1.36 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.81 0 81.95 1.36 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.33 0 87.47 1.36 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.21 0 54.35 1.36 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.17 0 89.31 1.36 ;
    END
  END chany_bottom_out[19]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 82.81 1.38 83.11 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 63.77 1.38 64.07 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.01 1.38 59.31 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.13 1.38 48.43 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 62.41 1.38 62.71 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 88.25 1.38 88.55 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 46.77 1.38 47.07 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.85 1.38 51.15 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 54.93 1.38 55.23 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.21 1.38 52.51 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 61.05 1.38 61.35 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 68.53 1.38 68.83 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.69 1.38 42.99 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 90.97 1.38 91.27 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.17 1.38 33.47 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 78.73 1.38 79.03 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.89 1.38 70.19 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.97 1.38 40.27 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 53.57 1.38 53.87 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 80.09 1.38 80.39 ;
    END
  END chanx_left_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 76.69 1.38 76.99 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 25.76 2.48 26.24 2.96 ;
        RECT 91.52 2.48 92 2.96 ;
        RECT 25.76 7.92 26.24 8.4 ;
        RECT 91.52 7.92 92 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 117.28 13.36 117.76 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 117.28 18.8 117.76 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 117.28 24.24 117.76 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 117.28 29.68 117.76 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 117.28 35.12 117.76 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 117.28 40.56 117.76 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 117.28 46 117.76 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 117.28 51.44 117.76 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 117.28 56.88 117.76 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 117.28 62.32 117.76 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 117.28 67.76 117.76 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 117.28 73.2 117.76 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 117.28 78.64 117.76 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 117.28 84.08 117.76 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 117.28 89.52 117.76 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 117.28 94.96 117.76 95.44 ;
        RECT 25.76 100.4 26.24 100.88 ;
        RECT 91.52 100.4 92 100.88 ;
        RECT 25.76 105.84 26.24 106.32 ;
        RECT 91.52 105.84 92 106.32 ;
      LAYER met4 ;
        RECT 36.5 0 37.1 0.6 ;
        RECT 65.94 0 66.54 0.6 ;
        RECT 106.42 10.88 107.02 11.48 ;
        RECT 106.42 97.32 107.02 97.92 ;
        RECT 36.5 108.2 37.1 108.8 ;
        RECT 65.94 108.2 66.54 108.8 ;
      LAYER met5 ;
        RECT 0 22.2 3.2 25.4 ;
        RECT 114.56 22.2 117.76 25.4 ;
        RECT 0 63 3.2 66.2 ;
        RECT 114.56 63 117.76 66.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 25.76 0 92 0.24 ;
        RECT 25.76 5.2 26.24 5.68 ;
        RECT 91.52 5.2 92 5.68 ;
        RECT 0 10.64 117.76 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 117.28 16.08 117.76 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 117.28 21.52 117.76 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 117.28 26.96 117.76 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 117.28 32.4 117.76 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 117.28 37.84 117.76 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 117.28 43.28 117.76 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 117.28 48.72 117.76 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 117.28 54.16 117.76 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 117.28 59.6 117.76 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 117.28 65.04 117.76 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 117.28 70.48 117.76 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 117.28 75.92 117.76 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 117.28 81.36 117.76 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 117.28 86.8 117.76 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 117.28 92.24 117.76 92.72 ;
        RECT 0 97.68 117.76 98.16 ;
        RECT 25.76 103.12 26.24 103.6 ;
        RECT 91.52 103.12 92 103.6 ;
        RECT 25.76 108.56 92 108.8 ;
      LAYER met4 ;
        RECT 51.22 0 51.82 0.6 ;
        RECT 80.66 0 81.26 0.6 ;
        RECT 10.74 10.88 11.34 11.48 ;
        RECT 10.74 97.32 11.34 97.92 ;
        RECT 51.22 108.2 51.82 108.8 ;
        RECT 80.66 108.2 81.26 108.8 ;
      LAYER met5 ;
        RECT 0 42.6 3.2 45.8 ;
        RECT 114.56 42.6 117.76 45.8 ;
        RECT 0 83.4 3.2 86.6 ;
        RECT 114.56 83.4 117.76 86.6 ;
    END
  END VSS
  PIN prog_clk__FEEDTHRU_1[0]
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 55.13 107.44 55.27 108.8 ;
    END
  END prog_clk__FEEDTHRU_1[0]
  PIN Test_en__FEEDTHRU_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.23 96.56 2.37 97.92 ;
    END
  END Test_en__FEEDTHRU_0[0]
  PIN Test_en__FEEDTHRU_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.23 10.88 2.37 12.24 ;
    END
  END Test_en__FEEDTHRU_1[0]
  PIN clk__FEEDTHRU_0[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 3.15 96.56 3.29 97.92 ;
    END
  END clk__FEEDTHRU_0[0]
  PIN clk__FEEDTHRU_1[0]
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 3.15 10.88 3.29 12.24 ;
    END
  END clk__FEEDTHRU_1[0]
  PIN grid_clb_0_bottom_width_0_height_0__pin_50___FEEDTHRU_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.33 10.88 18.47 12.24 ;
    END
  END grid_clb_0_bottom_width_0_height_0__pin_50___FEEDTHRU_0[0]
  PIN grid_clb_0_bottom_width_0_height_0__pin_50___FEEDTHRU_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.29 96.56 99.43 97.92 ;
    END
  END grid_clb_0_bottom_width_0_height_0__pin_50___FEEDTHRU_1[0]
  OBS
    LAYER li1 ;
      RECT 25.76 108.715 92 108.885 ;
      RECT 91.54 105.995 92 106.165 ;
      RECT 25.76 105.995 29.44 106.165 ;
      RECT 91.08 103.275 92 103.445 ;
      RECT 25.76 103.275 27.6 103.445 ;
      RECT 91.08 100.555 92 100.725 ;
      RECT 25.76 100.555 29.44 100.725 ;
      RECT 89.24 97.835 117.76 98.005 ;
      RECT 0 97.835 29.44 98.005 ;
      RECT 116.84 95.115 117.76 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 114.08 92.395 117.76 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 114.08 89.675 117.76 89.845 ;
      RECT 0 89.675 1.84 89.845 ;
      RECT 117.3 86.955 117.76 87.125 ;
      RECT 0 86.955 1.84 87.125 ;
      RECT 117.3 84.235 117.76 84.405 ;
      RECT 0 84.235 1.84 84.405 ;
      RECT 115.92 81.515 117.76 81.685 ;
      RECT 0 81.515 1.84 81.685 ;
      RECT 115.92 78.795 117.76 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 116.84 76.075 117.76 76.245 ;
      RECT 0 76.075 1.84 76.245 ;
      RECT 116.84 73.355 117.76 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 116.84 70.635 117.76 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 116.84 67.915 117.76 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 116.84 65.195 117.76 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 116.84 62.475 117.76 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 116.84 59.755 117.76 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 116.84 57.035 117.76 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 116.84 54.315 117.76 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 116.84 51.595 117.76 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 116.84 48.875 117.76 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 116.84 46.155 117.76 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 116.84 43.435 117.76 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 116.84 40.715 117.76 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 116.84 37.995 117.76 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 116.84 35.275 117.76 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 116.84 32.555 117.76 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 116.84 29.835 117.76 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 114.08 27.115 117.76 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 114.08 24.395 117.76 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 116.84 21.675 117.76 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 116.84 18.955 117.76 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 116.84 16.235 117.76 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 117.3 13.515 117.76 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 88.78 10.795 117.76 10.965 ;
      RECT 0 10.795 29.44 10.965 ;
      RECT 91.08 8.075 92 8.245 ;
      RECT 25.76 8.075 29.44 8.245 ;
      RECT 91.08 5.355 92 5.525 ;
      RECT 25.76 5.355 29.44 5.525 ;
      RECT 91.08 2.635 92 2.805 ;
      RECT 25.76 2.635 29.44 2.805 ;
      RECT 25.76 -0.085 92 0.085 ;
    LAYER met2 ;
      RECT 80.82 108.615 81.1 108.985 ;
      RECT 51.38 108.615 51.66 108.985 ;
      RECT 74.85 106.94 75.11 107.26 ;
      RECT 66.57 106.94 66.83 107.26 ;
      RECT 65.19 106.94 65.45 107.26 ;
      RECT 46.79 106.94 47.05 107.26 ;
      RECT 10.9 97.735 11.18 98.105 ;
      RECT 107.97 12.42 108.23 12.74 ;
      RECT 10.9 10.695 11.18 11.065 ;
      RECT 68.41 1.54 68.67 1.86 ;
      RECT 57.37 1.54 57.63 1.86 ;
      RECT 50.93 1.54 51.19 1.86 ;
      RECT 80.82 -0.185 81.1 0.185 ;
      RECT 51.38 -0.185 51.66 0.185 ;
      POLYGON 91.72 108.52 91.72 97.64 99.01 97.64 99.01 96.28 99.71 96.28 99.71 97.64 117.48 97.64 117.48 11.16 114.43 11.16 114.43 12.52 113.73 12.52 113.73 11.16 113.51 11.16 113.51 12.52 112.81 12.52 112.81 11.16 112.13 11.16 112.13 12.52 111.43 12.52 111.43 11.16 111.21 11.16 111.21 12.52 110.51 12.52 110.51 11.16 109.83 11.16 109.83 12.52 109.13 12.52 109.13 11.16 108.91 11.16 108.91 12.52 108.21 12.52 108.21 11.16 106.61 11.16 106.61 12.52 105.91 12.52 105.91 11.16 102.01 11.16 102.01 12.52 101.31 12.52 101.31 11.16 91.72 11.16 91.72 0.28 89.59 0.28 89.59 1.64 88.89 1.64 88.89 0.28 88.67 0.28 88.67 1.64 87.97 1.64 87.97 0.28 87.75 0.28 87.75 1.64 87.05 1.64 87.05 0.28 83.15 0.28 83.15 1.64 82.45 1.64 82.45 0.28 82.23 0.28 82.23 1.64 81.53 1.64 81.53 0.28 80.39 0.28 80.39 1.64 79.69 1.64 79.69 0.28 79.47 0.28 79.47 1.64 78.77 1.64 78.77 0.28 78.55 0.28 78.55 1.64 77.85 1.64 77.85 0.28 77.63 0.28 77.63 1.64 76.93 1.64 76.93 0.28 76.71 0.28 76.71 1.64 76.01 1.64 76.01 0.28 75.79 0.28 75.79 1.64 75.09 1.64 75.09 0.28 74.87 0.28 74.87 1.64 74.17 1.64 74.17 0.28 73.95 0.28 73.95 1.64 73.25 1.64 73.25 0.28 73.03 0.28 73.03 1.64 72.33 1.64 72.33 0.28 72.11 0.28 72.11 1.64 71.41 1.64 71.41 0.28 71.19 0.28 71.19 1.64 70.49 1.64 70.49 0.28 70.27 0.28 70.27 1.64 69.57 1.64 69.57 0.28 69.35 0.28 69.35 1.64 68.65 1.64 68.65 0.28 68.43 0.28 68.43 1.64 67.73 1.64 67.73 0.28 67.51 0.28 67.51 1.64 66.81 1.64 66.81 0.28 66.59 0.28 66.59 1.64 65.89 1.64 65.89 0.28 65.67 0.28 65.67 1.64 64.97 1.64 64.97 0.28 64.29 0.28 64.29 1.64 63.59 1.64 63.59 0.28 62.91 0.28 62.91 1.64 62.21 1.64 62.21 0.28 61.53 0.28 61.53 1.64 60.83 1.64 60.83 0.28 60.61 0.28 60.61 1.64 59.91 1.64 59.91 0.28 59.69 0.28 59.69 1.64 58.99 1.64 58.99 0.28 58.77 0.28 58.77 1.64 58.07 1.64 58.07 0.28 57.39 0.28 57.39 1.64 56.69 1.64 56.69 0.28 56.47 0.28 56.47 1.64 55.77 1.64 55.77 0.28 55.55 0.28 55.55 1.64 54.85 1.64 54.85 0.28 54.63 0.28 54.63 1.64 53.93 1.64 53.93 0.28 53.25 0.28 53.25 1.64 52.55 1.64 52.55 0.28 50.95 0.28 50.95 1.64 50.25 1.64 50.25 0.28 50.03 0.28 50.03 1.64 49.33 1.64 49.33 0.28 49.11 0.28 49.11 1.64 48.41 1.64 48.41 0.28 48.19 0.28 48.19 1.64 47.49 1.64 47.49 0.28 47.27 0.28 47.27 1.64 46.57 1.64 46.57 0.28 46.35 0.28 46.35 1.64 45.65 1.64 45.65 0.28 45.43 0.28 45.43 1.64 44.73 1.64 44.73 0.28 34.85 0.28 34.85 1.64 34.15 1.64 34.15 0.28 29.33 0.28 29.33 1.64 28.63 1.64 28.63 0.28 28.41 0.28 28.41 1.64 27.71 1.64 27.71 0.28 26.04 0.28 26.04 11.16 18.75 11.16 18.75 12.52 18.05 12.52 18.05 11.16 16.45 11.16 16.45 12.52 15.75 12.52 15.75 11.16 15.53 11.16 15.53 12.52 14.83 12.52 14.83 11.16 13.23 11.16 13.23 12.52 12.53 12.52 12.53 11.16 12.31 11.16 12.31 12.52 11.61 12.52 11.61 11.16 10.47 11.16 10.47 12.52 9.77 12.52 9.77 11.16 9.55 11.16 9.55 12.52 8.85 12.52 8.85 11.16 8.63 11.16 8.63 12.52 7.93 12.52 7.93 11.16 7.71 11.16 7.71 12.52 7.01 12.52 7.01 11.16 6.79 11.16 6.79 12.52 6.09 12.52 6.09 11.16 5.41 11.16 5.41 12.52 4.71 12.52 4.71 11.16 4.49 11.16 4.49 12.52 3.79 12.52 3.79 11.16 3.57 11.16 3.57 12.52 2.87 12.52 2.87 11.16 2.65 11.16 2.65 12.52 1.95 12.52 1.95 11.16 0.28 11.16 0.28 97.64 1.95 97.64 1.95 96.28 2.65 96.28 2.65 97.64 2.87 97.64 2.87 96.28 3.57 96.28 3.57 97.64 6.55 97.64 6.55 96.28 7.25 96.28 7.25 97.64 7.47 97.64 7.47 96.28 8.17 96.28 8.17 97.64 8.85 97.64 8.85 96.28 9.55 96.28 9.55 97.64 12.53 97.64 12.53 96.28 13.23 96.28 13.23 97.64 13.91 97.64 13.91 96.28 14.61 96.28 14.61 97.64 15.75 97.64 15.75 96.28 16.45 96.28 16.45 97.64 26.04 97.64 26.04 108.52 27.71 108.52 27.71 107.16 28.41 107.16 28.41 108.52 28.63 108.52 28.63 107.16 29.33 107.16 29.33 108.52 34.15 108.52 34.15 107.16 34.85 107.16 34.85 108.52 43.35 108.52 43.35 107.16 44.05 107.16 44.05 108.52 44.27 108.52 44.27 107.16 44.97 107.16 44.97 108.52 45.19 108.52 45.19 107.16 45.89 107.16 45.89 108.52 46.11 108.52 46.11 107.16 46.81 107.16 46.81 108.52 47.03 108.52 47.03 107.16 47.73 107.16 47.73 108.52 47.95 108.52 47.95 107.16 48.65 107.16 48.65 108.52 49.33 108.52 49.33 107.16 50.03 107.16 50.03 108.52 50.25 108.52 50.25 107.16 50.95 107.16 50.95 108.52 52.09 108.52 52.09 107.16 52.79 107.16 52.79 108.52 53.01 108.52 53.01 107.16 53.71 107.16 53.71 108.52 54.85 108.52 54.85 107.16 55.55 107.16 55.55 108.52 56.23 108.52 56.23 107.16 56.93 107.16 56.93 108.52 57.15 108.52 57.15 107.16 57.85 107.16 57.85 108.52 58.07 108.52 58.07 107.16 58.77 107.16 58.77 108.52 58.99 108.52 58.99 107.16 59.69 107.16 59.69 108.52 60.37 108.52 60.37 107.16 61.07 107.16 61.07 108.52 61.29 108.52 61.29 107.16 61.99 107.16 61.99 108.52 62.21 108.52 62.21 107.16 62.91 107.16 62.91 108.52 63.59 108.52 63.59 107.16 64.29 107.16 64.29 108.52 64.51 108.52 64.51 107.16 65.21 107.16 65.21 108.52 65.89 108.52 65.89 107.16 66.59 107.16 66.59 108.52 66.81 108.52 66.81 107.16 67.51 107.16 67.51 108.52 67.73 108.52 67.73 107.16 68.43 107.16 68.43 108.52 68.65 108.52 68.65 107.16 69.35 107.16 69.35 108.52 69.57 108.52 69.57 107.16 70.27 107.16 70.27 108.52 70.95 108.52 70.95 107.16 71.65 107.16 71.65 108.52 72.33 108.52 72.33 107.16 73.03 107.16 73.03 108.52 73.25 108.52 73.25 107.16 73.95 107.16 73.95 108.52 74.17 108.52 74.17 107.16 74.87 107.16 74.87 108.52 75.09 108.52 75.09 107.16 75.79 107.16 75.79 108.52 76.01 108.52 76.01 107.16 76.71 107.16 76.71 108.52 76.93 108.52 76.93 107.16 77.63 107.16 77.63 108.52 77.85 108.52 77.85 107.16 78.55 107.16 78.55 108.52 78.77 108.52 78.77 107.16 79.47 107.16 79.47 108.52 79.69 108.52 79.69 107.16 80.39 107.16 80.39 108.52 81.99 108.52 81.99 107.16 82.69 107.16 82.69 108.52 82.91 108.52 82.91 107.16 83.61 107.16 83.61 108.52 83.83 108.52 83.83 107.16 84.53 107.16 84.53 108.52 ;
    LAYER met4 ;
      POLYGON 91.6 108.4 91.6 97.52 106.02 97.52 106.02 96.92 107.42 96.92 107.42 97.52 117.36 97.52 117.36 11.28 107.42 11.28 107.42 11.88 106.02 11.88 106.02 11.28 91.6 11.28 91.6 0.4 81.66 0.4 81.66 1 80.26 1 80.26 0.4 66.94 0.4 66.94 1 65.54 1 65.54 0.4 52.22 0.4 52.22 1 50.82 1 50.82 0.4 37.5 0.4 37.5 1 36.1 1 36.1 0.4 26.16 0.4 26.16 11.28 13.43 11.28 13.43 12.64 12.33 12.64 12.33 11.28 11.74 11.28 11.74 11.88 10.34 11.88 10.34 11.28 9.75 11.28 9.75 12.64 8.65 12.64 8.65 11.28 5.15 11.28 5.15 12.64 4.05 12.64 4.05 11.28 0.4 11.28 0.4 97.52 10.34 97.52 10.34 96.92 11.74 96.92 11.74 97.52 26.16 97.52 26.16 108.4 36.1 108.4 36.1 107.8 37.5 107.8 37.5 108.4 50.82 108.4 50.82 107.8 52.22 107.8 52.22 108.4 62.93 108.4 62.93 107.04 64.03 107.04 64.03 108.4 65.54 108.4 65.54 107.8 66.94 107.8 66.94 108.4 67.53 108.4 67.53 107.04 68.63 107.04 68.63 108.4 80.26 108.4 80.26 107.8 81.66 107.8 81.66 108.4 ;
    LAYER met3 ;
      POLYGON 81.125 108.965 81.125 108.96 81.34 108.96 81.34 108.64 81.125 108.64 81.125 108.635 80.795 108.635 80.795 108.64 80.58 108.64 80.58 108.96 80.795 108.96 80.795 108.965 ;
      POLYGON 51.685 108.965 51.685 108.96 51.9 108.96 51.9 108.64 51.685 108.64 51.685 108.635 51.355 108.635 51.355 108.64 51.14 108.64 51.14 108.96 51.355 108.96 51.355 108.965 ;
      POLYGON 11.205 98.085 11.205 98.08 11.42 98.08 11.42 97.76 11.205 97.76 11.205 97.755 10.875 97.755 10.875 97.76 10.66 97.76 10.66 98.08 10.875 98.08 10.875 98.085 ;
      POLYGON 15.79 87.87 15.79 87.57 1.78 87.57 1.78 87.59 1.23 87.59 1.23 87.87 ;
      POLYGON 116.11 72.92 116.11 72.6 115.73 72.6 115.73 72.61 107.49 72.61 107.49 72.91 115.73 72.91 115.73 72.92 ;
      POLYGON 17.63 66.11 17.63 65.81 1.78 65.81 1.78 65.83 1.23 65.83 1.23 66.11 ;
      POLYGON 2.005 57.965 2.005 57.96 2.03 57.96 2.03 57.64 2.005 57.64 2.005 57.635 1.275 57.635 1.275 57.965 ;
      POLYGON 19.01 46.39 19.01 46.09 1.78 46.09 1.78 46.11 1.23 46.11 1.23 46.39 ;
      POLYGON 11.205 11.045 11.205 11.04 11.42 11.04 11.42 10.72 11.205 10.72 11.205 10.715 10.875 10.715 10.875 10.72 10.66 10.72 10.66 11.04 10.875 11.04 10.875 11.045 ;
      POLYGON 81.125 0.165 81.125 0.16 81.34 0.16 81.34 -0.16 81.125 -0.16 81.125 -0.165 80.795 -0.165 80.795 -0.16 80.58 -0.16 80.58 0.16 80.795 0.16 80.795 0.165 ;
      POLYGON 51.685 0.165 51.685 0.16 51.9 0.16 51.9 -0.16 51.685 -0.16 51.685 -0.165 51.355 -0.165 51.355 -0.16 51.14 -0.16 51.14 0.16 51.355 0.16 51.355 0.165 ;
      POLYGON 91.6 108.4 91.6 97.52 117.36 97.52 117.36 93.03 115.98 93.03 115.98 91.93 117.36 91.93 117.36 91.67 115.98 91.67 115.98 90.57 117.36 90.57 117.36 90.31 115.98 90.31 115.98 89.21 117.36 89.21 117.36 84.87 115.98 84.87 115.98 83.77 117.36 83.77 117.36 83.51 115.98 83.51 115.98 82.41 117.36 82.41 117.36 82.15 115.98 82.15 115.98 81.05 117.36 81.05 117.36 80.79 115.98 80.79 115.98 79.69 117.36 79.69 117.36 79.43 115.98 79.43 115.98 78.33 117.36 78.33 117.36 78.07 115.98 78.07 115.98 76.97 117.36 76.97 117.36 76.71 115.98 76.71 115.98 75.61 117.36 75.61 117.36 75.35 115.98 75.35 115.98 74.25 117.36 74.25 117.36 73.99 115.98 73.99 115.98 72.89 117.36 72.89 117.36 72.63 115.98 72.63 115.98 71.53 117.36 71.53 117.36 71.27 115.98 71.27 115.98 70.17 117.36 70.17 117.36 69.91 115.98 69.91 115.98 68.81 117.36 68.81 117.36 68.55 115.98 68.55 115.98 67.45 117.36 67.45 117.36 67.19 115.98 67.19 115.98 66.09 117.36 66.09 117.36 65.83 115.98 65.83 115.98 64.73 117.36 64.73 117.36 64.47 115.98 64.47 115.98 63.37 117.36 63.37 117.36 62.43 115.98 62.43 115.98 61.33 117.36 61.33 117.36 60.39 115.98 60.39 115.98 59.29 117.36 59.29 117.36 59.03 115.98 59.03 115.98 57.93 117.36 57.93 117.36 57.67 115.98 57.67 115.98 56.57 117.36 56.57 117.36 56.31 115.98 56.31 115.98 55.21 117.36 55.21 117.36 54.95 115.98 54.95 115.98 53.85 117.36 53.85 117.36 53.59 115.98 53.59 115.98 52.49 117.36 52.49 117.36 52.23 115.98 52.23 115.98 51.13 117.36 51.13 117.36 50.87 115.98 50.87 115.98 49.77 117.36 49.77 117.36 49.51 115.98 49.51 115.98 48.41 117.36 48.41 117.36 48.15 115.98 48.15 115.98 47.05 117.36 47.05 117.36 46.79 115.98 46.79 115.98 45.69 117.36 45.69 117.36 45.43 115.98 45.43 115.98 44.33 117.36 44.33 117.36 44.07 115.98 44.07 115.98 42.97 117.36 42.97 117.36 42.71 115.98 42.71 115.98 41.61 117.36 41.61 117.36 41.35 115.98 41.35 115.98 40.25 117.36 40.25 117.36 39.99 115.98 39.99 115.98 38.89 117.36 38.89 117.36 38.63 115.98 38.63 115.98 37.53 117.36 37.53 117.36 37.27 115.98 37.27 115.98 36.17 117.36 36.17 117.36 35.91 115.98 35.91 115.98 34.81 117.36 34.81 117.36 34.55 115.98 34.55 115.98 33.45 117.36 33.45 117.36 32.51 115.98 32.51 115.98 31.41 117.36 31.41 117.36 11.28 91.6 11.28 91.6 0.4 26.16 0.4 26.16 11.28 0.4 11.28 0.4 31.41 1.78 31.41 1.78 32.51 0.4 32.51 0.4 32.77 1.78 32.77 1.78 33.87 0.4 33.87 0.4 36.85 1.78 36.85 1.78 37.95 0.4 37.95 0.4 38.21 1.78 38.21 1.78 39.31 0.4 39.31 0.4 39.57 1.78 39.57 1.78 40.67 0.4 40.67 0.4 40.93 1.78 40.93 1.78 42.03 0.4 42.03 0.4 42.29 1.78 42.29 1.78 43.39 0.4 43.39 0.4 43.65 1.78 43.65 1.78 44.75 0.4 44.75 0.4 45.01 1.78 45.01 1.78 46.11 0.4 46.11 0.4 46.37 1.78 46.37 1.78 47.47 0.4 47.47 0.4 47.73 1.78 47.73 1.78 48.83 0.4 48.83 0.4 49.09 1.78 49.09 1.78 50.19 0.4 50.19 0.4 50.45 1.78 50.45 1.78 51.55 0.4 51.55 0.4 51.81 1.78 51.81 1.78 52.91 0.4 52.91 0.4 53.17 1.78 53.17 1.78 54.27 0.4 54.27 0.4 54.53 1.78 54.53 1.78 55.63 0.4 55.63 0.4 56.57 1.78 56.57 1.78 57.67 0.4 57.67 0.4 58.61 1.78 58.61 1.78 59.71 0.4 59.71 0.4 60.65 1.78 60.65 1.78 61.75 0.4 61.75 0.4 62.01 1.78 62.01 1.78 63.11 0.4 63.11 0.4 63.37 1.78 63.37 1.78 64.47 0.4 64.47 0.4 64.73 1.78 64.73 1.78 65.83 0.4 65.83 0.4 66.09 1.78 66.09 1.78 67.19 0.4 67.19 0.4 68.13 1.78 68.13 1.78 69.23 0.4 69.23 0.4 69.49 1.78 69.49 1.78 70.59 0.4 70.59 0.4 70.85 1.78 70.85 1.78 71.95 0.4 71.95 0.4 72.21 1.78 72.21 1.78 73.31 0.4 73.31 0.4 73.57 1.78 73.57 1.78 74.67 0.4 74.67 0.4 74.93 1.78 74.93 1.78 76.03 0.4 76.03 0.4 76.29 1.78 76.29 1.78 77.39 0.4 77.39 0.4 78.33 1.78 78.33 1.78 79.43 0.4 79.43 0.4 79.69 1.78 79.69 1.78 80.79 0.4 80.79 0.4 81.05 1.78 81.05 1.78 82.15 0.4 82.15 0.4 82.41 1.78 82.41 1.78 83.51 0.4 83.51 0.4 83.77 1.78 83.77 1.78 84.87 0.4 84.87 0.4 85.13 1.78 85.13 1.78 86.23 0.4 86.23 0.4 86.49 1.78 86.49 1.78 87.59 0.4 87.59 0.4 87.85 1.78 87.85 1.78 88.95 0.4 88.95 0.4 89.21 1.78 89.21 1.78 90.31 0.4 90.31 0.4 90.57 1.78 90.57 1.78 91.67 0.4 91.67 0.4 91.93 1.78 91.93 1.78 93.03 0.4 93.03 0.4 97.52 26.16 97.52 26.16 108.4 ;
    LAYER met5 ;
      POLYGON 90.4 107.2 90.4 96.32 116.16 96.32 116.16 88.2 112.96 88.2 112.96 81.8 116.16 81.8 116.16 67.8 112.96 67.8 112.96 61.4 116.16 61.4 116.16 47.4 112.96 47.4 112.96 41 116.16 41 116.16 27 112.96 27 112.96 20.6 116.16 20.6 116.16 12.48 90.4 12.48 90.4 1.6 27.36 1.6 27.36 12.48 1.6 12.48 1.6 20.6 4.8 20.6 4.8 27 1.6 27 1.6 41 4.8 41 4.8 47.4 1.6 47.4 1.6 61.4 4.8 61.4 4.8 67.8 1.6 67.8 1.6 81.8 4.8 81.8 4.8 88.2 1.6 88.2 1.6 96.32 27.36 96.32 27.36 107.2 ;
    LAYER met1 ;
      POLYGON 91.72 108.28 91.72 106.6 91.24 106.6 91.24 105.56 91.72 105.56 91.72 103.88 91.24 103.88 91.24 102.84 91.72 102.84 91.72 101.16 91.24 101.16 91.24 100.12 91.72 100.12 91.72 98.44 26.04 98.44 26.04 100.12 26.52 100.12 26.52 101.16 26.04 101.16 26.04 102.84 26.52 102.84 26.52 103.88 26.04 103.88 26.04 105.56 26.52 105.56 26.52 106.6 26.04 106.6 26.04 108.28 ;
      POLYGON 117.48 97.4 117.48 95.72 117 95.72 117 94.68 117.48 94.68 117.48 93 117 93 117 91.96 117.48 91.96 117.48 90.28 117 90.28 117 89.24 117.48 89.24 117.48 87.56 117 87.56 117 86.52 117.48 86.52 117.48 84.84 117 84.84 117 83.8 117.48 83.8 117.48 82.12 117 82.12 117 81.08 117.48 81.08 117.48 79.4 117 79.4 117 78.36 117.48 78.36 117.48 76.68 117 76.68 117 75.64 117.48 75.64 117.48 73.96 117 73.96 117 72.92 117.48 72.92 117.48 71.24 117 71.24 117 70.2 117.48 70.2 117.48 68.52 117 68.52 117 67.48 117.48 67.48 117.48 65.8 117 65.8 117 64.76 117.48 64.76 117.48 63.08 117 63.08 117 62.04 117.48 62.04 117.48 60.36 117 60.36 117 59.32 117.48 59.32 117.48 57.64 117 57.64 117 56.6 117.48 56.6 117.48 54.92 117 54.92 117 53.88 117.48 53.88 117.48 52.2 117 52.2 117 51.16 117.48 51.16 117.48 49.48 117 49.48 117 48.44 117.48 48.44 117.48 46.76 117 46.76 117 45.72 117.48 45.72 117.48 44.04 117 44.04 117 43 117.48 43 117.48 41.32 117 41.32 117 40.28 117.48 40.28 117.48 38.6 117 38.6 117 37.56 117.48 37.56 117.48 35.88 117 35.88 117 34.84 117.48 34.84 117.48 33.16 117 33.16 117 32.12 117.48 32.12 117.48 30.44 117 30.44 117 29.4 117.48 29.4 117.48 27.72 117 27.72 117 26.68 117.48 26.68 117.48 25 117 25 117 23.96 117.48 23.96 117.48 22.28 117 22.28 117 21.24 117.48 21.24 117.48 19.56 117 19.56 117 18.52 117.48 18.52 117.48 16.84 117 16.84 117 15.8 117.48 15.8 117.48 14.12 117 14.12 117 13.08 117.48 13.08 117.48 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 ;
      POLYGON 91.72 10.36 91.72 8.68 91.24 8.68 91.24 7.64 91.72 7.64 91.72 5.96 91.24 5.96 91.24 4.92 91.72 4.92 91.72 3.24 91.24 3.24 91.24 2.2 91.72 2.2 91.72 0.52 26.04 0.52 26.04 2.2 26.52 2.2 26.52 3.24 26.04 3.24 26.04 4.92 26.52 4.92 26.52 5.96 26.04 5.96 26.04 7.64 26.52 7.64 26.52 8.68 26.04 8.68 26.04 10.36 ;
    LAYER li1 ;
      POLYGON 91.83 108.63 91.83 97.75 117.59 97.75 117.59 11.05 91.83 11.05 91.83 0.17 25.93 0.17 25.93 11.05 0.17 11.05 0.17 97.75 25.93 97.75 25.93 108.63 ;
    LAYER mcon ;
      RECT 91.685 108.715 91.855 108.885 ;
      RECT 91.225 108.715 91.395 108.885 ;
      RECT 90.765 108.715 90.935 108.885 ;
      RECT 90.305 108.715 90.475 108.885 ;
      RECT 89.845 108.715 90.015 108.885 ;
      RECT 89.385 108.715 89.555 108.885 ;
      RECT 88.925 108.715 89.095 108.885 ;
      RECT 88.465 108.715 88.635 108.885 ;
      RECT 88.005 108.715 88.175 108.885 ;
      RECT 87.545 108.715 87.715 108.885 ;
      RECT 87.085 108.715 87.255 108.885 ;
      RECT 86.625 108.715 86.795 108.885 ;
      RECT 86.165 108.715 86.335 108.885 ;
      RECT 85.705 108.715 85.875 108.885 ;
      RECT 85.245 108.715 85.415 108.885 ;
      RECT 84.785 108.715 84.955 108.885 ;
      RECT 84.325 108.715 84.495 108.885 ;
      RECT 83.865 108.715 84.035 108.885 ;
      RECT 83.405 108.715 83.575 108.885 ;
      RECT 82.945 108.715 83.115 108.885 ;
      RECT 82.485 108.715 82.655 108.885 ;
      RECT 82.025 108.715 82.195 108.885 ;
      RECT 81.565 108.715 81.735 108.885 ;
      RECT 81.105 108.715 81.275 108.885 ;
      RECT 80.645 108.715 80.815 108.885 ;
      RECT 80.185 108.715 80.355 108.885 ;
      RECT 79.725 108.715 79.895 108.885 ;
      RECT 79.265 108.715 79.435 108.885 ;
      RECT 78.805 108.715 78.975 108.885 ;
      RECT 78.345 108.715 78.515 108.885 ;
      RECT 77.885 108.715 78.055 108.885 ;
      RECT 77.425 108.715 77.595 108.885 ;
      RECT 76.965 108.715 77.135 108.885 ;
      RECT 76.505 108.715 76.675 108.885 ;
      RECT 76.045 108.715 76.215 108.885 ;
      RECT 75.585 108.715 75.755 108.885 ;
      RECT 75.125 108.715 75.295 108.885 ;
      RECT 74.665 108.715 74.835 108.885 ;
      RECT 74.205 108.715 74.375 108.885 ;
      RECT 73.745 108.715 73.915 108.885 ;
      RECT 73.285 108.715 73.455 108.885 ;
      RECT 72.825 108.715 72.995 108.885 ;
      RECT 72.365 108.715 72.535 108.885 ;
      RECT 71.905 108.715 72.075 108.885 ;
      RECT 71.445 108.715 71.615 108.885 ;
      RECT 70.985 108.715 71.155 108.885 ;
      RECT 70.525 108.715 70.695 108.885 ;
      RECT 70.065 108.715 70.235 108.885 ;
      RECT 69.605 108.715 69.775 108.885 ;
      RECT 69.145 108.715 69.315 108.885 ;
      RECT 68.685 108.715 68.855 108.885 ;
      RECT 68.225 108.715 68.395 108.885 ;
      RECT 67.765 108.715 67.935 108.885 ;
      RECT 67.305 108.715 67.475 108.885 ;
      RECT 66.845 108.715 67.015 108.885 ;
      RECT 66.385 108.715 66.555 108.885 ;
      RECT 65.925 108.715 66.095 108.885 ;
      RECT 65.465 108.715 65.635 108.885 ;
      RECT 65.005 108.715 65.175 108.885 ;
      RECT 64.545 108.715 64.715 108.885 ;
      RECT 64.085 108.715 64.255 108.885 ;
      RECT 63.625 108.715 63.795 108.885 ;
      RECT 63.165 108.715 63.335 108.885 ;
      RECT 62.705 108.715 62.875 108.885 ;
      RECT 62.245 108.715 62.415 108.885 ;
      RECT 61.785 108.715 61.955 108.885 ;
      RECT 61.325 108.715 61.495 108.885 ;
      RECT 60.865 108.715 61.035 108.885 ;
      RECT 60.405 108.715 60.575 108.885 ;
      RECT 59.945 108.715 60.115 108.885 ;
      RECT 59.485 108.715 59.655 108.885 ;
      RECT 59.025 108.715 59.195 108.885 ;
      RECT 58.565 108.715 58.735 108.885 ;
      RECT 58.105 108.715 58.275 108.885 ;
      RECT 57.645 108.715 57.815 108.885 ;
      RECT 57.185 108.715 57.355 108.885 ;
      RECT 56.725 108.715 56.895 108.885 ;
      RECT 56.265 108.715 56.435 108.885 ;
      RECT 55.805 108.715 55.975 108.885 ;
      RECT 55.345 108.715 55.515 108.885 ;
      RECT 54.885 108.715 55.055 108.885 ;
      RECT 54.425 108.715 54.595 108.885 ;
      RECT 53.965 108.715 54.135 108.885 ;
      RECT 53.505 108.715 53.675 108.885 ;
      RECT 53.045 108.715 53.215 108.885 ;
      RECT 52.585 108.715 52.755 108.885 ;
      RECT 52.125 108.715 52.295 108.885 ;
      RECT 51.665 108.715 51.835 108.885 ;
      RECT 51.205 108.715 51.375 108.885 ;
      RECT 50.745 108.715 50.915 108.885 ;
      RECT 50.285 108.715 50.455 108.885 ;
      RECT 49.825 108.715 49.995 108.885 ;
      RECT 49.365 108.715 49.535 108.885 ;
      RECT 48.905 108.715 49.075 108.885 ;
      RECT 48.445 108.715 48.615 108.885 ;
      RECT 47.985 108.715 48.155 108.885 ;
      RECT 47.525 108.715 47.695 108.885 ;
      RECT 47.065 108.715 47.235 108.885 ;
      RECT 46.605 108.715 46.775 108.885 ;
      RECT 46.145 108.715 46.315 108.885 ;
      RECT 45.685 108.715 45.855 108.885 ;
      RECT 45.225 108.715 45.395 108.885 ;
      RECT 44.765 108.715 44.935 108.885 ;
      RECT 44.305 108.715 44.475 108.885 ;
      RECT 43.845 108.715 44.015 108.885 ;
      RECT 43.385 108.715 43.555 108.885 ;
      RECT 42.925 108.715 43.095 108.885 ;
      RECT 42.465 108.715 42.635 108.885 ;
      RECT 42.005 108.715 42.175 108.885 ;
      RECT 41.545 108.715 41.715 108.885 ;
      RECT 41.085 108.715 41.255 108.885 ;
      RECT 40.625 108.715 40.795 108.885 ;
      RECT 40.165 108.715 40.335 108.885 ;
      RECT 39.705 108.715 39.875 108.885 ;
      RECT 39.245 108.715 39.415 108.885 ;
      RECT 38.785 108.715 38.955 108.885 ;
      RECT 38.325 108.715 38.495 108.885 ;
      RECT 37.865 108.715 38.035 108.885 ;
      RECT 37.405 108.715 37.575 108.885 ;
      RECT 36.945 108.715 37.115 108.885 ;
      RECT 36.485 108.715 36.655 108.885 ;
      RECT 36.025 108.715 36.195 108.885 ;
      RECT 35.565 108.715 35.735 108.885 ;
      RECT 35.105 108.715 35.275 108.885 ;
      RECT 34.645 108.715 34.815 108.885 ;
      RECT 34.185 108.715 34.355 108.885 ;
      RECT 33.725 108.715 33.895 108.885 ;
      RECT 33.265 108.715 33.435 108.885 ;
      RECT 32.805 108.715 32.975 108.885 ;
      RECT 32.345 108.715 32.515 108.885 ;
      RECT 31.885 108.715 32.055 108.885 ;
      RECT 31.425 108.715 31.595 108.885 ;
      RECT 30.965 108.715 31.135 108.885 ;
      RECT 30.505 108.715 30.675 108.885 ;
      RECT 30.045 108.715 30.215 108.885 ;
      RECT 29.585 108.715 29.755 108.885 ;
      RECT 29.125 108.715 29.295 108.885 ;
      RECT 28.665 108.715 28.835 108.885 ;
      RECT 28.205 108.715 28.375 108.885 ;
      RECT 27.745 108.715 27.915 108.885 ;
      RECT 27.285 108.715 27.455 108.885 ;
      RECT 26.825 108.715 26.995 108.885 ;
      RECT 26.365 108.715 26.535 108.885 ;
      RECT 25.905 108.715 26.075 108.885 ;
      RECT 91.685 105.995 91.855 106.165 ;
      RECT 91.225 105.995 91.395 106.165 ;
      RECT 26.365 105.995 26.535 106.165 ;
      RECT 25.905 105.995 26.075 106.165 ;
      RECT 91.685 103.275 91.855 103.445 ;
      RECT 91.225 103.275 91.395 103.445 ;
      RECT 26.365 103.275 26.535 103.445 ;
      RECT 25.905 103.275 26.075 103.445 ;
      RECT 91.685 100.555 91.855 100.725 ;
      RECT 91.225 100.555 91.395 100.725 ;
      RECT 26.365 100.555 26.535 100.725 ;
      RECT 25.905 100.555 26.075 100.725 ;
      RECT 117.445 97.835 117.615 98.005 ;
      RECT 116.985 97.835 117.155 98.005 ;
      RECT 116.525 97.835 116.695 98.005 ;
      RECT 116.065 97.835 116.235 98.005 ;
      RECT 115.605 97.835 115.775 98.005 ;
      RECT 115.145 97.835 115.315 98.005 ;
      RECT 114.685 97.835 114.855 98.005 ;
      RECT 114.225 97.835 114.395 98.005 ;
      RECT 113.765 97.835 113.935 98.005 ;
      RECT 113.305 97.835 113.475 98.005 ;
      RECT 112.845 97.835 113.015 98.005 ;
      RECT 112.385 97.835 112.555 98.005 ;
      RECT 111.925 97.835 112.095 98.005 ;
      RECT 111.465 97.835 111.635 98.005 ;
      RECT 111.005 97.835 111.175 98.005 ;
      RECT 110.545 97.835 110.715 98.005 ;
      RECT 110.085 97.835 110.255 98.005 ;
      RECT 109.625 97.835 109.795 98.005 ;
      RECT 109.165 97.835 109.335 98.005 ;
      RECT 108.705 97.835 108.875 98.005 ;
      RECT 108.245 97.835 108.415 98.005 ;
      RECT 107.785 97.835 107.955 98.005 ;
      RECT 107.325 97.835 107.495 98.005 ;
      RECT 106.865 97.835 107.035 98.005 ;
      RECT 106.405 97.835 106.575 98.005 ;
      RECT 105.945 97.835 106.115 98.005 ;
      RECT 105.485 97.835 105.655 98.005 ;
      RECT 105.025 97.835 105.195 98.005 ;
      RECT 104.565 97.835 104.735 98.005 ;
      RECT 104.105 97.835 104.275 98.005 ;
      RECT 103.645 97.835 103.815 98.005 ;
      RECT 103.185 97.835 103.355 98.005 ;
      RECT 102.725 97.835 102.895 98.005 ;
      RECT 102.265 97.835 102.435 98.005 ;
      RECT 101.805 97.835 101.975 98.005 ;
      RECT 101.345 97.835 101.515 98.005 ;
      RECT 100.885 97.835 101.055 98.005 ;
      RECT 100.425 97.835 100.595 98.005 ;
      RECT 99.965 97.835 100.135 98.005 ;
      RECT 99.505 97.835 99.675 98.005 ;
      RECT 99.045 97.835 99.215 98.005 ;
      RECT 98.585 97.835 98.755 98.005 ;
      RECT 98.125 97.835 98.295 98.005 ;
      RECT 97.665 97.835 97.835 98.005 ;
      RECT 97.205 97.835 97.375 98.005 ;
      RECT 96.745 97.835 96.915 98.005 ;
      RECT 96.285 97.835 96.455 98.005 ;
      RECT 95.825 97.835 95.995 98.005 ;
      RECT 95.365 97.835 95.535 98.005 ;
      RECT 94.905 97.835 95.075 98.005 ;
      RECT 94.445 97.835 94.615 98.005 ;
      RECT 93.985 97.835 94.155 98.005 ;
      RECT 93.525 97.835 93.695 98.005 ;
      RECT 93.065 97.835 93.235 98.005 ;
      RECT 92.605 97.835 92.775 98.005 ;
      RECT 92.145 97.835 92.315 98.005 ;
      RECT 91.685 97.835 91.855 98.005 ;
      RECT 91.225 97.835 91.395 98.005 ;
      RECT 90.765 97.835 90.935 98.005 ;
      RECT 90.305 97.835 90.475 98.005 ;
      RECT 89.845 97.835 90.015 98.005 ;
      RECT 89.385 97.835 89.555 98.005 ;
      RECT 88.925 97.835 89.095 98.005 ;
      RECT 88.465 97.835 88.635 98.005 ;
      RECT 88.005 97.835 88.175 98.005 ;
      RECT 87.545 97.835 87.715 98.005 ;
      RECT 87.085 97.835 87.255 98.005 ;
      RECT 86.625 97.835 86.795 98.005 ;
      RECT 86.165 97.835 86.335 98.005 ;
      RECT 85.705 97.835 85.875 98.005 ;
      RECT 85.245 97.835 85.415 98.005 ;
      RECT 84.785 97.835 84.955 98.005 ;
      RECT 84.325 97.835 84.495 98.005 ;
      RECT 83.865 97.835 84.035 98.005 ;
      RECT 83.405 97.835 83.575 98.005 ;
      RECT 82.945 97.835 83.115 98.005 ;
      RECT 82.485 97.835 82.655 98.005 ;
      RECT 82.025 97.835 82.195 98.005 ;
      RECT 81.565 97.835 81.735 98.005 ;
      RECT 81.105 97.835 81.275 98.005 ;
      RECT 80.645 97.835 80.815 98.005 ;
      RECT 80.185 97.835 80.355 98.005 ;
      RECT 79.725 97.835 79.895 98.005 ;
      RECT 79.265 97.835 79.435 98.005 ;
      RECT 78.805 97.835 78.975 98.005 ;
      RECT 78.345 97.835 78.515 98.005 ;
      RECT 77.885 97.835 78.055 98.005 ;
      RECT 77.425 97.835 77.595 98.005 ;
      RECT 76.965 97.835 77.135 98.005 ;
      RECT 76.505 97.835 76.675 98.005 ;
      RECT 76.045 97.835 76.215 98.005 ;
      RECT 75.585 97.835 75.755 98.005 ;
      RECT 75.125 97.835 75.295 98.005 ;
      RECT 74.665 97.835 74.835 98.005 ;
      RECT 74.205 97.835 74.375 98.005 ;
      RECT 73.745 97.835 73.915 98.005 ;
      RECT 73.285 97.835 73.455 98.005 ;
      RECT 72.825 97.835 72.995 98.005 ;
      RECT 72.365 97.835 72.535 98.005 ;
      RECT 71.905 97.835 72.075 98.005 ;
      RECT 71.445 97.835 71.615 98.005 ;
      RECT 70.985 97.835 71.155 98.005 ;
      RECT 70.525 97.835 70.695 98.005 ;
      RECT 70.065 97.835 70.235 98.005 ;
      RECT 69.605 97.835 69.775 98.005 ;
      RECT 69.145 97.835 69.315 98.005 ;
      RECT 68.685 97.835 68.855 98.005 ;
      RECT 68.225 97.835 68.395 98.005 ;
      RECT 67.765 97.835 67.935 98.005 ;
      RECT 67.305 97.835 67.475 98.005 ;
      RECT 66.845 97.835 67.015 98.005 ;
      RECT 66.385 97.835 66.555 98.005 ;
      RECT 65.925 97.835 66.095 98.005 ;
      RECT 65.465 97.835 65.635 98.005 ;
      RECT 65.005 97.835 65.175 98.005 ;
      RECT 64.545 97.835 64.715 98.005 ;
      RECT 64.085 97.835 64.255 98.005 ;
      RECT 63.625 97.835 63.795 98.005 ;
      RECT 63.165 97.835 63.335 98.005 ;
      RECT 62.705 97.835 62.875 98.005 ;
      RECT 62.245 97.835 62.415 98.005 ;
      RECT 61.785 97.835 61.955 98.005 ;
      RECT 61.325 97.835 61.495 98.005 ;
      RECT 60.865 97.835 61.035 98.005 ;
      RECT 60.405 97.835 60.575 98.005 ;
      RECT 59.945 97.835 60.115 98.005 ;
      RECT 59.485 97.835 59.655 98.005 ;
      RECT 59.025 97.835 59.195 98.005 ;
      RECT 58.565 97.835 58.735 98.005 ;
      RECT 58.105 97.835 58.275 98.005 ;
      RECT 57.645 97.835 57.815 98.005 ;
      RECT 57.185 97.835 57.355 98.005 ;
      RECT 56.725 97.835 56.895 98.005 ;
      RECT 56.265 97.835 56.435 98.005 ;
      RECT 55.805 97.835 55.975 98.005 ;
      RECT 55.345 97.835 55.515 98.005 ;
      RECT 54.885 97.835 55.055 98.005 ;
      RECT 54.425 97.835 54.595 98.005 ;
      RECT 53.965 97.835 54.135 98.005 ;
      RECT 53.505 97.835 53.675 98.005 ;
      RECT 53.045 97.835 53.215 98.005 ;
      RECT 52.585 97.835 52.755 98.005 ;
      RECT 52.125 97.835 52.295 98.005 ;
      RECT 51.665 97.835 51.835 98.005 ;
      RECT 51.205 97.835 51.375 98.005 ;
      RECT 50.745 97.835 50.915 98.005 ;
      RECT 50.285 97.835 50.455 98.005 ;
      RECT 49.825 97.835 49.995 98.005 ;
      RECT 49.365 97.835 49.535 98.005 ;
      RECT 48.905 97.835 49.075 98.005 ;
      RECT 48.445 97.835 48.615 98.005 ;
      RECT 47.985 97.835 48.155 98.005 ;
      RECT 47.525 97.835 47.695 98.005 ;
      RECT 47.065 97.835 47.235 98.005 ;
      RECT 46.605 97.835 46.775 98.005 ;
      RECT 46.145 97.835 46.315 98.005 ;
      RECT 45.685 97.835 45.855 98.005 ;
      RECT 45.225 97.835 45.395 98.005 ;
      RECT 44.765 97.835 44.935 98.005 ;
      RECT 44.305 97.835 44.475 98.005 ;
      RECT 43.845 97.835 44.015 98.005 ;
      RECT 43.385 97.835 43.555 98.005 ;
      RECT 42.925 97.835 43.095 98.005 ;
      RECT 42.465 97.835 42.635 98.005 ;
      RECT 42.005 97.835 42.175 98.005 ;
      RECT 41.545 97.835 41.715 98.005 ;
      RECT 41.085 97.835 41.255 98.005 ;
      RECT 40.625 97.835 40.795 98.005 ;
      RECT 40.165 97.835 40.335 98.005 ;
      RECT 39.705 97.835 39.875 98.005 ;
      RECT 39.245 97.835 39.415 98.005 ;
      RECT 38.785 97.835 38.955 98.005 ;
      RECT 38.325 97.835 38.495 98.005 ;
      RECT 37.865 97.835 38.035 98.005 ;
      RECT 37.405 97.835 37.575 98.005 ;
      RECT 36.945 97.835 37.115 98.005 ;
      RECT 36.485 97.835 36.655 98.005 ;
      RECT 36.025 97.835 36.195 98.005 ;
      RECT 35.565 97.835 35.735 98.005 ;
      RECT 35.105 97.835 35.275 98.005 ;
      RECT 34.645 97.835 34.815 98.005 ;
      RECT 34.185 97.835 34.355 98.005 ;
      RECT 33.725 97.835 33.895 98.005 ;
      RECT 33.265 97.835 33.435 98.005 ;
      RECT 32.805 97.835 32.975 98.005 ;
      RECT 32.345 97.835 32.515 98.005 ;
      RECT 31.885 97.835 32.055 98.005 ;
      RECT 31.425 97.835 31.595 98.005 ;
      RECT 30.965 97.835 31.135 98.005 ;
      RECT 30.505 97.835 30.675 98.005 ;
      RECT 30.045 97.835 30.215 98.005 ;
      RECT 29.585 97.835 29.755 98.005 ;
      RECT 29.125 97.835 29.295 98.005 ;
      RECT 28.665 97.835 28.835 98.005 ;
      RECT 28.205 97.835 28.375 98.005 ;
      RECT 27.745 97.835 27.915 98.005 ;
      RECT 27.285 97.835 27.455 98.005 ;
      RECT 26.825 97.835 26.995 98.005 ;
      RECT 26.365 97.835 26.535 98.005 ;
      RECT 25.905 97.835 26.075 98.005 ;
      RECT 25.445 97.835 25.615 98.005 ;
      RECT 24.985 97.835 25.155 98.005 ;
      RECT 24.525 97.835 24.695 98.005 ;
      RECT 24.065 97.835 24.235 98.005 ;
      RECT 23.605 97.835 23.775 98.005 ;
      RECT 23.145 97.835 23.315 98.005 ;
      RECT 22.685 97.835 22.855 98.005 ;
      RECT 22.225 97.835 22.395 98.005 ;
      RECT 21.765 97.835 21.935 98.005 ;
      RECT 21.305 97.835 21.475 98.005 ;
      RECT 20.845 97.835 21.015 98.005 ;
      RECT 20.385 97.835 20.555 98.005 ;
      RECT 19.925 97.835 20.095 98.005 ;
      RECT 19.465 97.835 19.635 98.005 ;
      RECT 19.005 97.835 19.175 98.005 ;
      RECT 18.545 97.835 18.715 98.005 ;
      RECT 18.085 97.835 18.255 98.005 ;
      RECT 17.625 97.835 17.795 98.005 ;
      RECT 17.165 97.835 17.335 98.005 ;
      RECT 16.705 97.835 16.875 98.005 ;
      RECT 16.245 97.835 16.415 98.005 ;
      RECT 15.785 97.835 15.955 98.005 ;
      RECT 15.325 97.835 15.495 98.005 ;
      RECT 14.865 97.835 15.035 98.005 ;
      RECT 14.405 97.835 14.575 98.005 ;
      RECT 13.945 97.835 14.115 98.005 ;
      RECT 13.485 97.835 13.655 98.005 ;
      RECT 13.025 97.835 13.195 98.005 ;
      RECT 12.565 97.835 12.735 98.005 ;
      RECT 12.105 97.835 12.275 98.005 ;
      RECT 11.645 97.835 11.815 98.005 ;
      RECT 11.185 97.835 11.355 98.005 ;
      RECT 10.725 97.835 10.895 98.005 ;
      RECT 10.265 97.835 10.435 98.005 ;
      RECT 9.805 97.835 9.975 98.005 ;
      RECT 9.345 97.835 9.515 98.005 ;
      RECT 8.885 97.835 9.055 98.005 ;
      RECT 8.425 97.835 8.595 98.005 ;
      RECT 7.965 97.835 8.135 98.005 ;
      RECT 7.505 97.835 7.675 98.005 ;
      RECT 7.045 97.835 7.215 98.005 ;
      RECT 6.585 97.835 6.755 98.005 ;
      RECT 6.125 97.835 6.295 98.005 ;
      RECT 5.665 97.835 5.835 98.005 ;
      RECT 5.205 97.835 5.375 98.005 ;
      RECT 4.745 97.835 4.915 98.005 ;
      RECT 4.285 97.835 4.455 98.005 ;
      RECT 3.825 97.835 3.995 98.005 ;
      RECT 3.365 97.835 3.535 98.005 ;
      RECT 2.905 97.835 3.075 98.005 ;
      RECT 2.445 97.835 2.615 98.005 ;
      RECT 1.985 97.835 2.155 98.005 ;
      RECT 1.525 97.835 1.695 98.005 ;
      RECT 1.065 97.835 1.235 98.005 ;
      RECT 0.605 97.835 0.775 98.005 ;
      RECT 0.145 97.835 0.315 98.005 ;
      RECT 117.445 95.115 117.615 95.285 ;
      RECT 116.985 95.115 117.155 95.285 ;
      RECT 0.605 95.115 0.775 95.285 ;
      RECT 0.145 95.115 0.315 95.285 ;
      RECT 117.445 92.395 117.615 92.565 ;
      RECT 116.985 92.395 117.155 92.565 ;
      RECT 0.605 92.395 0.775 92.565 ;
      RECT 0.145 92.395 0.315 92.565 ;
      RECT 117.445 89.675 117.615 89.845 ;
      RECT 116.985 89.675 117.155 89.845 ;
      RECT 0.605 89.675 0.775 89.845 ;
      RECT 0.145 89.675 0.315 89.845 ;
      RECT 117.445 86.955 117.615 87.125 ;
      RECT 116.985 86.955 117.155 87.125 ;
      RECT 0.605 86.955 0.775 87.125 ;
      RECT 0.145 86.955 0.315 87.125 ;
      RECT 117.445 84.235 117.615 84.405 ;
      RECT 116.985 84.235 117.155 84.405 ;
      RECT 0.605 84.235 0.775 84.405 ;
      RECT 0.145 84.235 0.315 84.405 ;
      RECT 117.445 81.515 117.615 81.685 ;
      RECT 116.985 81.515 117.155 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 117.445 78.795 117.615 78.965 ;
      RECT 116.985 78.795 117.155 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 117.445 76.075 117.615 76.245 ;
      RECT 116.985 76.075 117.155 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 117.445 73.355 117.615 73.525 ;
      RECT 116.985 73.355 117.155 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 117.445 70.635 117.615 70.805 ;
      RECT 116.985 70.635 117.155 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 117.445 67.915 117.615 68.085 ;
      RECT 116.985 67.915 117.155 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 117.445 65.195 117.615 65.365 ;
      RECT 116.985 65.195 117.155 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 117.445 62.475 117.615 62.645 ;
      RECT 116.985 62.475 117.155 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 117.445 59.755 117.615 59.925 ;
      RECT 116.985 59.755 117.155 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 117.445 57.035 117.615 57.205 ;
      RECT 116.985 57.035 117.155 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 117.445 54.315 117.615 54.485 ;
      RECT 116.985 54.315 117.155 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 117.445 51.595 117.615 51.765 ;
      RECT 116.985 51.595 117.155 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 117.445 48.875 117.615 49.045 ;
      RECT 116.985 48.875 117.155 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 117.445 46.155 117.615 46.325 ;
      RECT 116.985 46.155 117.155 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 117.445 43.435 117.615 43.605 ;
      RECT 116.985 43.435 117.155 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 117.445 40.715 117.615 40.885 ;
      RECT 116.985 40.715 117.155 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 117.445 37.995 117.615 38.165 ;
      RECT 116.985 37.995 117.155 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 117.445 35.275 117.615 35.445 ;
      RECT 116.985 35.275 117.155 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 117.445 32.555 117.615 32.725 ;
      RECT 116.985 32.555 117.155 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 117.445 29.835 117.615 30.005 ;
      RECT 116.985 29.835 117.155 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 117.445 27.115 117.615 27.285 ;
      RECT 116.985 27.115 117.155 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 117.445 24.395 117.615 24.565 ;
      RECT 116.985 24.395 117.155 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 117.445 21.675 117.615 21.845 ;
      RECT 116.985 21.675 117.155 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 117.445 18.955 117.615 19.125 ;
      RECT 116.985 18.955 117.155 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 117.445 16.235 117.615 16.405 ;
      RECT 116.985 16.235 117.155 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 117.445 13.515 117.615 13.685 ;
      RECT 116.985 13.515 117.155 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 117.445 10.795 117.615 10.965 ;
      RECT 116.985 10.795 117.155 10.965 ;
      RECT 116.525 10.795 116.695 10.965 ;
      RECT 116.065 10.795 116.235 10.965 ;
      RECT 115.605 10.795 115.775 10.965 ;
      RECT 115.145 10.795 115.315 10.965 ;
      RECT 114.685 10.795 114.855 10.965 ;
      RECT 114.225 10.795 114.395 10.965 ;
      RECT 113.765 10.795 113.935 10.965 ;
      RECT 113.305 10.795 113.475 10.965 ;
      RECT 112.845 10.795 113.015 10.965 ;
      RECT 112.385 10.795 112.555 10.965 ;
      RECT 111.925 10.795 112.095 10.965 ;
      RECT 111.465 10.795 111.635 10.965 ;
      RECT 111.005 10.795 111.175 10.965 ;
      RECT 110.545 10.795 110.715 10.965 ;
      RECT 110.085 10.795 110.255 10.965 ;
      RECT 109.625 10.795 109.795 10.965 ;
      RECT 109.165 10.795 109.335 10.965 ;
      RECT 108.705 10.795 108.875 10.965 ;
      RECT 108.245 10.795 108.415 10.965 ;
      RECT 107.785 10.795 107.955 10.965 ;
      RECT 107.325 10.795 107.495 10.965 ;
      RECT 106.865 10.795 107.035 10.965 ;
      RECT 106.405 10.795 106.575 10.965 ;
      RECT 105.945 10.795 106.115 10.965 ;
      RECT 105.485 10.795 105.655 10.965 ;
      RECT 105.025 10.795 105.195 10.965 ;
      RECT 104.565 10.795 104.735 10.965 ;
      RECT 104.105 10.795 104.275 10.965 ;
      RECT 103.645 10.795 103.815 10.965 ;
      RECT 103.185 10.795 103.355 10.965 ;
      RECT 102.725 10.795 102.895 10.965 ;
      RECT 102.265 10.795 102.435 10.965 ;
      RECT 101.805 10.795 101.975 10.965 ;
      RECT 101.345 10.795 101.515 10.965 ;
      RECT 100.885 10.795 101.055 10.965 ;
      RECT 100.425 10.795 100.595 10.965 ;
      RECT 99.965 10.795 100.135 10.965 ;
      RECT 99.505 10.795 99.675 10.965 ;
      RECT 99.045 10.795 99.215 10.965 ;
      RECT 98.585 10.795 98.755 10.965 ;
      RECT 98.125 10.795 98.295 10.965 ;
      RECT 97.665 10.795 97.835 10.965 ;
      RECT 97.205 10.795 97.375 10.965 ;
      RECT 96.745 10.795 96.915 10.965 ;
      RECT 96.285 10.795 96.455 10.965 ;
      RECT 95.825 10.795 95.995 10.965 ;
      RECT 95.365 10.795 95.535 10.965 ;
      RECT 94.905 10.795 95.075 10.965 ;
      RECT 94.445 10.795 94.615 10.965 ;
      RECT 93.985 10.795 94.155 10.965 ;
      RECT 93.525 10.795 93.695 10.965 ;
      RECT 93.065 10.795 93.235 10.965 ;
      RECT 92.605 10.795 92.775 10.965 ;
      RECT 92.145 10.795 92.315 10.965 ;
      RECT 91.685 10.795 91.855 10.965 ;
      RECT 91.225 10.795 91.395 10.965 ;
      RECT 90.765 10.795 90.935 10.965 ;
      RECT 90.305 10.795 90.475 10.965 ;
      RECT 89.845 10.795 90.015 10.965 ;
      RECT 89.385 10.795 89.555 10.965 ;
      RECT 88.925 10.795 89.095 10.965 ;
      RECT 88.465 10.795 88.635 10.965 ;
      RECT 88.005 10.795 88.175 10.965 ;
      RECT 87.545 10.795 87.715 10.965 ;
      RECT 87.085 10.795 87.255 10.965 ;
      RECT 86.625 10.795 86.795 10.965 ;
      RECT 86.165 10.795 86.335 10.965 ;
      RECT 85.705 10.795 85.875 10.965 ;
      RECT 85.245 10.795 85.415 10.965 ;
      RECT 84.785 10.795 84.955 10.965 ;
      RECT 84.325 10.795 84.495 10.965 ;
      RECT 83.865 10.795 84.035 10.965 ;
      RECT 83.405 10.795 83.575 10.965 ;
      RECT 82.945 10.795 83.115 10.965 ;
      RECT 82.485 10.795 82.655 10.965 ;
      RECT 82.025 10.795 82.195 10.965 ;
      RECT 81.565 10.795 81.735 10.965 ;
      RECT 81.105 10.795 81.275 10.965 ;
      RECT 80.645 10.795 80.815 10.965 ;
      RECT 80.185 10.795 80.355 10.965 ;
      RECT 79.725 10.795 79.895 10.965 ;
      RECT 79.265 10.795 79.435 10.965 ;
      RECT 78.805 10.795 78.975 10.965 ;
      RECT 78.345 10.795 78.515 10.965 ;
      RECT 77.885 10.795 78.055 10.965 ;
      RECT 77.425 10.795 77.595 10.965 ;
      RECT 76.965 10.795 77.135 10.965 ;
      RECT 76.505 10.795 76.675 10.965 ;
      RECT 76.045 10.795 76.215 10.965 ;
      RECT 75.585 10.795 75.755 10.965 ;
      RECT 75.125 10.795 75.295 10.965 ;
      RECT 74.665 10.795 74.835 10.965 ;
      RECT 74.205 10.795 74.375 10.965 ;
      RECT 73.745 10.795 73.915 10.965 ;
      RECT 73.285 10.795 73.455 10.965 ;
      RECT 72.825 10.795 72.995 10.965 ;
      RECT 72.365 10.795 72.535 10.965 ;
      RECT 71.905 10.795 72.075 10.965 ;
      RECT 71.445 10.795 71.615 10.965 ;
      RECT 70.985 10.795 71.155 10.965 ;
      RECT 70.525 10.795 70.695 10.965 ;
      RECT 70.065 10.795 70.235 10.965 ;
      RECT 69.605 10.795 69.775 10.965 ;
      RECT 69.145 10.795 69.315 10.965 ;
      RECT 68.685 10.795 68.855 10.965 ;
      RECT 68.225 10.795 68.395 10.965 ;
      RECT 67.765 10.795 67.935 10.965 ;
      RECT 67.305 10.795 67.475 10.965 ;
      RECT 66.845 10.795 67.015 10.965 ;
      RECT 66.385 10.795 66.555 10.965 ;
      RECT 65.925 10.795 66.095 10.965 ;
      RECT 65.465 10.795 65.635 10.965 ;
      RECT 65.005 10.795 65.175 10.965 ;
      RECT 64.545 10.795 64.715 10.965 ;
      RECT 64.085 10.795 64.255 10.965 ;
      RECT 63.625 10.795 63.795 10.965 ;
      RECT 63.165 10.795 63.335 10.965 ;
      RECT 62.705 10.795 62.875 10.965 ;
      RECT 62.245 10.795 62.415 10.965 ;
      RECT 61.785 10.795 61.955 10.965 ;
      RECT 61.325 10.795 61.495 10.965 ;
      RECT 60.865 10.795 61.035 10.965 ;
      RECT 60.405 10.795 60.575 10.965 ;
      RECT 59.945 10.795 60.115 10.965 ;
      RECT 59.485 10.795 59.655 10.965 ;
      RECT 59.025 10.795 59.195 10.965 ;
      RECT 58.565 10.795 58.735 10.965 ;
      RECT 58.105 10.795 58.275 10.965 ;
      RECT 57.645 10.795 57.815 10.965 ;
      RECT 57.185 10.795 57.355 10.965 ;
      RECT 56.725 10.795 56.895 10.965 ;
      RECT 56.265 10.795 56.435 10.965 ;
      RECT 55.805 10.795 55.975 10.965 ;
      RECT 55.345 10.795 55.515 10.965 ;
      RECT 54.885 10.795 55.055 10.965 ;
      RECT 54.425 10.795 54.595 10.965 ;
      RECT 53.965 10.795 54.135 10.965 ;
      RECT 53.505 10.795 53.675 10.965 ;
      RECT 53.045 10.795 53.215 10.965 ;
      RECT 52.585 10.795 52.755 10.965 ;
      RECT 52.125 10.795 52.295 10.965 ;
      RECT 51.665 10.795 51.835 10.965 ;
      RECT 51.205 10.795 51.375 10.965 ;
      RECT 50.745 10.795 50.915 10.965 ;
      RECT 50.285 10.795 50.455 10.965 ;
      RECT 49.825 10.795 49.995 10.965 ;
      RECT 49.365 10.795 49.535 10.965 ;
      RECT 48.905 10.795 49.075 10.965 ;
      RECT 48.445 10.795 48.615 10.965 ;
      RECT 47.985 10.795 48.155 10.965 ;
      RECT 47.525 10.795 47.695 10.965 ;
      RECT 47.065 10.795 47.235 10.965 ;
      RECT 46.605 10.795 46.775 10.965 ;
      RECT 46.145 10.795 46.315 10.965 ;
      RECT 45.685 10.795 45.855 10.965 ;
      RECT 45.225 10.795 45.395 10.965 ;
      RECT 44.765 10.795 44.935 10.965 ;
      RECT 44.305 10.795 44.475 10.965 ;
      RECT 43.845 10.795 44.015 10.965 ;
      RECT 43.385 10.795 43.555 10.965 ;
      RECT 42.925 10.795 43.095 10.965 ;
      RECT 42.465 10.795 42.635 10.965 ;
      RECT 42.005 10.795 42.175 10.965 ;
      RECT 41.545 10.795 41.715 10.965 ;
      RECT 41.085 10.795 41.255 10.965 ;
      RECT 40.625 10.795 40.795 10.965 ;
      RECT 40.165 10.795 40.335 10.965 ;
      RECT 39.705 10.795 39.875 10.965 ;
      RECT 39.245 10.795 39.415 10.965 ;
      RECT 38.785 10.795 38.955 10.965 ;
      RECT 38.325 10.795 38.495 10.965 ;
      RECT 37.865 10.795 38.035 10.965 ;
      RECT 37.405 10.795 37.575 10.965 ;
      RECT 36.945 10.795 37.115 10.965 ;
      RECT 36.485 10.795 36.655 10.965 ;
      RECT 36.025 10.795 36.195 10.965 ;
      RECT 35.565 10.795 35.735 10.965 ;
      RECT 35.105 10.795 35.275 10.965 ;
      RECT 34.645 10.795 34.815 10.965 ;
      RECT 34.185 10.795 34.355 10.965 ;
      RECT 33.725 10.795 33.895 10.965 ;
      RECT 33.265 10.795 33.435 10.965 ;
      RECT 32.805 10.795 32.975 10.965 ;
      RECT 32.345 10.795 32.515 10.965 ;
      RECT 31.885 10.795 32.055 10.965 ;
      RECT 31.425 10.795 31.595 10.965 ;
      RECT 30.965 10.795 31.135 10.965 ;
      RECT 30.505 10.795 30.675 10.965 ;
      RECT 30.045 10.795 30.215 10.965 ;
      RECT 29.585 10.795 29.755 10.965 ;
      RECT 29.125 10.795 29.295 10.965 ;
      RECT 28.665 10.795 28.835 10.965 ;
      RECT 28.205 10.795 28.375 10.965 ;
      RECT 27.745 10.795 27.915 10.965 ;
      RECT 27.285 10.795 27.455 10.965 ;
      RECT 26.825 10.795 26.995 10.965 ;
      RECT 26.365 10.795 26.535 10.965 ;
      RECT 25.905 10.795 26.075 10.965 ;
      RECT 25.445 10.795 25.615 10.965 ;
      RECT 24.985 10.795 25.155 10.965 ;
      RECT 24.525 10.795 24.695 10.965 ;
      RECT 24.065 10.795 24.235 10.965 ;
      RECT 23.605 10.795 23.775 10.965 ;
      RECT 23.145 10.795 23.315 10.965 ;
      RECT 22.685 10.795 22.855 10.965 ;
      RECT 22.225 10.795 22.395 10.965 ;
      RECT 21.765 10.795 21.935 10.965 ;
      RECT 21.305 10.795 21.475 10.965 ;
      RECT 20.845 10.795 21.015 10.965 ;
      RECT 20.385 10.795 20.555 10.965 ;
      RECT 19.925 10.795 20.095 10.965 ;
      RECT 19.465 10.795 19.635 10.965 ;
      RECT 19.005 10.795 19.175 10.965 ;
      RECT 18.545 10.795 18.715 10.965 ;
      RECT 18.085 10.795 18.255 10.965 ;
      RECT 17.625 10.795 17.795 10.965 ;
      RECT 17.165 10.795 17.335 10.965 ;
      RECT 16.705 10.795 16.875 10.965 ;
      RECT 16.245 10.795 16.415 10.965 ;
      RECT 15.785 10.795 15.955 10.965 ;
      RECT 15.325 10.795 15.495 10.965 ;
      RECT 14.865 10.795 15.035 10.965 ;
      RECT 14.405 10.795 14.575 10.965 ;
      RECT 13.945 10.795 14.115 10.965 ;
      RECT 13.485 10.795 13.655 10.965 ;
      RECT 13.025 10.795 13.195 10.965 ;
      RECT 12.565 10.795 12.735 10.965 ;
      RECT 12.105 10.795 12.275 10.965 ;
      RECT 11.645 10.795 11.815 10.965 ;
      RECT 11.185 10.795 11.355 10.965 ;
      RECT 10.725 10.795 10.895 10.965 ;
      RECT 10.265 10.795 10.435 10.965 ;
      RECT 9.805 10.795 9.975 10.965 ;
      RECT 9.345 10.795 9.515 10.965 ;
      RECT 8.885 10.795 9.055 10.965 ;
      RECT 8.425 10.795 8.595 10.965 ;
      RECT 7.965 10.795 8.135 10.965 ;
      RECT 7.505 10.795 7.675 10.965 ;
      RECT 7.045 10.795 7.215 10.965 ;
      RECT 6.585 10.795 6.755 10.965 ;
      RECT 6.125 10.795 6.295 10.965 ;
      RECT 5.665 10.795 5.835 10.965 ;
      RECT 5.205 10.795 5.375 10.965 ;
      RECT 4.745 10.795 4.915 10.965 ;
      RECT 4.285 10.795 4.455 10.965 ;
      RECT 3.825 10.795 3.995 10.965 ;
      RECT 3.365 10.795 3.535 10.965 ;
      RECT 2.905 10.795 3.075 10.965 ;
      RECT 2.445 10.795 2.615 10.965 ;
      RECT 1.985 10.795 2.155 10.965 ;
      RECT 1.525 10.795 1.695 10.965 ;
      RECT 1.065 10.795 1.235 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 91.685 8.075 91.855 8.245 ;
      RECT 91.225 8.075 91.395 8.245 ;
      RECT 26.365 8.075 26.535 8.245 ;
      RECT 25.905 8.075 26.075 8.245 ;
      RECT 91.685 5.355 91.855 5.525 ;
      RECT 91.225 5.355 91.395 5.525 ;
      RECT 26.365 5.355 26.535 5.525 ;
      RECT 25.905 5.355 26.075 5.525 ;
      RECT 91.685 2.635 91.855 2.805 ;
      RECT 91.225 2.635 91.395 2.805 ;
      RECT 26.365 2.635 26.535 2.805 ;
      RECT 25.905 2.635 26.075 2.805 ;
      RECT 91.685 -0.085 91.855 0.085 ;
      RECT 91.225 -0.085 91.395 0.085 ;
      RECT 90.765 -0.085 90.935 0.085 ;
      RECT 90.305 -0.085 90.475 0.085 ;
      RECT 89.845 -0.085 90.015 0.085 ;
      RECT 89.385 -0.085 89.555 0.085 ;
      RECT 88.925 -0.085 89.095 0.085 ;
      RECT 88.465 -0.085 88.635 0.085 ;
      RECT 88.005 -0.085 88.175 0.085 ;
      RECT 87.545 -0.085 87.715 0.085 ;
      RECT 87.085 -0.085 87.255 0.085 ;
      RECT 86.625 -0.085 86.795 0.085 ;
      RECT 86.165 -0.085 86.335 0.085 ;
      RECT 85.705 -0.085 85.875 0.085 ;
      RECT 85.245 -0.085 85.415 0.085 ;
      RECT 84.785 -0.085 84.955 0.085 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
    LAYER via ;
      RECT 80.885 108.725 81.035 108.875 ;
      RECT 51.445 108.725 51.595 108.875 ;
      RECT 63.865 107.025 64.015 107.175 ;
      RECT 49.605 107.025 49.755 107.175 ;
      RECT 43.625 107.025 43.775 107.175 ;
      RECT 80.885 97.845 81.035 97.995 ;
      RECT 51.445 97.845 51.595 97.995 ;
      RECT 10.965 97.845 11.115 97.995 ;
      RECT 14.185 96.145 14.335 96.295 ;
      RECT 9.125 96.145 9.275 96.295 ;
      RECT 114.005 12.505 114.155 12.655 ;
      RECT 4.985 12.505 5.135 12.655 ;
      RECT 80.885 10.805 81.035 10.955 ;
      RECT 51.445 10.805 51.595 10.955 ;
      RECT 10.965 10.805 11.115 10.955 ;
      RECT 69.845 1.625 69.995 1.775 ;
      RECT 65.245 1.625 65.395 1.775 ;
      RECT 80.885 -0.075 81.035 0.075 ;
      RECT 51.445 -0.075 51.595 0.075 ;
    LAYER via2 ;
      RECT 80.86 108.7 81.06 108.9 ;
      RECT 51.42 108.7 51.62 108.9 ;
      RECT 10.94 97.82 11.14 98.02 ;
      RECT 1.28 85.58 1.48 85.78 ;
      RECT 1.74 80.14 1.94 80.34 ;
      RECT 1.74 61.1 1.94 61.3 ;
      RECT 1.28 59.06 1.48 59.26 ;
      RECT 116.28 54.3 116.48 54.5 ;
      RECT 115.82 47.5 116.02 47.7 ;
      RECT 1.28 33.22 1.48 33.42 ;
      RECT 116.28 31.86 116.48 32.06 ;
      RECT 10.94 10.78 11.14 10.98 ;
      RECT 80.86 -0.1 81.06 0.1 ;
      RECT 51.42 -0.1 51.62 0.1 ;
    LAYER via3 ;
      RECT 80.86 108.7 81.06 108.9 ;
      RECT 51.42 108.7 51.62 108.9 ;
      RECT 10.94 97.82 11.14 98.02 ;
      RECT 1.74 53.62 1.94 53.82 ;
      RECT 115.82 43.42 116.02 43.62 ;
      RECT 10.94 10.78 11.14 10.98 ;
      RECT 80.86 -0.1 81.06 0.1 ;
      RECT 51.42 -0.1 51.62 0.1 ;
    LAYER OVERLAP ;
      POLYGON 25.76 0 25.76 10.88 0 10.88 0 97.92 25.76 97.92 25.76 108.8 92 108.8 92 97.92 117.76 97.92 117.76 10.88 92 10.88 92 0 ;
  END
END sb_1__1_

END LIBRARY
