//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module sky130_fd_sc_hd__inv_2
(
    A,
    Y
);

    input A;
    output Y;

    wire A;
    wire Y;

endmodule

