VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_0__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 103.96 BY 130.56 ;
  SYMMETRY X Y ;
  PIN pReset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 64.36 0.595 64.5 ;
    END
  END pReset[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 19.63 129.76 19.93 130.56 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.7 130.075 68.84 130.56 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.36 130.075 55.5 130.56 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.74 130.075 10.88 130.56 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.98 130.075 8.12 130.56 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5 130.075 59.64 130.56 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.66 130.075 11.8 130.56 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.5 130.075 13.64 130.56 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.46 130.075 25.6 130.56 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.54 130.075 24.68 130.56 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.5 130.075 36.64 130.56 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 130.075 61.48 130.56 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.06 130.075 53.2 130.56 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.86 130.075 67 130.56 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.08 130.075 70.22 130.56 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.2 130.075 57.34 130.56 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.42 130.075 60.56 130.56 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.3 130.075 27.44 130.56 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 130.075 35.72 130.56 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 130.075 65.16 130.56 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.94 130.075 66.08 130.56 ;
    END
  END chany_top_in[20]
  PIN chany_top_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.12 130.075 58.26 130.56 ;
    END
  END chany_top_in[21]
  PIN chany_top_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.58 130.075 12.72 130.56 ;
    END
  END chany_top_in[22]
  PIN chany_top_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.42 130.075 14.56 130.56 ;
    END
  END chany_top_in[23]
  PIN chany_top_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.06 130.075 30.2 130.56 ;
    END
  END chany_top_in[24]
  PIN chany_top_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.82 130.075 9.96 130.56 ;
    END
  END chany_top_in[25]
  PIN chany_top_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 130.075 64.24 130.56 ;
    END
  END chany_top_in[26]
  PIN chany_top_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 130.075 56.42 130.56 ;
    END
  END chany_top_in[27]
  PIN chany_top_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71 130.075 71.14 130.56 ;
    END
  END chany_top_in[28]
  PIN chany_top_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.54 130.075 47.68 130.56 ;
    END
  END chany_top_in[29]
  PIN top_left_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.84 130.075 3.98 130.56 ;
    END
  END top_left_grid_pin_1_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 47.11 103.96 47.41 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 60.71 103.96 61.01 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 67.51 103.96 67.81 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 45.75 103.96 46.05 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 37.16 103.96 37.3 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 34.1 103.96 34.24 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 52.46 103.96 52.6 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 44.39 103.96 44.69 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 59.35 103.96 59.65 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 26.71 103.96 27.01 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 15.4 103.96 15.54 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 44.64 103.96 44.78 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 58.24 103.96 58.38 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 64.79 103.96 65.09 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 42.6 103.96 42.74 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 50.42 103.96 50.56 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 14.72 103.96 14.86 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 39.88 103.96 40.02 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 41.92 103.96 42.06 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 62.07 103.96 62.37 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 33.42 103.96 33.56 ;
    END
  END chanx_right_in[20]
  PIN chanx_right_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 23.99 103.96 24.29 ;
    END
  END chanx_right_in[21]
  PIN chanx_right_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 47.02 103.96 47.16 ;
    END
  END chanx_right_in[22]
  PIN chanx_right_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 45.32 103.96 45.46 ;
    END
  END chanx_right_in[23]
  PIN chanx_right_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 63.68 103.96 63.82 ;
    END
  END chanx_right_in[24]
  PIN chanx_right_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 49.74 103.96 49.88 ;
    END
  END chanx_right_in[25]
  PIN chanx_right_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 39.2 103.96 39.34 ;
    END
  END chanx_right_in[26]
  PIN chanx_right_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 21.27 103.96 21.57 ;
    END
  END chanx_right_in[27]
  PIN chanx_right_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 36.48 103.96 36.62 ;
    END
  END chanx_right_in[28]
  PIN chanx_right_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 47.7 103.96 47.84 ;
    END
  END chanx_right_in[29]
  PIN right_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94 5.44 94.14 5.925 ;
    END
  END right_bottom_grid_pin_36_[0]
  PIN right_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.76 5.44 96.9 5.925 ;
    END
  END right_bottom_grid_pin_37_[0]
  PIN right_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.84 5.44 95.98 5.925 ;
    END
  END right_bottom_grid_pin_38_[0]
  PIN right_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.92 5.44 95.06 5.925 ;
    END
  END right_bottom_grid_pin_39_[0]
  PIN right_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.4 5.44 89.54 5.925 ;
    END
  END right_bottom_grid_pin_40_[0]
  PIN right_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.32 5.44 90.46 5.925 ;
    END
  END right_bottom_grid_pin_41_[0]
  PIN right_bottom_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.08 5.44 93.22 5.925 ;
    END
  END right_bottom_grid_pin_42_[0]
  PIN right_bottom_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.24 5.44 91.38 5.925 ;
    END
  END right_bottom_grid_pin_43_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.82 0 32.96 0.485 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5 0 59.64 0.485 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.94 0 66.08 0.485 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 0 35.72 0.485 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 0 39.4 0.485 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.86 0 67 0.485 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.74 0 33.88 0.485 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.44 0 54.58 0.485 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.54 0 47.68 0.485 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 0 61.48 0.485 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.82 0 9.96 0.485 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.98 0 8.12 0.485 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.46 0 48.6 0.485 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.12 0 58.26 0.485 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.42 0 60.56 0.485 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.7 0 68.84 0.485 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71 0 71.14 0.485 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.84 0 3.98 0.485 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.66 0 34.8 0.485 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.78 0 44.92 0.485 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.36 0 55.5 0.485 ;
    END
  END chany_bottom_in[20]
  PIN chany_bottom_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.78 0 67.92 0.485 ;
    END
  END chany_bottom_in[21]
  PIN chany_bottom_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 0 56.42 0.485 ;
    END
  END chany_bottom_in[22]
  PIN chany_bottom_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.42 0 37.56 0.485 ;
    END
  END chany_bottom_in[23]
  PIN chany_bottom_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.9 0 9.04 0.485 ;
    END
  END chany_bottom_in[24]
  PIN chany_bottom_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.2 0 57.34 0.485 ;
    END
  END chany_bottom_in[25]
  PIN chany_bottom_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.5 0 36.64 0.485 ;
    END
  END chany_bottom_in[26]
  PIN chany_bottom_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.62 0 46.76 0.485 ;
    END
  END chany_bottom_in[27]
  PIN chany_bottom_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.52 0 53.66 0.485 ;
    END
  END chany_bottom_in[28]
  PIN chany_bottom_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 0 65.16 0.485 ;
    END
  END chany_bottom_in[29]
  PIN bottom_left_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.06 0 7.2 0.485 ;
    END
  END bottom_left_grid_pin_1_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 66.4 103.96 66.54 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.34 130.075 15.48 130.56 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 130.075 62.4 130.56 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.26 130.075 16.4 130.56 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.06 130.075 7.2 130.56 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.62 130.075 46.76 130.56 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.62 130.075 23.76 130.56 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.9 130.075 9.04 130.56 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.42 130.075 37.56 130.56 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.18 130.075 63.32 130.56 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.18 130.075 17.32 130.56 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.7 130.075 45.84 130.56 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.7 130.075 22.84 130.56 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.38 130.075 26.52 130.56 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.1 130.075 18.24 130.56 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.78 130.075 67.92 130.56 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 130.075 38.48 130.56 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.78 130.075 44.92 130.56 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.78 130.075 21.92 130.56 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.76 130.075 4.9 130.56 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 130.075 39.4 130.56 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.86 130.075 44 130.56 ;
    END
  END chany_top_out[20]
  PIN chany_top_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.02 130.075 19.16 130.56 ;
    END
  END chany_top_out[21]
  PIN chany_top_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.14 130.075 6.28 130.56 ;
    END
  END chany_top_out[22]
  PIN chany_top_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.18 130.075 40.32 130.56 ;
    END
  END chany_top_out[23]
  PIN chany_top_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.22 130.075 28.36 130.56 ;
    END
  END chany_top_out[24]
  PIN chany_top_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.94 130.075 43.08 130.56 ;
    END
  END chany_top_out[25]
  PIN chany_top_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 130.075 41.24 130.56 ;
    END
  END chany_top_out[26]
  PIN chany_top_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.86 130.075 21 130.56 ;
    END
  END chany_top_out[27]
  PIN chany_top_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.94 130.075 20.08 130.56 ;
    END
  END chany_top_out[28]
  PIN chany_top_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.02 130.075 42.16 130.56 ;
    END
  END chany_top_out[29]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 61.64 103.96 61.78 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 20.16 103.96 20.3 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 27.98 103.96 28.12 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 64.36 103.96 64.5 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 25.35 103.96 25.65 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 30.7 103.96 30.84 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 66.15 103.96 66.45 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 13.79 103.96 14.09 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 22.63 103.96 22.93 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 58.92 103.96 59.06 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 56.2 103.96 56.34 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 18.12 103.96 18.26 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 60.96 103.96 61.1 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 12.43 103.96 12.73 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 31.38 103.96 31.52 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 55.52 103.96 55.66 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 11.07 103.96 11.37 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 22.88 103.96 23.02 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 63.43 103.96 63.73 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 11.66 103.96 11.8 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 17.44 103.96 17.58 ;
    END
  END chanx_right_out[20]
  PIN chanx_right_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 67.08 103.96 67.22 ;
    END
  END chanx_right_out[21]
  PIN chanx_right_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 20.84 103.96 20.98 ;
    END
  END chanx_right_out[22]
  PIN chanx_right_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 25.26 103.96 25.4 ;
    END
  END chanx_right_out[23]
  PIN chanx_right_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 88.84 103.96 88.98 ;
    END
  END chanx_right_out[24]
  PIN chanx_right_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 12.34 103.96 12.48 ;
    END
  END chanx_right_out[25]
  PIN chanx_right_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 28.66 103.96 28.8 ;
    END
  END chanx_right_out[26]
  PIN chanx_right_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 53.48 103.96 53.62 ;
    END
  END chanx_right_out[27]
  PIN chanx_right_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 25.94 103.96 26.08 ;
    END
  END chanx_right_out[28]
  PIN chanx_right_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 23.56 103.96 23.7 ;
    END
  END chanx_right_out[29]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.66 0 11.8 0.485 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 0 64.24 0.485 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.86 0 44 0.485 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.68 0 5.82 0.485 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.38 0 26.52 0.485 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.18 0 40.32 0.485 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.74 0 10.88 0.485 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.42 0 14.56 0.485 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.46 0 25.6 0.485 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 0 62.4 0.485 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.94 0 43.08 0.485 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 0 41.24 0.485 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.3 0 27.44 0.485 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.34 0 15.48 0.485 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.62 0 69.76 0.485 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.54 0 24.68 0.485 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.76 0 4.9 0.485 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.26 0 16.4 0.485 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.58 0 12.72 0.485 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.62 0 23.76 0.485 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.18 0 17.32 0.485 ;
    END
  END chany_bottom_out[20]
  PIN chany_bottom_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.7 0 22.84 0.485 ;
    END
  END chany_bottom_out[21]
  PIN chany_bottom_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.7 0 45.84 0.485 ;
    END
  END chany_bottom_out[22]
  PIN chany_bottom_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.1 0 18.24 0.485 ;
    END
  END chany_bottom_out[23]
  PIN chany_bottom_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 0 38.48 0.485 ;
    END
  END chany_bottom_out[24]
  PIN chany_bottom_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.78 0 21.92 0.485 ;
    END
  END chany_bottom_out[25]
  PIN chany_bottom_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.18 0 63.32 0.485 ;
    END
  END chany_bottom_out[26]
  PIN chany_bottom_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.02 0 19.16 0.485 ;
    END
  END chany_bottom_out[27]
  PIN chany_bottom_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.86 0 21 0.485 ;
    END
  END chany_bottom_out[28]
  PIN chany_bottom_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.94 0 20.08 0.485 ;
    END
  END chany_bottom_out[29]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.5 0 13.64 0.485 ;
    END
  END ccff_tail[0]
  PIN pReset_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 80.34 103.96 80.48 ;
    END
  END pReset_E_in
  PIN pReset_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.02 0 42.16 0.485 ;
    END
  END pReset_S_out
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 103.365 115.02 103.96 115.16 ;
    END
  END prog_clk_0_E_in
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 22.88 3.2 26.08 ;
        RECT 100.76 22.88 103.96 26.08 ;
        RECT 0 63.68 3.2 66.88 ;
        RECT 100.76 63.68 103.96 66.88 ;
        RECT 0 104.48 3.2 107.68 ;
        RECT 100.76 104.48 103.96 107.68 ;
      LAYER met4 ;
        RECT 14.42 0 15.02 0.6 ;
        RECT 43.86 0 44.46 0.6 ;
        RECT 89.86 5.44 90.46 6.04 ;
        RECT 89.86 124.52 90.46 125.12 ;
        RECT 14.42 129.96 15.02 130.56 ;
        RECT 43.86 129.96 44.46 130.56 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 73.12 2.48 73.6 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 103.48 7.92 103.96 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 103.48 13.36 103.96 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 103.48 18.8 103.96 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 103.48 24.24 103.96 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 103.48 29.68 103.96 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 103.48 35.12 103.96 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 103.48 40.56 103.96 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 103.48 46 103.96 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 103.48 51.44 103.96 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 103.48 56.88 103.96 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 103.48 62.32 103.96 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 103.48 67.76 103.96 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 103.48 73.2 103.96 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 103.48 78.64 103.96 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 103.48 84.08 103.96 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 103.48 89.52 103.96 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 103.48 94.96 103.96 95.44 ;
        RECT 0 100.4 0.48 100.88 ;
        RECT 103.48 100.4 103.96 100.88 ;
        RECT 0 105.84 0.48 106.32 ;
        RECT 103.48 105.84 103.96 106.32 ;
        RECT 0 111.28 0.48 111.76 ;
        RECT 103.48 111.28 103.96 111.76 ;
        RECT 0 116.72 0.48 117.2 ;
        RECT 103.48 116.72 103.96 117.2 ;
        RECT 0 122.16 0.48 122.64 ;
        RECT 103.48 122.16 103.96 122.64 ;
        RECT 0 127.6 0.48 128.08 ;
        RECT 73.12 127.6 73.6 128.08 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 43.28 3.2 46.48 ;
        RECT 100.76 43.28 103.96 46.48 ;
        RECT 0 84.08 3.2 87.28 ;
        RECT 100.76 84.08 103.96 87.28 ;
      LAYER met4 ;
        RECT 29.14 0 29.74 0.6 ;
        RECT 58.58 0 59.18 0.6 ;
        RECT 29.14 129.96 29.74 130.56 ;
        RECT 58.58 129.96 59.18 130.56 ;
      LAYER met1 ;
        RECT 0 -0.24 0.48 0.24 ;
        RECT 73.12 -0.24 73.6 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 103.48 5.2 103.96 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 103.48 10.64 103.96 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 103.48 16.08 103.96 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 103.48 21.52 103.96 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 103.48 26.96 103.96 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 103.48 32.4 103.96 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 103.48 37.84 103.96 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 103.48 43.28 103.96 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 103.48 48.72 103.96 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 103.48 54.16 103.96 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 103.48 59.6 103.96 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 103.48 65.04 103.96 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 103.48 70.48 103.96 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 103.48 75.92 103.96 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 103.48 81.36 103.96 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 103.48 86.8 103.96 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 103.48 92.24 103.96 92.72 ;
        RECT 0 97.68 0.48 98.16 ;
        RECT 103.48 97.68 103.96 98.16 ;
        RECT 0 103.12 0.48 103.6 ;
        RECT 103.48 103.12 103.96 103.6 ;
        RECT 0 108.56 0.48 109.04 ;
        RECT 103.48 108.56 103.96 109.04 ;
        RECT 0 114 0.48 114.48 ;
        RECT 103.48 114 103.96 114.48 ;
        RECT 0 119.44 0.48 119.92 ;
        RECT 103.48 119.44 103.96 119.92 ;
        RECT 0 124.88 0.48 125.36 ;
        RECT 103.48 124.88 103.96 125.36 ;
        RECT 0 130.32 0.48 130.8 ;
        RECT 73.12 130.32 73.6 130.8 ;
    END
  END VSS
  OBS
    LAYER met1 ;
      POLYGON 72.84 130.8 72.84 130.32 59.04 130.32 59.04 130.31 58.72 130.31 58.72 130.32 29.6 130.32 29.6 130.31 29.28 130.31 29.28 130.32 0.76 130.32 0.76 130.8 ;
      RECT 53.96 124.88 103.2 125.36 ;
      POLYGON 103.435 26.76 103.435 26.36 103.295 26.36 103.295 26.62 97.22 26.62 97.22 26.76 ;
      RECT 53.96 5.2 103.2 5.68 ;
      POLYGON 59.04 0.25 59.04 0.24 72.84 0.24 72.84 -0.24 0.76 -0.24 0.76 0.24 29.28 0.24 29.28 0.25 29.6 0.25 29.6 0.24 58.72 0.24 58.72 0.25 ;
      POLYGON 72.84 130.28 72.84 130.04 73.32 130.04 73.32 128.36 72.84 128.36 72.84 127.32 73.32 127.32 73.32 124.84 103.2 124.84 103.2 124.6 103.68 124.6 103.68 122.92 103.2 122.92 103.2 121.88 103.68 121.88 103.68 120.2 103.2 120.2 103.2 119.16 103.68 119.16 103.68 117.48 103.2 117.48 103.2 116.44 103.68 116.44 103.68 115.44 103.085 115.44 103.085 114.74 103.2 114.74 103.2 113.72 103.68 113.72 103.68 112.04 103.2 112.04 103.2 111 103.68 111 103.68 109.32 103.2 109.32 103.2 108.28 103.68 108.28 103.68 106.6 103.2 106.6 103.2 105.56 103.68 105.56 103.68 103.88 103.2 103.88 103.2 102.84 103.68 102.84 103.68 101.16 103.2 101.16 103.2 100.12 103.68 100.12 103.68 98.44 103.2 98.44 103.2 97.4 103.68 97.4 103.68 95.72 103.2 95.72 103.2 94.68 103.68 94.68 103.68 93 103.2 93 103.2 91.96 103.68 91.96 103.68 90.28 103.2 90.28 103.2 89.26 103.085 89.26 103.085 88.56 103.68 88.56 103.68 87.56 103.2 87.56 103.2 86.52 103.68 86.52 103.68 84.84 103.2 84.84 103.2 83.8 103.68 83.8 103.68 82.12 103.2 82.12 103.2 81.08 103.68 81.08 103.68 80.76 103.085 80.76 103.085 80.06 103.68 80.06 103.68 79.4 103.2 79.4 103.2 78.36 103.68 78.36 103.68 76.68 103.2 76.68 103.2 75.64 103.68 75.64 103.68 73.96 103.2 73.96 103.2 72.92 103.68 72.92 103.68 71.24 103.2 71.24 103.2 70.2 103.68 70.2 103.68 68.52 103.2 68.52 103.2 67.5 103.085 67.5 103.085 66.12 103.68 66.12 103.68 65.8 103.2 65.8 103.2 64.78 103.085 64.78 103.085 63.4 103.68 63.4 103.68 63.08 103.2 63.08 103.2 62.06 103.085 62.06 103.085 60.68 103.68 60.68 103.68 60.36 103.2 60.36 103.2 59.34 103.085 59.34 103.085 57.96 103.68 57.96 103.68 57.64 103.2 57.64 103.2 56.62 103.085 56.62 103.085 55.24 103.68 55.24 103.68 54.92 103.2 54.92 103.2 53.9 103.085 53.9 103.085 53.2 103.68 53.2 103.68 52.88 103.085 52.88 103.085 52.18 103.2 52.18 103.2 51.16 103.68 51.16 103.68 50.84 103.085 50.84 103.085 49.46 103.2 49.46 103.2 48.44 103.68 48.44 103.68 48.12 103.085 48.12 103.085 46.74 103.2 46.74 103.2 45.74 103.085 45.74 103.085 44.36 103.68 44.36 103.68 44.04 103.2 44.04 103.2 43.02 103.085 43.02 103.085 41.64 103.68 41.64 103.68 41.32 103.2 41.32 103.2 40.3 103.085 40.3 103.085 38.92 103.68 38.92 103.68 38.6 103.2 38.6 103.2 37.58 103.085 37.58 103.085 36.2 103.68 36.2 103.68 35.88 103.2 35.88 103.2 34.84 103.68 34.84 103.68 34.52 103.085 34.52 103.085 33.14 103.2 33.14 103.2 32.12 103.68 32.12 103.68 31.8 103.085 31.8 103.085 30.42 103.2 30.42 103.2 29.4 103.68 29.4 103.68 29.08 103.085 29.08 103.085 27.7 103.2 27.7 103.2 26.68 103.68 26.68 103.68 26.36 103.085 26.36 103.085 24.98 103.2 24.98 103.2 23.98 103.085 23.98 103.085 22.6 103.68 22.6 103.68 22.28 103.2 22.28 103.2 21.26 103.085 21.26 103.085 19.88 103.68 19.88 103.68 19.56 103.2 19.56 103.2 18.54 103.085 18.54 103.085 17.16 103.68 17.16 103.68 16.84 103.2 16.84 103.2 15.82 103.085 15.82 103.085 14.44 103.68 14.44 103.68 14.12 103.2 14.12 103.2 13.08 103.68 13.08 103.68 12.76 103.085 12.76 103.085 11.38 103.2 11.38 103.2 10.36 103.68 10.36 103.68 8.68 103.2 8.68 103.2 7.64 103.68 7.64 103.68 5.96 103.2 5.96 103.2 5.72 73.32 5.72 73.32 3.24 72.84 3.24 72.84 2.2 73.32 2.2 73.32 0.52 72.84 0.52 72.84 0.28 0.76 0.28 0.76 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.08 0.875 64.08 0.875 64.78 0.76 64.78 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 0.76 97.4 0.76 98.44 0.28 98.44 0.28 100.12 0.76 100.12 0.76 101.16 0.28 101.16 0.28 102.84 0.76 102.84 0.76 103.88 0.28 103.88 0.28 105.56 0.76 105.56 0.76 106.6 0.28 106.6 0.28 108.28 0.76 108.28 0.76 109.32 0.28 109.32 0.28 111 0.76 111 0.76 112.04 0.28 112.04 0.28 113.72 0.76 113.72 0.76 114.76 0.28 114.76 0.28 116.44 0.76 116.44 0.76 117.48 0.28 117.48 0.28 119.16 0.76 119.16 0.76 120.2 0.28 120.2 0.28 121.88 0.76 121.88 0.76 122.92 0.28 122.92 0.28 124.6 0.76 124.6 0.76 125.64 0.28 125.64 0.28 127.32 0.76 127.32 0.76 128.36 0.28 128.36 0.28 130.04 0.76 130.04 0.76 130.28 ;
    LAYER met4 ;
      POLYGON 20.85 130.37 20.85 96.24 20.55 96.24 20.55 130.07 20.33 130.07 20.33 130.37 ;
      POLYGON 86.17 16.98 86.17 5.945 86.185 5.945 86.185 5.615 85.855 5.615 85.855 5.945 85.87 5.945 85.87 16.98 ;
      POLYGON 73.2 130.16 73.2 124.72 89.46 124.72 89.46 124.12 90.86 124.12 90.86 124.72 103.56 124.72 103.56 5.84 90.86 5.84 90.86 6.44 89.46 6.44 89.46 5.84 73.2 5.84 73.2 0.4 59.58 0.4 59.58 1 58.18 1 58.18 0.4 44.86 0.4 44.86 1 43.46 1 43.46 0.4 30.14 0.4 30.14 1 28.74 1 28.74 0.4 15.42 0.4 15.42 1 14.02 1 14.02 0.4 0.4 0.4 0.4 130.16 14.02 130.16 14.02 129.56 15.42 129.56 15.42 130.16 19.23 130.16 19.23 129.36 20.33 129.36 20.33 130.16 28.74 130.16 28.74 129.56 30.14 129.56 30.14 130.16 43.46 130.16 43.46 129.56 44.86 129.56 44.86 130.16 58.18 130.16 58.18 129.56 59.58 129.56 59.58 130.16 ;
    LAYER met2 ;
      RECT 58.74 130.255 59.02 130.625 ;
      RECT 29.3 130.255 29.58 130.625 ;
      POLYGON 39.86 130.46 39.86 104.48 39.72 104.48 39.72 130.32 39.68 130.32 39.68 130.46 ;
      POLYGON 73.51 124.965 73.51 124.595 73.44 124.595 73.44 114.51 73.3 114.51 73.3 124.595 73.23 124.595 73.23 124.965 ;
      POLYGON 22.38 27.1 22.38 0.24 22.42 0.24 22.42 0.1 22.24 0.1 22.24 27.1 ;
      POLYGON 86.32 12.82 86.32 5.85 88.94 5.85 88.94 6.13 88.88 6.13 88.88 6.45 89.14 6.45 89.14 6.13 89.08 6.13 89.08 5.71 86.18 5.71 86.18 12.82 ;
      RECT 58.74 -0.065 59.02 0.305 ;
      RECT 29.3 -0.065 29.58 0.305 ;
      POLYGON 73.32 130.28 73.32 124.84 103.68 124.84 103.68 5.72 97.18 5.72 97.18 6.205 96.48 6.205 96.48 5.72 96.26 5.72 96.26 6.205 95.56 6.205 95.56 5.72 95.34 5.72 95.34 6.205 94.64 6.205 94.64 5.72 94.42 5.72 94.42 6.205 93.72 6.205 93.72 5.72 93.5 5.72 93.5 6.205 92.8 6.205 92.8 5.72 91.66 5.72 91.66 6.205 90.96 6.205 90.96 5.72 90.74 5.72 90.74 6.205 90.04 6.205 90.04 5.72 89.82 5.72 89.82 6.205 89.12 6.205 89.12 5.72 73.32 5.72 73.32 0.28 71.42 0.28 71.42 0.765 70.72 0.765 70.72 0.28 70.04 0.28 70.04 0.765 69.34 0.765 69.34 0.28 69.12 0.28 69.12 0.765 68.42 0.765 68.42 0.28 68.2 0.28 68.2 0.765 67.5 0.765 67.5 0.28 67.28 0.28 67.28 0.765 66.58 0.765 66.58 0.28 66.36 0.28 66.36 0.765 65.66 0.765 65.66 0.28 65.44 0.28 65.44 0.765 64.74 0.765 64.74 0.28 64.52 0.28 64.52 0.765 63.82 0.765 63.82 0.28 63.6 0.28 63.6 0.765 62.9 0.765 62.9 0.28 62.68 0.28 62.68 0.765 61.98 0.765 61.98 0.28 61.76 0.28 61.76 0.765 61.06 0.765 61.06 0.28 60.84 0.28 60.84 0.765 60.14 0.765 60.14 0.28 59.92 0.28 59.92 0.765 59.22 0.765 59.22 0.28 58.54 0.28 58.54 0.765 57.84 0.765 57.84 0.28 57.62 0.28 57.62 0.765 56.92 0.765 56.92 0.28 56.7 0.28 56.7 0.765 56 0.765 56 0.28 55.78 0.28 55.78 0.765 55.08 0.765 55.08 0.28 54.86 0.28 54.86 0.765 54.16 0.765 54.16 0.28 53.94 0.28 53.94 0.765 53.24 0.765 53.24 0.28 48.88 0.28 48.88 0.765 48.18 0.765 48.18 0.28 47.96 0.28 47.96 0.765 47.26 0.765 47.26 0.28 47.04 0.28 47.04 0.765 46.34 0.765 46.34 0.28 46.12 0.28 46.12 0.765 45.42 0.765 45.42 0.28 45.2 0.28 45.2 0.765 44.5 0.765 44.5 0.28 44.28 0.28 44.28 0.765 43.58 0.765 43.58 0.28 43.36 0.28 43.36 0.765 42.66 0.765 42.66 0.28 42.44 0.28 42.44 0.765 41.74 0.765 41.74 0.28 41.52 0.28 41.52 0.765 40.82 0.765 40.82 0.28 40.6 0.28 40.6 0.765 39.9 0.765 39.9 0.28 39.68 0.28 39.68 0.765 38.98 0.765 38.98 0.28 38.76 0.28 38.76 0.765 38.06 0.765 38.06 0.28 37.84 0.28 37.84 0.765 37.14 0.765 37.14 0.28 36.92 0.28 36.92 0.765 36.22 0.765 36.22 0.28 36 0.28 36 0.765 35.3 0.765 35.3 0.28 35.08 0.28 35.08 0.765 34.38 0.765 34.38 0.28 34.16 0.28 34.16 0.765 33.46 0.765 33.46 0.28 33.24 0.28 33.24 0.765 32.54 0.765 32.54 0.28 27.72 0.28 27.72 0.765 27.02 0.765 27.02 0.28 26.8 0.28 26.8 0.765 26.1 0.765 26.1 0.28 25.88 0.28 25.88 0.765 25.18 0.765 25.18 0.28 24.96 0.28 24.96 0.765 24.26 0.765 24.26 0.28 24.04 0.28 24.04 0.765 23.34 0.765 23.34 0.28 23.12 0.28 23.12 0.765 22.42 0.765 22.42 0.28 22.2 0.28 22.2 0.765 21.5 0.765 21.5 0.28 21.28 0.28 21.28 0.765 20.58 0.765 20.58 0.28 20.36 0.28 20.36 0.765 19.66 0.765 19.66 0.28 19.44 0.28 19.44 0.765 18.74 0.765 18.74 0.28 18.52 0.28 18.52 0.765 17.82 0.765 17.82 0.28 17.6 0.28 17.6 0.765 16.9 0.765 16.9 0.28 16.68 0.28 16.68 0.765 15.98 0.765 15.98 0.28 15.76 0.28 15.76 0.765 15.06 0.765 15.06 0.28 14.84 0.28 14.84 0.765 14.14 0.765 14.14 0.28 13.92 0.28 13.92 0.765 13.22 0.765 13.22 0.28 13 0.28 13 0.765 12.3 0.765 12.3 0.28 12.08 0.28 12.08 0.765 11.38 0.765 11.38 0.28 11.16 0.28 11.16 0.765 10.46 0.765 10.46 0.28 10.24 0.28 10.24 0.765 9.54 0.765 9.54 0.28 9.32 0.28 9.32 0.765 8.62 0.765 8.62 0.28 8.4 0.28 8.4 0.765 7.7 0.765 7.7 0.28 7.48 0.28 7.48 0.765 6.78 0.765 6.78 0.28 6.1 0.28 6.1 0.765 5.4 0.765 5.4 0.28 5.18 0.28 5.18 0.765 4.48 0.765 4.48 0.28 4.26 0.28 4.26 0.765 3.56 0.765 3.56 0.28 0.28 0.28 0.28 130.28 3.56 130.28 3.56 129.795 4.26 129.795 4.26 130.28 4.48 130.28 4.48 129.795 5.18 129.795 5.18 130.28 5.86 130.28 5.86 129.795 6.56 129.795 6.56 130.28 6.78 130.28 6.78 129.795 7.48 129.795 7.48 130.28 7.7 130.28 7.7 129.795 8.4 129.795 8.4 130.28 8.62 130.28 8.62 129.795 9.32 129.795 9.32 130.28 9.54 130.28 9.54 129.795 10.24 129.795 10.24 130.28 10.46 130.28 10.46 129.795 11.16 129.795 11.16 130.28 11.38 130.28 11.38 129.795 12.08 129.795 12.08 130.28 12.3 130.28 12.3 129.795 13 129.795 13 130.28 13.22 130.28 13.22 129.795 13.92 129.795 13.92 130.28 14.14 130.28 14.14 129.795 14.84 129.795 14.84 130.28 15.06 130.28 15.06 129.795 15.76 129.795 15.76 130.28 15.98 130.28 15.98 129.795 16.68 129.795 16.68 130.28 16.9 130.28 16.9 129.795 17.6 129.795 17.6 130.28 17.82 130.28 17.82 129.795 18.52 129.795 18.52 130.28 18.74 130.28 18.74 129.795 19.44 129.795 19.44 130.28 19.66 130.28 19.66 129.795 20.36 129.795 20.36 130.28 20.58 130.28 20.58 129.795 21.28 129.795 21.28 130.28 21.5 130.28 21.5 129.795 22.2 129.795 22.2 130.28 22.42 130.28 22.42 129.795 23.12 129.795 23.12 130.28 23.34 130.28 23.34 129.795 24.04 129.795 24.04 130.28 24.26 130.28 24.26 129.795 24.96 129.795 24.96 130.28 25.18 130.28 25.18 129.795 25.88 129.795 25.88 130.28 26.1 130.28 26.1 129.795 26.8 129.795 26.8 130.28 27.02 130.28 27.02 129.795 27.72 129.795 27.72 130.28 27.94 130.28 27.94 129.795 28.64 129.795 28.64 130.28 29.78 130.28 29.78 129.795 30.48 129.795 30.48 130.28 35.3 130.28 35.3 129.795 36 129.795 36 130.28 36.22 130.28 36.22 129.795 36.92 129.795 36.92 130.28 37.14 130.28 37.14 129.795 37.84 129.795 37.84 130.28 38.06 130.28 38.06 129.795 38.76 129.795 38.76 130.28 38.98 130.28 38.98 129.795 39.68 129.795 39.68 130.28 39.9 130.28 39.9 129.795 40.6 129.795 40.6 130.28 40.82 130.28 40.82 129.795 41.52 129.795 41.52 130.28 41.74 130.28 41.74 129.795 42.44 129.795 42.44 130.28 42.66 130.28 42.66 129.795 43.36 129.795 43.36 130.28 43.58 130.28 43.58 129.795 44.28 129.795 44.28 130.28 44.5 130.28 44.5 129.795 45.2 129.795 45.2 130.28 45.42 130.28 45.42 129.795 46.12 129.795 46.12 130.28 46.34 130.28 46.34 129.795 47.04 129.795 47.04 130.28 47.26 130.28 47.26 129.795 47.96 129.795 47.96 130.28 52.78 130.28 52.78 129.795 53.48 129.795 53.48 130.28 55.08 130.28 55.08 129.795 55.78 129.795 55.78 130.28 56 130.28 56 129.795 56.7 129.795 56.7 130.28 56.92 130.28 56.92 129.795 57.62 129.795 57.62 130.28 57.84 130.28 57.84 129.795 58.54 129.795 58.54 130.28 59.22 130.28 59.22 129.795 59.92 129.795 59.92 130.28 60.14 130.28 60.14 129.795 60.84 129.795 60.84 130.28 61.06 130.28 61.06 129.795 61.76 129.795 61.76 130.28 61.98 130.28 61.98 129.795 62.68 129.795 62.68 130.28 62.9 130.28 62.9 129.795 63.6 129.795 63.6 130.28 63.82 130.28 63.82 129.795 64.52 129.795 64.52 130.28 64.74 130.28 64.74 129.795 65.44 129.795 65.44 130.28 65.66 130.28 65.66 129.795 66.36 129.795 66.36 130.28 66.58 130.28 66.58 129.795 67.28 129.795 67.28 130.28 67.5 130.28 67.5 129.795 68.2 129.795 68.2 130.28 68.42 130.28 68.42 129.795 69.12 129.795 69.12 130.28 69.8 130.28 69.8 129.795 70.5 129.795 70.5 130.28 70.72 130.28 70.72 129.795 71.42 129.795 71.42 130.28 ;
    LAYER met3 ;
      POLYGON 59.045 130.605 59.045 130.6 59.26 130.6 59.26 130.28 59.045 130.28 59.045 130.275 58.715 130.275 58.715 130.28 58.5 130.28 58.5 130.6 58.715 130.6 58.715 130.605 ;
      POLYGON 29.605 130.605 29.605 130.6 29.82 130.6 29.82 130.28 29.605 130.28 29.605 130.275 29.275 130.275 29.275 130.28 29.06 130.28 29.06 130.6 29.275 130.6 29.275 130.605 ;
      POLYGON 73.535 124.945 73.535 124.615 73.205 124.615 73.205 124.63 68.39 124.63 68.39 124.93 73.205 124.93 73.205 124.945 ;
      POLYGON 95.155 5.945 95.155 5.615 94.825 5.615 94.825 5.63 86.21 5.63 86.21 5.62 85.83 5.62 85.83 5.94 86.21 5.94 86.21 5.93 94.825 5.93 94.825 5.945 ;
      POLYGON 59.045 0.285 59.045 0.28 59.26 0.28 59.26 -0.04 59.045 -0.04 59.045 -0.045 58.715 -0.045 58.715 -0.04 58.5 -0.04 58.5 0.28 58.715 0.28 58.715 0.285 ;
      POLYGON 29.605 0.285 29.605 0.28 29.82 0.28 29.82 -0.04 29.605 -0.04 29.605 -0.045 29.275 -0.045 29.275 -0.04 29.06 -0.04 29.06 0.28 29.275 0.28 29.275 0.285 ;
      POLYGON 73.2 130.16 73.2 124.72 103.56 124.72 103.56 68.21 102.76 68.21 102.76 67.11 103.56 67.11 103.56 66.85 102.76 66.85 102.76 65.75 103.56 65.75 103.56 65.49 102.76 65.49 102.76 64.39 103.56 64.39 103.56 64.13 102.76 64.13 102.76 63.03 103.56 63.03 103.56 62.77 102.76 62.77 102.76 61.67 103.56 61.67 103.56 61.41 102.76 61.41 102.76 60.31 103.56 60.31 103.56 60.05 102.76 60.05 102.76 58.95 103.56 58.95 103.56 47.81 102.76 47.81 102.76 46.71 103.56 46.71 103.56 46.45 102.76 46.45 102.76 45.35 103.56 45.35 103.56 45.09 102.76 45.09 102.76 43.99 103.56 43.99 103.56 27.41 102.76 27.41 102.76 26.31 103.56 26.31 103.56 26.05 102.76 26.05 102.76 24.95 103.56 24.95 103.56 24.69 102.76 24.69 102.76 23.59 103.56 23.59 103.56 23.33 102.76 23.33 102.76 22.23 103.56 22.23 103.56 21.97 102.76 21.97 102.76 20.87 103.56 20.87 103.56 14.49 102.76 14.49 102.76 13.39 103.56 13.39 103.56 13.13 102.76 13.13 102.76 12.03 103.56 12.03 103.56 11.77 102.76 11.77 102.76 10.67 103.56 10.67 103.56 5.84 73.2 5.84 73.2 0.4 0.4 0.4 0.4 130.16 ;
    LAYER met5 ;
      POLYGON 72 128.96 72 123.52 102.36 123.52 102.36 109.28 99.16 109.28 99.16 102.88 102.36 102.88 102.36 88.88 99.16 88.88 99.16 82.48 102.36 82.48 102.36 68.48 99.16 68.48 99.16 62.08 102.36 62.08 102.36 48.08 99.16 48.08 99.16 41.68 102.36 41.68 102.36 27.68 99.16 27.68 99.16 21.28 102.36 21.28 102.36 7.04 72 7.04 72 1.6 1.6 1.6 1.6 21.28 4.8 21.28 4.8 27.68 1.6 27.68 1.6 41.68 4.8 41.68 4.8 48.08 1.6 48.08 1.6 62.08 4.8 62.08 4.8 68.48 1.6 68.48 1.6 82.48 4.8 82.48 4.8 88.88 1.6 88.88 1.6 102.88 4.8 102.88 4.8 109.28 1.6 109.28 1.6 128.96 ;
    LAYER li1 ;
      POLYGON 73.6 130.645 73.6 130.475 70.125 130.475 70.125 130.015 69.87 130.015 69.87 130.475 69.2 130.475 69.2 130.015 69.03 130.015 69.03 130.475 68.36 130.475 68.36 130.015 68.19 130.015 68.19 130.475 67.52 130.475 67.52 130.015 67.35 130.015 67.35 130.475 66.68 130.475 66.68 130.015 66.375 130.015 66.375 130.475 65.805 130.475 65.805 129.995 65.635 129.995 65.635 130.475 64.965 130.475 64.965 129.995 64.795 129.995 64.795 130.475 64.205 130.475 64.205 129.995 63.875 129.995 63.875 130.475 63.365 130.475 63.365 129.995 63.035 129.995 63.035 130.475 62.525 130.475 62.525 129.675 62.195 129.675 62.195 130.475 56.525 130.475 56.525 129.995 56.195 129.995 56.195 130.475 55.685 130.475 55.685 129.995 55.355 129.995 55.355 130.475 54.845 130.475 54.845 129.995 54.515 129.995 54.515 130.475 54.005 130.475 54.005 129.995 53.675 129.995 53.675 130.475 53.165 130.475 53.165 129.995 52.835 129.995 52.835 130.475 52.325 130.475 52.325 129.675 51.995 129.675 51.995 130.475 50.085 130.475 50.085 129.995 49.755 129.995 49.755 130.475 49.245 130.475 49.245 129.995 48.915 129.995 48.915 130.475 48.405 130.475 48.405 129.995 48.075 129.995 48.075 130.475 47.565 130.475 47.565 129.995 47.235 129.995 47.235 130.475 46.725 130.475 46.725 129.995 46.395 129.995 46.395 130.475 45.885 130.475 45.885 129.675 45.555 129.675 45.555 130.475 44.025 130.475 44.025 130.015 43.72 130.015 43.72 130.475 43.05 130.475 43.05 130.015 42.88 130.015 42.88 130.475 42.21 130.475 42.21 130.015 42.04 130.015 42.04 130.475 41.37 130.475 41.37 130.015 41.2 130.015 41.2 130.475 40.53 130.475 40.53 130.015 40.275 130.015 40.275 130.475 37.665 130.475 37.665 129.995 37.335 129.995 37.335 130.475 36.825 130.475 36.825 129.995 36.495 129.995 36.495 130.475 35.985 130.475 35.985 129.995 35.655 129.995 35.655 130.475 35.145 130.475 35.145 129.995 34.815 129.995 34.815 130.475 34.305 130.475 34.305 129.995 33.975 129.995 33.975 130.475 33.465 130.475 33.465 129.675 33.135 129.675 33.135 130.475 31.265 130.475 31.265 129.675 30.935 129.675 30.935 130.475 30.425 130.475 30.425 129.995 30.095 129.995 30.095 130.475 29.585 130.475 29.585 129.995 29.255 129.995 29.255 130.475 28.745 130.475 28.745 129.995 28.415 129.995 28.415 130.475 27.905 130.475 27.905 129.995 27.575 129.995 27.575 130.475 27.065 130.475 27.065 129.995 26.735 129.995 26.735 130.475 25.285 130.475 25.285 129.675 24.955 129.675 24.955 130.475 24.445 130.475 24.445 129.995 24.115 129.995 24.115 130.475 23.605 130.475 23.605 129.995 23.275 129.995 23.275 130.475 22.765 130.475 22.765 129.995 22.435 129.995 22.435 130.475 21.925 130.475 21.925 129.995 21.595 129.995 21.595 130.475 21.085 130.475 21.085 129.995 20.755 129.995 20.755 130.475 18.845 130.475 18.845 129.675 18.515 129.675 18.515 130.475 18.005 130.475 18.005 129.995 17.675 129.995 17.675 130.475 17.165 130.475 17.165 129.995 16.835 129.995 16.835 130.475 16.325 130.475 16.325 129.995 15.995 129.995 15.995 130.475 15.485 130.475 15.485 129.995 15.155 129.995 15.155 130.475 14.645 130.475 14.645 129.995 14.315 129.995 14.315 130.475 11.985 130.475 11.985 129.995 11.815 129.995 11.815 130.475 11.145 130.475 11.145 129.995 10.975 129.995 10.975 130.475 10.385 130.475 10.385 129.995 10.055 129.995 10.055 130.475 9.545 130.475 9.545 129.995 9.215 129.995 9.215 130.475 8.705 130.475 8.705 129.675 8.375 129.675 8.375 130.475 0 130.475 0 130.645 ;
      RECT 72.68 127.755 73.6 127.925 ;
      RECT 0 127.755 3.68 127.925 ;
      POLYGON 103.96 125.205 103.96 125.035 97.435 125.035 97.435 124.235 97.125 124.235 97.125 125.035 95.135 125.035 95.135 124.53 94.85 124.53 94.85 125.035 92.825 125.035 92.825 124.225 92.555 124.225 92.555 125.035 91.885 125.035 91.885 124.225 91.645 124.225 91.645 125.035 90.25 125.035 90.25 124.215 90.02 124.215 90.02 125.035 87.77 125.035 87.77 124.53 87.485 124.53 87.485 125.035 86.855 125.035 86.855 124.53 86.57 124.53 86.57 125.035 84.14 125.035 84.14 124.3 83.8 124.3 83.8 125.035 83.045 125.035 83.045 124.3 82.705 124.3 82.705 125.035 74.605 125.035 74.605 124.3 74.275 124.3 74.275 125.035 72.68 125.035 72.68 125.205 ;
      RECT 0 125.035 3.68 125.205 ;
      RECT 103.04 122.315 103.96 122.485 ;
      RECT 0 122.315 1.84 122.485 ;
      RECT 103.5 119.595 103.96 119.765 ;
      RECT 0 119.595 1.84 119.765 ;
      RECT 103.5 116.875 103.96 117.045 ;
      RECT 0 116.875 3.68 117.045 ;
      RECT 103.5 114.155 103.96 114.325 ;
      RECT 0 114.155 3.68 114.325 ;
      RECT 103.5 111.435 103.96 111.605 ;
      RECT 0 111.435 1.84 111.605 ;
      RECT 103.5 108.715 103.96 108.885 ;
      RECT 0 108.715 3.68 108.885 ;
      RECT 100.28 105.995 103.96 106.165 ;
      RECT 0 105.995 3.68 106.165 ;
      RECT 100.28 103.275 103.96 103.445 ;
      RECT 0 103.275 3.68 103.445 ;
      RECT 100.28 100.555 103.96 100.725 ;
      RECT 0 100.555 1.84 100.725 ;
      RECT 100.28 97.835 103.96 98.005 ;
      RECT 0 97.835 1.84 98.005 ;
      RECT 100.28 95.115 103.96 95.285 ;
      RECT 0 95.115 1.84 95.285 ;
      RECT 103.04 92.395 103.96 92.565 ;
      RECT 0 92.395 1.84 92.565 ;
      RECT 103.04 89.675 103.96 89.845 ;
      RECT 0 89.675 1.84 89.845 ;
      RECT 103.04 86.955 103.96 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 103.04 84.235 103.96 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 103.04 81.515 103.96 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 103.04 78.795 103.96 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 103.04 76.075 103.96 76.245 ;
      RECT 0 76.075 1.84 76.245 ;
      RECT 103.04 73.355 103.96 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 103.04 70.635 103.96 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 103.04 67.915 103.96 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 103.04 65.195 103.96 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 103.04 62.475 103.96 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 103.04 59.755 103.96 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 103.04 57.035 103.96 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 103.04 54.315 103.96 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 103.04 51.595 103.96 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 100.28 48.875 103.96 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 100.28 46.155 103.96 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 100.28 43.435 103.96 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 103.04 40.715 103.96 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 103.04 37.995 103.96 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 103.04 35.275 103.96 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 103.04 32.555 103.96 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 103.04 29.835 103.96 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 103.04 27.115 103.96 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 103.04 24.395 103.96 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 103.04 21.675 103.96 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 103.04 18.955 103.96 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 103.04 16.235 103.96 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 103.04 13.515 103.96 13.685 ;
      RECT 0 13.515 1.84 13.685 ;
      RECT 103.04 10.795 103.96 10.965 ;
      RECT 0 10.795 1.84 10.965 ;
      RECT 103.5 8.075 103.96 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      POLYGON 100.645 6.325 100.645 5.525 103.96 5.525 103.96 5.355 73.14 5.355 73.14 5.525 73.655 5.525 73.655 6.005 73.985 6.005 73.985 5.525 74.495 5.525 74.495 6.005 74.825 6.005 74.825 5.525 75.335 5.525 75.335 6.005 75.665 6.005 75.665 5.525 76.175 5.525 76.175 6.005 76.505 6.005 76.505 5.525 77.015 5.525 77.015 6.005 77.345 6.005 77.345 5.525 77.855 5.525 77.855 6.325 78.185 6.325 78.185 5.525 79.945 5.525 79.945 6.06 80.455 6.06 80.455 5.525 82.415 5.525 82.415 5.925 82.745 5.925 82.745 5.525 87.305 5.525 87.305 6.06 87.815 6.06 87.815 5.525 89.775 5.525 89.775 5.925 90.105 5.925 90.105 5.525 91.975 5.525 91.975 6.005 92.145 6.005 92.145 5.525 92.815 5.525 92.815 6.005 92.985 6.005 92.985 5.525 93.575 5.525 93.575 6.005 93.905 6.005 93.905 5.525 94.415 5.525 94.415 6.005 94.745 6.005 94.745 5.525 95.255 5.525 95.255 6.325 95.585 6.325 95.585 5.525 97.035 5.525 97.035 6.005 97.205 6.005 97.205 5.525 97.875 5.525 97.875 6.005 98.045 6.005 98.045 5.525 98.635 5.525 98.635 6.005 98.965 6.005 98.965 5.525 99.475 5.525 99.475 6.005 99.805 6.005 99.805 5.525 100.315 5.525 100.315 6.325 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 73.14 2.635 73.6 2.805 ;
      RECT 0 2.635 1.84 2.805 ;
      POLYGON 65.665 0.885 65.665 0.085 66.175 0.085 66.175 0.565 66.505 0.565 66.505 0.085 67.015 0.085 67.015 0.565 67.345 0.565 67.345 0.085 67.855 0.085 67.855 0.565 68.185 0.565 68.185 0.085 68.695 0.085 68.695 0.565 69.025 0.565 69.025 0.085 69.535 0.085 69.535 0.565 69.865 0.565 69.865 0.085 73.6 0.085 73.6 -0.085 0 -0.085 0 0.085 2.855 0.085 2.855 0.885 3.185 0.885 3.185 0.085 3.695 0.085 3.695 0.565 4.025 0.565 4.025 0.085 4.535 0.085 4.535 0.565 4.865 0.565 4.865 0.085 5.455 0.085 5.455 0.565 5.625 0.565 5.625 0.085 6.295 0.085 6.295 0.565 6.465 0.565 6.465 0.085 7.875 0.085 7.875 0.565 8.205 0.565 8.205 0.085 8.715 0.085 8.715 0.565 9.045 0.565 9.045 0.085 9.555 0.085 9.555 0.565 9.885 0.565 9.885 0.085 10.395 0.085 10.395 0.565 10.725 0.565 10.725 0.085 11.235 0.085 11.235 0.565 11.565 0.565 11.565 0.085 12.075 0.085 12.075 0.885 12.405 0.885 12.405 0.085 13.435 0.085 13.435 0.885 13.765 0.885 13.765 0.085 14.275 0.085 14.275 0.565 14.605 0.565 14.605 0.085 15.115 0.085 15.115 0.565 15.445 0.565 15.445 0.085 16.035 0.085 16.035 0.565 16.205 0.565 16.205 0.085 16.875 0.085 16.875 0.565 17.045 0.565 17.045 0.085 17.575 0.085 17.575 0.885 17.905 0.885 17.905 0.085 18.415 0.085 18.415 0.565 18.745 0.565 18.745 0.085 19.255 0.085 19.255 0.565 19.585 0.565 19.585 0.085 20.175 0.085 20.175 0.565 20.345 0.565 20.345 0.085 21.015 0.085 21.015 0.565 21.185 0.565 21.185 0.085 24.055 0.085 24.055 0.545 24.36 0.545 24.36 0.085 25.03 0.085 25.03 0.545 25.2 0.545 25.2 0.085 25.87 0.085 25.87 0.545 26.04 0.545 26.04 0.085 26.71 0.085 26.71 0.545 26.88 0.545 26.88 0.085 27.55 0.085 27.55 0.545 27.805 0.545 27.805 0.085 29.455 0.085 29.455 0.885 29.785 0.885 29.785 0.085 30.295 0.085 30.295 0.565 30.625 0.565 30.625 0.085 31.135 0.085 31.135 0.565 31.465 0.565 31.465 0.085 31.975 0.085 31.975 0.565 32.305 0.565 32.305 0.085 32.815 0.085 32.815 0.565 33.145 0.565 33.145 0.085 33.655 0.085 33.655 0.565 33.985 0.565 33.985 0.085 35.895 0.085 35.895 0.885 36.225 0.885 36.225 0.085 36.735 0.085 36.735 0.565 37.065 0.565 37.065 0.085 37.575 0.085 37.575 0.565 37.905 0.565 37.905 0.085 38.415 0.085 38.415 0.565 38.745 0.565 38.745 0.085 39.255 0.085 39.255 0.565 39.585 0.565 39.585 0.085 40.095 0.085 40.095 0.565 40.425 0.565 40.425 0.085 41.875 0.085 41.875 0.885 42.205 0.885 42.205 0.085 42.715 0.085 42.715 0.565 43.045 0.565 43.045 0.085 43.555 0.085 43.555 0.565 43.885 0.565 43.885 0.085 44.395 0.085 44.395 0.565 44.725 0.565 44.725 0.085 45.235 0.085 45.235 0.565 45.565 0.565 45.565 0.085 46.075 0.085 46.075 0.565 46.405 0.565 46.405 0.085 47.635 0.085 47.635 0.545 47.89 0.545 47.89 0.085 48.56 0.085 48.56 0.545 48.73 0.545 48.73 0.085 49.4 0.085 49.4 0.545 49.57 0.545 49.57 0.085 50.24 0.085 50.24 0.545 50.41 0.545 50.41 0.085 51.08 0.085 51.08 0.545 51.385 0.545 51.385 0.085 53.415 0.085 53.415 0.565 53.745 0.565 53.745 0.085 54.255 0.085 54.255 0.565 54.585 0.565 54.585 0.085 55.095 0.085 55.095 0.565 55.425 0.565 55.425 0.085 55.935 0.085 55.935 0.565 56.265 0.565 56.265 0.085 56.775 0.085 56.775 0.565 57.105 0.565 57.105 0.085 57.615 0.085 57.615 0.885 57.945 0.885 57.945 0.085 59.595 0.085 59.595 0.545 59.85 0.545 59.85 0.085 60.52 0.085 60.52 0.545 60.69 0.545 60.69 0.085 61.36 0.085 61.36 0.545 61.53 0.545 61.53 0.085 62.2 0.085 62.2 0.545 62.37 0.545 62.37 0.085 63.04 0.085 63.04 0.545 63.345 0.545 63.345 0.085 65.335 0.085 65.335 0.885 ;
      POLYGON 73.43 130.39 73.43 124.95 103.79 124.95 103.79 5.61 73.43 5.61 73.43 0.17 0.17 0.17 0.17 130.39 ;
    LAYER mcon ;
      RECT 84.325 125.035 84.495 125.205 ;
      RECT 83.865 125.035 84.035 125.205 ;
      RECT 83.405 125.035 83.575 125.205 ;
      RECT 82.945 125.035 83.115 125.205 ;
      RECT 82.485 125.035 82.655 125.205 ;
      RECT 82.025 125.035 82.195 125.205 ;
      RECT 81.565 125.035 81.735 125.205 ;
      RECT 81.105 125.035 81.275 125.205 ;
      RECT 80.645 125.035 80.815 125.205 ;
      RECT 80.185 125.035 80.355 125.205 ;
      RECT 79.725 125.035 79.895 125.205 ;
      RECT 79.265 125.035 79.435 125.205 ;
      RECT 78.805 125.035 78.975 125.205 ;
      RECT 78.345 125.035 78.515 125.205 ;
      RECT 77.885 125.035 78.055 125.205 ;
      RECT 77.425 125.035 77.595 125.205 ;
      RECT 76.965 125.035 77.135 125.205 ;
      RECT 76.505 125.035 76.675 125.205 ;
      RECT 76.045 125.035 76.215 125.205 ;
      RECT 75.585 125.035 75.755 125.205 ;
      RECT 75.125 125.035 75.295 125.205 ;
      RECT 74.665 125.035 74.835 125.205 ;
      RECT 74.205 125.035 74.375 125.205 ;
    LAYER via ;
      RECT 58.805 130.365 58.955 130.515 ;
      RECT 29.365 130.365 29.515 130.515 ;
      RECT 67.775 129.975 67.925 130.125 ;
      RECT 27.295 129.975 27.445 130.125 ;
      RECT 25.455 129.975 25.605 130.125 ;
      RECT 89.395 5.875 89.545 6.025 ;
      RECT 42.015 0.435 42.165 0.585 ;
      RECT 11.655 0.435 11.805 0.585 ;
      RECT 58.805 0.045 58.955 0.195 ;
      RECT 29.365 0.045 29.515 0.195 ;
    LAYER via2 ;
      RECT 58.78 130.34 58.98 130.54 ;
      RECT 29.34 130.34 29.54 130.54 ;
      RECT 73.27 124.68 73.47 124.88 ;
      RECT 102.71 47.16 102.91 47.36 ;
      RECT 94.89 5.68 95.09 5.88 ;
      RECT 58.78 0.02 58.98 0.22 ;
      RECT 29.34 0.02 29.54 0.22 ;
    LAYER via3 ;
      RECT 58.78 130.34 58.98 130.54 ;
      RECT 29.34 130.34 29.54 130.54 ;
      RECT 85.92 5.68 86.12 5.88 ;
      RECT 58.78 0.02 58.98 0.22 ;
      RECT 29.34 0.02 29.54 0.22 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 130.56 73.6 130.56 73.6 125.12 103.96 125.12 103.96 5.44 73.6 5.44 73.6 0 ;
  END
END sb_0__1_

END LIBRARY
