//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module sky130_fd_sc_hd__buf_4
(
    A,
    X
);

    input A;
    output X;

    wire A;
    wire X;

endmodule

