//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module sb_8__8_
(
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
    bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
    bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
    bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
    ccff_head,
    chanx_left_in,
    chany_bottom_in,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_,
    left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
    left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
    left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
    left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
    pReset,
    prog_clk,
    ccff_tail,
    chanx_left_out,
    chany_bottom_out
);

    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
    input bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
    input bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
    input bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
    input bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
    input ccff_head;
    input [0:29]chanx_left_in;
    input [0:29]chany_bottom_in;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_;
    input left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
    input left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
    input left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
    input left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
    input pReset;
    input prog_clk;
    output ccff_tail;
    output [0:29]chanx_left_out;
    output [0:29]chany_bottom_out;

    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
    wire bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
    wire bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
    wire bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
    wire bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
    wire ccff_head;
    wire ccff_tail;
    wire [0:29]chanx_left_in;
    wire [0:29]chanx_left_out;
    wire [0:29]chany_bottom_in;
    wire [0:29]chany_bottom_out;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_;
    wire left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
    wire left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
    wire left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
    wire left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
    wire [0:2]mux_bottom_track_11_undriven_sram_inv;
    wire [0:1]mux_bottom_track_13_undriven_sram_inv;
    wire [0:1]mux_bottom_track_15_undriven_sram_inv;
    wire [0:1]mux_bottom_track_17_undriven_sram_inv;
    wire [0:1]mux_bottom_track_19_undriven_sram_inv;
    wire [0:2]mux_bottom_track_1_undriven_sram_inv;
    wire [0:1]mux_bottom_track_21_undriven_sram_inv;
    wire [0:1]mux_bottom_track_23_undriven_sram_inv;
    wire [0:1]mux_bottom_track_25_undriven_sram_inv;
    wire [0:1]mux_bottom_track_27_undriven_sram_inv;
    wire [0:1]mux_bottom_track_29_undriven_sram_inv;
    wire [0:1]mux_bottom_track_31_undriven_sram_inv;
    wire [0:1]mux_bottom_track_33_undriven_sram_inv;
    wire [0:1]mux_bottom_track_35_undriven_sram_inv;
    wire [0:2]mux_bottom_track_3_undriven_sram_inv;
    wire [0:1]mux_bottom_track_45_undriven_sram_inv;
    wire [0:1]mux_bottom_track_47_undriven_sram_inv;
    wire [0:1]mux_bottom_track_49_undriven_sram_inv;
    wire [0:1]mux_bottom_track_51_undriven_sram_inv;
    wire [0:1]mux_bottom_track_53_undriven_sram_inv;
    wire [0:1]mux_bottom_track_55_undriven_sram_inv;
    wire [0:1]mux_bottom_track_57_undriven_sram_inv;
    wire [0:1]mux_bottom_track_59_undriven_sram_inv;
    wire [0:2]mux_bottom_track_5_undriven_sram_inv;
    wire [0:2]mux_bottom_track_7_undriven_sram_inv;
    wire [0:2]mux_bottom_track_9_undriven_sram_inv;
    wire [0:2]mux_left_track_11_undriven_sram_inv;
    wire [0:1]mux_left_track_13_undriven_sram_inv;
    wire [0:1]mux_left_track_15_undriven_sram_inv;
    wire [0:1]mux_left_track_17_undriven_sram_inv;
    wire [0:1]mux_left_track_19_undriven_sram_inv;
    wire [0:2]mux_left_track_1_undriven_sram_inv;
    wire [0:1]mux_left_track_21_undriven_sram_inv;
    wire [0:1]mux_left_track_23_undriven_sram_inv;
    wire [0:1]mux_left_track_25_undriven_sram_inv;
    wire [0:1]mux_left_track_27_undriven_sram_inv;
    wire [0:1]mux_left_track_29_undriven_sram_inv;
    wire [0:1]mux_left_track_31_undriven_sram_inv;
    wire [0:1]mux_left_track_33_undriven_sram_inv;
    wire [0:1]mux_left_track_35_undriven_sram_inv;
    wire [0:1]mux_left_track_37_undriven_sram_inv;
    wire [0:1]mux_left_track_39_undriven_sram_inv;
    wire [0:2]mux_left_track_3_undriven_sram_inv;
    wire [0:1]mux_left_track_41_undriven_sram_inv;
    wire [0:1]mux_left_track_43_undriven_sram_inv;
    wire [0:1]mux_left_track_45_undriven_sram_inv;
    wire [0:1]mux_left_track_47_undriven_sram_inv;
    wire [0:1]mux_left_track_49_undriven_sram_inv;
    wire [0:1]mux_left_track_51_undriven_sram_inv;
    wire [0:1]mux_left_track_53_undriven_sram_inv;
    wire [0:1]mux_left_track_55_undriven_sram_inv;
    wire [0:1]mux_left_track_57_undriven_sram_inv;
    wire [0:1]mux_left_track_59_undriven_sram_inv;
    wire [0:2]mux_left_track_5_undriven_sram_inv;
    wire [0:2]mux_left_track_7_undriven_sram_inv;
    wire [0:2]mux_left_track_9_undriven_sram_inv;
    wire [0:1]mux_tree_tapbuf_size2_0_sram;
    wire [0:1]mux_tree_tapbuf_size2_10_sram;
    wire [0:1]mux_tree_tapbuf_size2_11_sram;
    wire [0:1]mux_tree_tapbuf_size2_12_sram;
    wire [0:1]mux_tree_tapbuf_size2_13_sram;
    wire [0:1]mux_tree_tapbuf_size2_14_sram;
    wire [0:1]mux_tree_tapbuf_size2_15_sram;
    wire [0:1]mux_tree_tapbuf_size2_16_sram;
    wire [0:1]mux_tree_tapbuf_size2_17_sram;
    wire [0:1]mux_tree_tapbuf_size2_18_sram;
    wire [0:1]mux_tree_tapbuf_size2_19_sram;
    wire [0:1]mux_tree_tapbuf_size2_1_sram;
    wire [0:1]mux_tree_tapbuf_size2_20_sram;
    wire [0:1]mux_tree_tapbuf_size2_21_sram;
    wire [0:1]mux_tree_tapbuf_size2_22_sram;
    wire [0:1]mux_tree_tapbuf_size2_23_sram;
    wire [0:1]mux_tree_tapbuf_size2_24_sram;
    wire [0:1]mux_tree_tapbuf_size2_2_sram;
    wire [0:1]mux_tree_tapbuf_size2_3_sram;
    wire [0:1]mux_tree_tapbuf_size2_4_sram;
    wire [0:1]mux_tree_tapbuf_size2_5_sram;
    wire [0:1]mux_tree_tapbuf_size2_6_sram;
    wire [0:1]mux_tree_tapbuf_size2_7_sram;
    wire [0:1]mux_tree_tapbuf_size2_8_sram;
    wire [0:1]mux_tree_tapbuf_size2_9_sram;
    wire mux_tree_tapbuf_size2_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_10_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_11_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_12_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_13_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_14_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_15_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_16_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_17_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_18_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_19_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_20_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_21_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_22_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_23_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_24_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_2_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_3_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_4_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_5_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_6_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_7_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_8_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_9_ccff_tail;
    wire [0:1]mux_tree_tapbuf_size3_0_sram;
    wire [0:1]mux_tree_tapbuf_size3_10_sram;
    wire [0:1]mux_tree_tapbuf_size3_11_sram;
    wire [0:1]mux_tree_tapbuf_size3_12_sram;
    wire [0:1]mux_tree_tapbuf_size3_13_sram;
    wire [0:1]mux_tree_tapbuf_size3_14_sram;
    wire [0:1]mux_tree_tapbuf_size3_15_sram;
    wire [0:1]mux_tree_tapbuf_size3_16_sram;
    wire [0:1]mux_tree_tapbuf_size3_17_sram;
    wire [0:1]mux_tree_tapbuf_size3_18_sram;
    wire [0:1]mux_tree_tapbuf_size3_1_sram;
    wire [0:1]mux_tree_tapbuf_size3_2_sram;
    wire [0:1]mux_tree_tapbuf_size3_3_sram;
    wire [0:1]mux_tree_tapbuf_size3_4_sram;
    wire [0:1]mux_tree_tapbuf_size3_5_sram;
    wire [0:1]mux_tree_tapbuf_size3_6_sram;
    wire [0:1]mux_tree_tapbuf_size3_7_sram;
    wire [0:1]mux_tree_tapbuf_size3_8_sram;
    wire [0:1]mux_tree_tapbuf_size3_9_sram;
    wire mux_tree_tapbuf_size3_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_10_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_11_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_12_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_13_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_14_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_15_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_16_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_17_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_2_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_3_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_4_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_5_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_6_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_7_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_8_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_9_ccff_tail;
    wire [0:2]mux_tree_tapbuf_size5_0_sram;
    wire [0:2]mux_tree_tapbuf_size5_10_sram;
    wire [0:2]mux_tree_tapbuf_size5_11_sram;
    wire [0:2]mux_tree_tapbuf_size5_1_sram;
    wire [0:2]mux_tree_tapbuf_size5_2_sram;
    wire [0:2]mux_tree_tapbuf_size5_3_sram;
    wire [0:2]mux_tree_tapbuf_size5_4_sram;
    wire [0:2]mux_tree_tapbuf_size5_5_sram;
    wire [0:2]mux_tree_tapbuf_size5_6_sram;
    wire [0:2]mux_tree_tapbuf_size5_7_sram;
    wire [0:2]mux_tree_tapbuf_size5_8_sram;
    wire [0:2]mux_tree_tapbuf_size5_9_sram;
    wire mux_tree_tapbuf_size5_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_10_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_11_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_2_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_3_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_4_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_5_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_6_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_7_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_8_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_9_ccff_tail;
    wire pReset;
    wire prog_clk;

assign chany_bottom_out[18] = chanx_left_in[19];
assign chany_bottom_out[19] = chanx_left_in[20];
assign chany_bottom_out[20] = chanx_left_in[21];
assign chany_bottom_out[21] = chanx_left_in[22];
    mux_tree_tapbuf_size5_mem mem_bottom_track_1
    (
        .ccff_head(ccff_head),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_0_sram)
    );
    mux_tree_tapbuf_size5_mem mem_bottom_track_11
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_5_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_13
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_0_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_15
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_0_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_1_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_17
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_1_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_2_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_19
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_2_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_3_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_3_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_21
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_3_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_4_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_4_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_23
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_4_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_5_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_5_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_25
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_5_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_6_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_6_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_27
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_6_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_7_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_7_sram)
    );
    mux_tree_tapbuf_size3_mem mem_bottom_track_29
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_7_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_0_sram)
    );
    mux_tree_tapbuf_size5_mem mem_bottom_track_3
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_1_sram)
    );
    mux_tree_tapbuf_size3_mem mem_bottom_track_31
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_0_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_1_sram)
    );
    mux_tree_tapbuf_size3_mem mem_bottom_track_33
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_1_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_2_sram)
    );
    mux_tree_tapbuf_size3_mem mem_bottom_track_35
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_2_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_3_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_3_sram)
    );
    mux_tree_tapbuf_size3_mem mem_bottom_track_45
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_3_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_4_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_4_sram)
    );
    mux_tree_tapbuf_size3_mem mem_bottom_track_47
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_4_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_5_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_5_sram)
    );
    mux_tree_tapbuf_size3_mem mem_bottom_track_49
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_5_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_6_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_6_sram)
    );
    mux_tree_tapbuf_size5_mem mem_bottom_track_5
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_2_sram)
    );
    mux_tree_tapbuf_size3_mem mem_bottom_track_51
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_6_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_7_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_7_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_53
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_7_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_8_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_8_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_55
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_8_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_9_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_9_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_57
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_9_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_10_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_10_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_59
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_10_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_11_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_11_sram)
    );
    mux_tree_tapbuf_size5_mem mem_bottom_track_7
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_3_sram)
    );
    mux_tree_tapbuf_size5_mem mem_bottom_track_9
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_4_sram)
    );
    mux_tree_tapbuf_size5_mem mem_left_track_1
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_11_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_6_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_6_sram)
    );
    mux_tree_tapbuf_size5_mem mem_left_track_11
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_10_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_11_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_11_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_13
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_11_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_8_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_8_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_15
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_8_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_9_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_9_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_17
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_9_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_10_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_10_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_19
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_10_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_12_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_12_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_21
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_12_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_13_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_13_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_23
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_13_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_14_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_14_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_25
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_14_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_15_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_15_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_27
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_15_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_16_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_16_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_29
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_16_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_11_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_11_sram)
    );
    mux_tree_tapbuf_size5_mem mem_left_track_3
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_6_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_7_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_7_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_31
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_11_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_12_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_12_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_33
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_12_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_13_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_13_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_35
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_13_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_14_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_14_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_37
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_14_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_17_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_17_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_39
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_17_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_18_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_18_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_41
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_18_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_19_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_19_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_43
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_19_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_20_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_20_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_45
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_20_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_15_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_15_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_47
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_15_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_16_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_16_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_49
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_16_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_17_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_17_sram)
    );
    mux_tree_tapbuf_size5_mem mem_left_track_5
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_7_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_8_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_8_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_51
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_17_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_21_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_21_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_53
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_21_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_22_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_22_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_55
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_22_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_23_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_23_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_57
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_23_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_24_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_24_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_59
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_24_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_18_sram)
    );
    mux_tree_tapbuf_size5_mem mem_left_track_7
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_8_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_9_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_9_sram)
    );
    mux_tree_tapbuf_size5_mem mem_left_track_9
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_9_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_10_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_10_sram)
    );
    mux_tree_tapbuf_size5 mux_bottom_track_1
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[1]}),
        .sram(mux_tree_tapbuf_size5_0_sram),
        .sram_inv(mux_bottom_track_1_undriven_sram_inv),
        .out(chany_bottom_out[0])
    );
    mux_tree_tapbuf_size5 mux_bottom_track_11
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[6]}),
        .sram(mux_tree_tapbuf_size5_5_sram),
        .sram_inv(mux_bottom_track_11_undriven_sram_inv),
        .out(chany_bottom_out[5])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_13
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[7]}),
        .sram(mux_tree_tapbuf_size2_0_sram),
        .sram_inv(mux_bottom_track_13_undriven_sram_inv),
        .out(chany_bottom_out[6])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_15
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[8]}),
        .sram(mux_tree_tapbuf_size2_1_sram),
        .sram_inv(mux_bottom_track_15_undriven_sram_inv),
        .out(chany_bottom_out[7])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_17
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[9]}),
        .sram(mux_tree_tapbuf_size2_2_sram),
        .sram_inv(mux_bottom_track_17_undriven_sram_inv),
        .out(chany_bottom_out[8])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_19
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[10]}),
        .sram(mux_tree_tapbuf_size2_3_sram),
        .sram_inv(mux_bottom_track_19_undriven_sram_inv),
        .out(chany_bottom_out[9])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_21
    (
        .in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[11]}),
        .sram(mux_tree_tapbuf_size2_4_sram),
        .sram_inv(mux_bottom_track_21_undriven_sram_inv),
        .out(chany_bottom_out[10])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_23
    (
        .in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[12]}),
        .sram(mux_tree_tapbuf_size2_5_sram),
        .sram_inv(mux_bottom_track_23_undriven_sram_inv),
        .out(chany_bottom_out[11])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_25
    (
        .in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, chanx_left_in[13]}),
        .sram(mux_tree_tapbuf_size2_6_sram),
        .sram_inv(mux_bottom_track_25_undriven_sram_inv),
        .out(chany_bottom_out[12])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_27
    (
        .in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, chanx_left_in[14]}),
        .sram(mux_tree_tapbuf_size2_7_sram),
        .sram_inv(mux_bottom_track_27_undriven_sram_inv),
        .out(chany_bottom_out[13])
    );
    mux_tree_tapbuf_size3 mux_bottom_track_29
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, chanx_left_in[15]}),
        .sram(mux_tree_tapbuf_size3_0_sram),
        .sram_inv(mux_bottom_track_29_undriven_sram_inv),
        .out(chany_bottom_out[14])
    );
    mux_tree_tapbuf_size5 mux_bottom_track_3
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, chanx_left_in[2]}),
        .sram(mux_tree_tapbuf_size5_1_sram),
        .sram_inv(mux_bottom_track_3_undriven_sram_inv),
        .out(chany_bottom_out[1])
    );
    mux_tree_tapbuf_size3 mux_bottom_track_31
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[16]}),
        .sram(mux_tree_tapbuf_size3_1_sram),
        .sram_inv(mux_bottom_track_31_undriven_sram_inv),
        .out(chany_bottom_out[15])
    );
    mux_tree_tapbuf_size3 mux_bottom_track_33
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, chanx_left_in[17]}),
        .sram(mux_tree_tapbuf_size3_2_sram),
        .sram_inv(mux_bottom_track_33_undriven_sram_inv),
        .out(chany_bottom_out[16])
    );
    mux_tree_tapbuf_size3 mux_bottom_track_35
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[18]}),
        .sram(mux_tree_tapbuf_size3_3_sram),
        .sram_inv(mux_bottom_track_35_undriven_sram_inv),
        .out(chany_bottom_out[17])
    );
    mux_tree_tapbuf_size3 mux_bottom_track_45
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[23]}),
        .sram(mux_tree_tapbuf_size3_4_sram),
        .sram_inv(mux_bottom_track_45_undriven_sram_inv),
        .out(chany_bottom_out[22])
    );
    mux_tree_tapbuf_size3 mux_bottom_track_47
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[24]}),
        .sram(mux_tree_tapbuf_size3_5_sram),
        .sram_inv(mux_bottom_track_47_undriven_sram_inv),
        .out(chany_bottom_out[23])
    );
    mux_tree_tapbuf_size3 mux_bottom_track_49
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, chanx_left_in[25]}),
        .sram(mux_tree_tapbuf_size3_6_sram),
        .sram_inv(mux_bottom_track_49_undriven_sram_inv),
        .out(chany_bottom_out[24])
    );
    mux_tree_tapbuf_size5 mux_bottom_track_5
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[3]}),
        .sram(mux_tree_tapbuf_size5_2_sram),
        .sram_inv(mux_bottom_track_5_undriven_sram_inv),
        .out(chany_bottom_out[2])
    );
    mux_tree_tapbuf_size3 mux_bottom_track_51
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, chanx_left_in[26]}),
        .sram(mux_tree_tapbuf_size3_7_sram),
        .sram_inv(mux_bottom_track_51_undriven_sram_inv),
        .out(chany_bottom_out[25])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_53
    (
        .in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, chanx_left_in[27]}),
        .sram(mux_tree_tapbuf_size2_8_sram),
        .sram_inv(mux_bottom_track_53_undriven_sram_inv),
        .out(chany_bottom_out[26])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_55
    (
        .in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[28]}),
        .sram(mux_tree_tapbuf_size2_9_sram),
        .sram_inv(mux_bottom_track_55_undriven_sram_inv),
        .out(chany_bottom_out[27])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_57
    (
        .in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, chanx_left_in[29]}),
        .sram(mux_tree_tapbuf_size2_10_sram),
        .sram_inv(mux_bottom_track_57_undriven_sram_inv),
        .out(chany_bottom_out[28])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_59
    (
        .in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[0]}),
        .sram(mux_tree_tapbuf_size2_11_sram),
        .sram_inv(mux_bottom_track_59_undriven_sram_inv),
        .out(chany_bottom_out[29])
    );
    mux_tree_tapbuf_size5 mux_bottom_track_7
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[4]}),
        .sram(mux_tree_tapbuf_size5_3_sram),
        .sram_inv(mux_bottom_track_7_undriven_sram_inv),
        .out(chany_bottom_out[3])
    );
    mux_tree_tapbuf_size5 mux_bottom_track_9
    (
        .in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, chanx_left_in[5]}),
        .sram(mux_tree_tapbuf_size5_4_sram),
        .sram_inv(mux_bottom_track_9_undriven_sram_inv),
        .out(chany_bottom_out[4])
    );
    mux_tree_tapbuf_size5 mux_left_track_1
    (
        .in({chany_bottom_in[29], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
        .sram(mux_tree_tapbuf_size5_6_sram),
        .sram_inv(mux_left_track_1_undriven_sram_inv),
        .out(chanx_left_out[0])
    );
    mux_tree_tapbuf_size5 mux_left_track_11
    (
        .in({chany_bottom_in[4], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_}),
        .sram(mux_tree_tapbuf_size5_11_sram),
        .sram_inv(mux_left_track_11_undriven_sram_inv),
        .out(chanx_left_out[5])
    );
    mux_tree_tapbuf_size3 mux_left_track_13
    (
        .in({chany_bottom_in[5], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
        .sram(mux_tree_tapbuf_size3_8_sram),
        .sram_inv(mux_left_track_13_undriven_sram_inv),
        .out(chanx_left_out[6])
    );
    mux_tree_tapbuf_size3 mux_left_track_15
    (
        .in({chany_bottom_in[6], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
        .sram(mux_tree_tapbuf_size3_9_sram),
        .sram_inv(mux_left_track_15_undriven_sram_inv),
        .out(chanx_left_out[7])
    );
    mux_tree_tapbuf_size3 mux_left_track_17
    (
        .in({chany_bottom_in[7], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
        .sram(mux_tree_tapbuf_size3_10_sram),
        .sram_inv(mux_left_track_17_undriven_sram_inv),
        .out(chanx_left_out[8])
    );
    mux_tree_tapbuf_size2 mux_left_track_19
    (
        .in({chany_bottom_in[8], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_12_sram),
        .sram_inv(mux_left_track_19_undriven_sram_inv),
        .out(chanx_left_out[9])
    );
    mux_tree_tapbuf_size2 mux_left_track_21
    (
        .in({chany_bottom_in[9], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
        .sram(mux_tree_tapbuf_size2_13_sram),
        .sram_inv(mux_left_track_21_undriven_sram_inv),
        .out(chanx_left_out[10])
    );
    mux_tree_tapbuf_size2 mux_left_track_23
    (
        .in({chany_bottom_in[10], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_}),
        .sram(mux_tree_tapbuf_size2_14_sram),
        .sram_inv(mux_left_track_23_undriven_sram_inv),
        .out(chanx_left_out[11])
    );
    mux_tree_tapbuf_size2 mux_left_track_25
    (
        .in({chany_bottom_in[11], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
        .sram(mux_tree_tapbuf_size2_15_sram),
        .sram_inv(mux_left_track_25_undriven_sram_inv),
        .out(chanx_left_out[12])
    );
    mux_tree_tapbuf_size2 mux_left_track_27
    (
        .in({chany_bottom_in[12], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_}),
        .sram(mux_tree_tapbuf_size2_16_sram),
        .sram_inv(mux_left_track_27_undriven_sram_inv),
        .out(chanx_left_out[13])
    );
    mux_tree_tapbuf_size3 mux_left_track_29
    (
        .in({chany_bottom_in[13], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
        .sram(mux_tree_tapbuf_size3_11_sram),
        .sram_inv(mux_left_track_29_undriven_sram_inv),
        .out(chanx_left_out[14])
    );
    mux_tree_tapbuf_size5 mux_left_track_3
    (
        .in({chany_bottom_in[0], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
        .sram(mux_tree_tapbuf_size5_7_sram),
        .sram_inv(mux_left_track_3_undriven_sram_inv),
        .out(chanx_left_out[1])
    );
    mux_tree_tapbuf_size3 mux_left_track_31
    (
        .in({chany_bottom_in[14], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
        .sram(mux_tree_tapbuf_size3_12_sram),
        .sram_inv(mux_left_track_31_undriven_sram_inv),
        .out(chanx_left_out[15])
    );
    mux_tree_tapbuf_size3 mux_left_track_33
    (
        .in({chany_bottom_in[15], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
        .sram(mux_tree_tapbuf_size3_13_sram),
        .sram_inv(mux_left_track_33_undriven_sram_inv),
        .out(chanx_left_out[16])
    );
    mux_tree_tapbuf_size3 mux_left_track_35
    (
        .in({chany_bottom_in[16], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_}),
        .sram(mux_tree_tapbuf_size3_14_sram),
        .sram_inv(mux_left_track_35_undriven_sram_inv),
        .out(chanx_left_out[17])
    );
    mux_tree_tapbuf_size2 mux_left_track_37
    (
        .in({chany_bottom_in[17], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
        .sram(mux_tree_tapbuf_size2_17_sram),
        .sram_inv(mux_left_track_37_undriven_sram_inv),
        .out(chanx_left_out[18])
    );
    mux_tree_tapbuf_size2 mux_left_track_39
    (
        .in({chany_bottom_in[18], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_}),
        .sram(mux_tree_tapbuf_size2_18_sram),
        .sram_inv(mux_left_track_39_undriven_sram_inv),
        .out(chanx_left_out[19])
    );
    mux_tree_tapbuf_size2 mux_left_track_41
    (
        .in({chany_bottom_in[19], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
        .sram(mux_tree_tapbuf_size2_19_sram),
        .sram_inv(mux_left_track_41_undriven_sram_inv),
        .out(chanx_left_out[20])
    );
    mux_tree_tapbuf_size2 mux_left_track_43
    (
        .in({chany_bottom_in[20], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_}),
        .sram(mux_tree_tapbuf_size2_20_sram),
        .sram_inv(mux_left_track_43_undriven_sram_inv),
        .out(chanx_left_out[21])
    );
    mux_tree_tapbuf_size3 mux_left_track_45
    (
        .in({chany_bottom_in[21], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
        .sram(mux_tree_tapbuf_size3_15_sram),
        .sram_inv(mux_left_track_45_undriven_sram_inv),
        .out(chanx_left_out[22])
    );
    mux_tree_tapbuf_size3 mux_left_track_47
    (
        .in({chany_bottom_in[22], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
        .sram(mux_tree_tapbuf_size3_16_sram),
        .sram_inv(mux_left_track_47_undriven_sram_inv),
        .out(chanx_left_out[23])
    );
    mux_tree_tapbuf_size3 mux_left_track_49
    (
        .in({chany_bottom_in[23], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
        .sram(mux_tree_tapbuf_size3_17_sram),
        .sram_inv(mux_left_track_49_undriven_sram_inv),
        .out(chanx_left_out[24])
    );
    mux_tree_tapbuf_size5 mux_left_track_5
    (
        .in({chany_bottom_in[1], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_}),
        .sram(mux_tree_tapbuf_size5_8_sram),
        .sram_inv(mux_left_track_5_undriven_sram_inv),
        .out(chanx_left_out[2])
    );
    mux_tree_tapbuf_size2 mux_left_track_51
    (
        .in({chany_bottom_in[24], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_21_sram),
        .sram_inv(mux_left_track_51_undriven_sram_inv),
        .out(chanx_left_out[25])
    );
    mux_tree_tapbuf_size2 mux_left_track_53
    (
        .in({chany_bottom_in[25], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
        .sram(mux_tree_tapbuf_size2_22_sram),
        .sram_inv(mux_left_track_53_undriven_sram_inv),
        .out(chanx_left_out[26])
    );
    mux_tree_tapbuf_size2 mux_left_track_55
    (
        .in({chany_bottom_in[26], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_}),
        .sram(mux_tree_tapbuf_size2_23_sram),
        .sram_inv(mux_left_track_55_undriven_sram_inv),
        .out(chanx_left_out[27])
    );
    mux_tree_tapbuf_size2 mux_left_track_57
    (
        .in({chany_bottom_in[27], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
        .sram(mux_tree_tapbuf_size2_24_sram),
        .sram_inv(mux_left_track_57_undriven_sram_inv),
        .out(chanx_left_out[28])
    );
    mux_tree_tapbuf_size3 mux_left_track_59
    (
        .in({chany_bottom_in[28], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_}),
        .sram(mux_tree_tapbuf_size3_18_sram),
        .sram_inv(mux_left_track_59_undriven_sram_inv),
        .out(chanx_left_out[29])
    );
    mux_tree_tapbuf_size5 mux_left_track_7
    (
        .in({chany_bottom_in[2], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
        .sram(mux_tree_tapbuf_size5_9_sram),
        .sram_inv(mux_left_track_7_undriven_sram_inv),
        .out(chanx_left_out[3])
    );
    mux_tree_tapbuf_size5 mux_left_track_9
    (
        .in({chany_bottom_in[3], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
        .sram(mux_tree_tapbuf_size5_10_sram),
        .sram_inv(mux_left_track_9_undriven_sram_inv),
        .out(chanx_left_out[4])
    );
endmodule

