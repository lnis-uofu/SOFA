VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_1__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 134.32 BY 130.56 ;
  SYMMETRY X Y ;
  PIN pReset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.04 130.075 59.18 130.56 ;
    END
  END pReset[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 75.75 129.76 76.05 130.56 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 79.43 129.76 79.73 130.56 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.1 130.075 87.24 130.56 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.79 129.76 87.09 130.56 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.79 129.76 64.09 130.56 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71 130.075 71.14 130.56 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.62 130.075 92.76 130.56 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.59 129.76 77.89 130.56 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.23 129.76 70.53 130.56 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.66 130.075 34.8 130.56 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 130.075 35.72 130.56 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.84 130.075 95.98 130.56 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.58 130.075 81.72 130.56 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.36 130.075 78.5 130.56 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.95 129.76 62.25 130.56 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.07 129.76 72.37 130.56 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.18 130.075 86.32 130.56 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94 130.075 94.14 130.56 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.11 129.76 83.41 130.56 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.2 130.075 80.34 130.56 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.02 130.075 42.16 130.56 ;
    END
  END chany_top_in[20]
  PIN chany_top_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 65.63 129.76 65.93 130.56 ;
    END
  END chany_top_in[21]
  PIN chany_top_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.39 129.76 68.69 130.56 ;
    END
  END chany_top_in[22]
  PIN chany_top_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.42 130.075 83.56 130.56 ;
    END
  END chany_top_in[23]
  PIN chany_top_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.27 129.76 81.57 130.56 ;
    END
  END chany_top_in[24]
  PIN chany_top_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.95 129.76 85.25 130.56 ;
    END
  END chany_top_in[25]
  PIN chany_top_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.02 130.075 88.16 130.56 ;
    END
  END chany_top_in[26]
  PIN chany_top_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.86 130.075 90 130.56 ;
    END
  END chany_top_in[27]
  PIN chany_top_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.7 130.075 91.84 130.56 ;
    END
  END chany_top_in[28]
  PIN chany_top_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.5 130.075 82.64 130.56 ;
    END
  END chany_top_in[29]
  PIN top_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.18 124.635 17.32 125.12 ;
    END
  END top_left_grid_pin_44_[0]
  PIN top_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.12 124.635 12.26 125.12 ;
    END
  END top_left_grid_pin_45_[0]
  PIN top_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.02 124.635 19.16 125.12 ;
    END
  END top_left_grid_pin_46_[0]
  PIN top_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.4 124.635 20.54 125.12 ;
    END
  END top_left_grid_pin_47_[0]
  PIN top_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.84 124.635 3.98 125.12 ;
    END
  END top_left_grid_pin_48_[0]
  PIN top_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.42 124.635 14.56 125.12 ;
    END
  END top_left_grid_pin_49_[0]
  PIN top_left_grid_pin_50_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.2 124.635 11.34 125.12 ;
    END
  END top_left_grid_pin_50_[0]
  PIN top_left_grid_pin_51_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.1 124.635 18.24 125.12 ;
    END
  END top_left_grid_pin_51_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 47.11 134.32 47.41 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 60.71 134.32 61.01 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 67.51 134.32 67.81 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 45.75 134.32 46.05 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 37.16 134.32 37.3 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 34.1 134.32 34.24 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 52.46 134.32 52.6 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 44.39 134.32 44.69 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 59.35 134.32 59.65 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 26.71 134.32 27.01 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 15.4 134.32 15.54 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 44.64 134.32 44.78 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 58.24 134.32 58.38 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 64.79 134.32 65.09 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 42.6 134.32 42.74 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 50.42 134.32 50.56 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 14.72 134.32 14.86 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 39.88 134.32 40.02 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 41.92 134.32 42.06 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 62.07 134.32 62.37 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 33.42 134.32 33.56 ;
    END
  END chanx_right_in[20]
  PIN chanx_right_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 23.99 134.32 24.29 ;
    END
  END chanx_right_in[21]
  PIN chanx_right_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 47.02 134.32 47.16 ;
    END
  END chanx_right_in[22]
  PIN chanx_right_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 45.32 134.32 45.46 ;
    END
  END chanx_right_in[23]
  PIN chanx_right_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 63.68 134.32 63.82 ;
    END
  END chanx_right_in[24]
  PIN chanx_right_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 49.74 134.32 49.88 ;
    END
  END chanx_right_in[25]
  PIN chanx_right_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 39.2 134.32 39.34 ;
    END
  END chanx_right_in[26]
  PIN chanx_right_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 21.27 134.32 21.57 ;
    END
  END chanx_right_in[27]
  PIN chanx_right_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 36.48 134.32 36.62 ;
    END
  END chanx_right_in[28]
  PIN chanx_right_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 47.7 134.32 47.84 ;
    END
  END chanx_right_in[29]
  PIN right_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.36 5.44 124.5 5.925 ;
    END
  END right_bottom_grid_pin_36_[0]
  PIN right_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.12 5.44 127.26 5.925 ;
    END
  END right_bottom_grid_pin_37_[0]
  PIN right_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.2 5.44 126.34 5.925 ;
    END
  END right_bottom_grid_pin_38_[0]
  PIN right_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.28 5.44 125.42 5.925 ;
    END
  END right_bottom_grid_pin_39_[0]
  PIN right_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.76 5.44 119.9 5.925 ;
    END
  END right_bottom_grid_pin_40_[0]
  PIN right_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.68 5.44 120.82 5.925 ;
    END
  END right_bottom_grid_pin_41_[0]
  PIN right_bottom_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.44 5.44 123.58 5.925 ;
    END
  END right_bottom_grid_pin_42_[0]
  PIN right_bottom_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.6 5.44 121.74 5.925 ;
    END
  END right_bottom_grid_pin_43_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.23 0 70.53 0.8 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.47 0 90.77 0.8 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.55 0 66.85 0.8 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.31 0 92.61 0.8 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.79 0 87.09 0.8 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.87 0 63.17 0.8 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.04 0 59.18 0.485 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.72 0 39.86 0.485 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.62 0 92.76 0.485 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.6 0 75.74 0.485 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 75.75 0 76.05 0.8 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.07 0 72.37 0.8 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.99 0 96.29 0.8 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.22 0 97.36 0.485 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.46 0 94.6 0.485 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.52 0 76.66 0.485 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 64.71 0 65.01 0.8 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.03 0 61.33 0.8 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.15 0 94.45 0.8 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.27 0 81.57 0.8 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.3 0 96.44 0.485 ;
    END
  END chany_bottom_in[20]
  PIN chany_bottom_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.38 0 95.52 0.485 ;
    END
  END chany_bottom_in[21]
  PIN chany_bottom_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.64 0 40.78 0.485 ;
    END
  END chany_bottom_in[22]
  PIN chany_bottom_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.68 0 74.82 0.485 ;
    END
  END chany_bottom_in[23]
  PIN chany_bottom_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.83 0 98.13 0.8 ;
    END
  END chany_bottom_in[24]
  PIN chany_bottom_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.2 0 80.34 0.485 ;
    END
  END chany_bottom_in[25]
  PIN chany_bottom_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.39 0 68.69 0.8 ;
    END
  END chany_bottom_in[26]
  PIN chany_bottom_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.78 0 90.92 0.485 ;
    END
  END chany_bottom_in[27]
  PIN chany_bottom_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.59 0 77.89 0.8 ;
    END
  END chany_bottom_in[28]
  PIN chany_bottom_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 79.43 0 79.73 0.8 ;
    END
  END chany_bottom_in[29]
  PIN bottom_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.72 5.44 16.86 5.925 ;
    END
  END bottom_left_grid_pin_44_[0]
  PIN bottom_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.84 5.44 3.98 5.925 ;
    END
  END bottom_left_grid_pin_45_[0]
  PIN bottom_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.56 5.44 18.7 5.925 ;
    END
  END bottom_left_grid_pin_46_[0]
  PIN bottom_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.64 5.44 17.78 5.925 ;
    END
  END bottom_left_grid_pin_47_[0]
  PIN bottom_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.28 5.44 10.42 5.925 ;
    END
  END bottom_left_grid_pin_48_[0]
  PIN bottom_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.5 5.44 13.64 5.925 ;
    END
  END bottom_left_grid_pin_49_[0]
  PIN bottom_left_grid_pin_50_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.34 5.44 15.48 5.925 ;
    END
  END bottom_left_grid_pin_50_[0]
  PIN bottom_left_grid_pin_51_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.42 5.44 14.56 5.925 ;
    END
  END bottom_left_grid_pin_51_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 39.2 0.595 39.34 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.39 0.8 44.69 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 64.79 0.8 65.09 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.47 0.8 48.77 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 53.91 0.8 54.21 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 12.68 0.595 12.82 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 64.36 0.595 64.5 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 41.92 0.595 42.06 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 52.46 0.595 52.6 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 67.51 0.8 67.81 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 58.24 0.595 58.38 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 55.18 0.595 55.32 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 62.07 0.8 62.37 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 39.88 0.595 40.02 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 49.83 0.8 50.13 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.03 0.8 43.33 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 55.27 0.8 55.57 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 37.16 0.595 37.3 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 66.15 0.8 66.45 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 47.11 0.8 47.41 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 60.71 0.8 61.01 ;
    END
  END chanx_left_in[20]
  PIN chanx_left_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 61.64 0.595 61.78 ;
    END
  END chanx_left_in[21]
  PIN chanx_left_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 58.92 0.595 59.06 ;
    END
  END chanx_left_in[22]
  PIN chanx_left_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 49.74 0.595 49.88 ;
    END
  END chanx_left_in[23]
  PIN chanx_left_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 63.43 0.8 63.73 ;
    END
  END chanx_left_in[24]
  PIN chanx_left_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 47.7 0.595 47.84 ;
    END
  END chanx_left_in[25]
  PIN chanx_left_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 50.42 0.595 50.56 ;
    END
  END chanx_left_in[26]
  PIN chanx_left_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 55.86 0.595 56 ;
    END
  END chanx_left_in[27]
  PIN chanx_left_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.35 0.8 59.65 ;
    END
  END chanx_left_in[28]
  PIN chanx_left_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 45.75 0.8 46.05 ;
    END
  END chanx_left_in[29]
  PIN left_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.12 5.44 12.26 5.925 ;
    END
  END left_bottom_grid_pin_36_[0]
  PIN left_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 7.24 0.595 7.38 ;
    END
  END left_bottom_grid_pin_37_[0]
  PIN left_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.36 5.44 9.5 5.925 ;
    END
  END left_bottom_grid_pin_38_[0]
  PIN left_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.44 5.44 8.58 5.925 ;
    END
  END left_bottom_grid_pin_39_[0]
  PIN left_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.52 5.44 7.66 5.925 ;
    END
  END left_bottom_grid_pin_40_[0]
  PIN left_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.92 5.44 3.06 5.925 ;
    END
  END left_bottom_grid_pin_41_[0]
  PIN left_bottom_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.2 5.44 11.34 5.925 ;
    END
  END left_bottom_grid_pin_42_[0]
  PIN left_bottom_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 8.94 0.595 9.08 ;
    END
  END left_bottom_grid_pin_43_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 66.4 134.32 66.54 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.52 130.075 76.66 130.56 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.24 130.075 45.38 130.56 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 130.075 41.24 130.56 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.28 130.075 79.42 130.56 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48 130.075 48.14 130.56 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.8 130.075 61.94 130.56 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.6 130.075 75.74 130.56 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.68 130.075 74.82 130.56 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.64 130.075 63.78 130.56 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.16 130.075 69.3 130.56 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.24 130.075 68.38 130.56 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.4 130.075 66.54 130.56 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.72 130.075 62.86 130.56 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.84 130.075 49.98 130.56 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.88 130.075 61.02 130.56 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.08 130.075 70.22 130.56 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.16 130.075 46.3 130.56 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.56 130.075 64.7 130.56 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.92 130.075 72.06 130.56 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.92 130.075 49.06 130.56 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.31 129.76 92.61 130.56 ;
    END
  END chany_top_out[20]
  PIN chany_top_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.44 130.075 77.58 130.56 ;
    END
  END chany_top_out[21]
  PIN chany_top_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.08 130.075 47.22 130.56 ;
    END
  END chany_top_out[22]
  PIN chany_top_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.42 130.075 37.56 130.56 ;
    END
  END chany_top_out[23]
  PIN chany_top_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.92 130.075 95.06 130.56 ;
    END
  END chany_top_out[24]
  PIN chany_top_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.32 130.075 44.46 130.56 ;
    END
  END chany_top_out[25]
  PIN chany_top_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.48 130.075 65.62 130.56 ;
    END
  END chany_top_out[26]
  PIN chany_top_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.8 130.075 38.94 130.56 ;
    END
  END chany_top_out[27]
  PIN chany_top_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.32 130.075 67.46 130.56 ;
    END
  END chany_top_out[28]
  PIN chany_top_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.4 130.075 43.54 130.56 ;
    END
  END chany_top_out[29]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 61.64 134.32 61.78 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 20.16 134.32 20.3 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 27.98 134.32 28.12 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 64.36 134.32 64.5 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 25.35 134.32 25.65 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 30.7 134.32 30.84 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 66.15 134.32 66.45 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 13.79 134.32 14.09 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 22.63 134.32 22.93 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 58.92 134.32 59.06 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 56.2 134.32 56.34 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 18.12 134.32 18.26 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 60.96 134.32 61.1 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 12.43 134.32 12.73 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 31.38 134.32 31.52 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 55.52 134.32 55.66 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 11.07 134.32 11.37 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 22.88 134.32 23.02 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.52 63.43 134.32 63.73 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 11.66 134.32 11.8 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 17.44 134.32 17.58 ;
    END
  END chanx_right_out[20]
  PIN chanx_right_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 67.08 134.32 67.22 ;
    END
  END chanx_right_out[21]
  PIN chanx_right_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 20.84 134.32 20.98 ;
    END
  END chanx_right_out[22]
  PIN chanx_right_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 25.26 134.32 25.4 ;
    END
  END chanx_right_out[23]
  PIN chanx_right_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 88.84 134.32 88.98 ;
    END
  END chanx_right_out[24]
  PIN chanx_right_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 12.34 134.32 12.48 ;
    END
  END chanx_right_out[25]
  PIN chanx_right_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 28.66 134.32 28.8 ;
    END
  END chanx_right_out[26]
  PIN chanx_right_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 53.48 134.32 53.62 ;
    END
  END chanx_right_out[27]
  PIN chanx_right_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 25.94 134.32 26.08 ;
    END
  END chanx_right_out[28]
  PIN chanx_right_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 23.56 134.32 23.7 ;
    END
  END chanx_right_out[29]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.18 0 86.32 0.485 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.32 0 44.46 0.485 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.48 0 42.62 0.485 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.54 0 93.68 0.485 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.12 0 81.26 0.485 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.16 0 46.3 0.485 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.46 0 71.6 0.485 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48 0 48.14 0.485 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.08 0 47.22 0.485 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.32 0 67.46 0.485 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.4 0 66.54 0.485 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.7 0 91.84 0.485 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.02 0 88.16 0.485 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.28 0 79.42 0.485 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.56 0 64.7 0.485 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.7 0 68.84 0.485 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.54 0 70.68 0.485 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.48 0 65.62 0.485 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.36 0 78.5 0.485 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.44 0 77.58 0.485 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.86 0 90 0.485 ;
    END
  END chany_bottom_out[20]
  PIN chany_bottom_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.8 0 61.94 0.485 ;
    END
  END chany_bottom_out[21]
  PIN chany_bottom_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.4 0 43.54 0.485 ;
    END
  END chany_bottom_out[22]
  PIN chany_bottom_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.88 0 61.02 0.485 ;
    END
  END chany_bottom_out[23]
  PIN chany_bottom_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.1 0 87.24 0.485 ;
    END
  END chany_bottom_out[24]
  PIN chany_bottom_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.72 0 62.86 0.485 ;
    END
  END chany_bottom_out[25]
  PIN chany_bottom_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.64 0 63.78 0.485 ;
    END
  END chany_bottom_out[26]
  PIN chany_bottom_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.92 0 49.06 0.485 ;
    END
  END chany_bottom_out[27]
  PIN chany_bottom_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.62 0 69.76 0.485 ;
    END
  END chany_bottom_out[28]
  PIN chany_bottom_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.24 0 45.38 0.485 ;
    END
  END chany_bottom_out[29]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 47.02 0.595 47.16 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 15.4 0.595 15.54 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 18.12 0.595 18.26 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 44.64 0.595 44.78 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 17.44 0.595 17.58 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 28.66 0.595 28.8 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 23.99 0.8 24.29 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 11.66 0.595 11.8 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 30.7 0.595 30.84 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 57.99 0.8 58.29 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 27.98 0.595 28.12 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 14.72 0.595 14.86 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.63 0.8 56.93 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 11.07 0.8 11.37 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 22.88 0.595 23.02 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 60.96 0.595 61.1 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 25.94 0.595 26.08 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 25.26 0.595 25.4 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 66.4 0.595 66.54 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 13.79 0.8 14.09 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 36.14 0.595 36.28 ;
    END
  END chanx_left_out[20]
  PIN chanx_left_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 67.08 0.595 67.22 ;
    END
  END chanx_left_out[21]
  PIN chanx_left_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 42.6 0.595 42.74 ;
    END
  END chanx_left_out[22]
  PIN chanx_left_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 23.56 0.595 23.7 ;
    END
  END chanx_left_out[23]
  PIN chanx_left_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 88.84 0.595 88.98 ;
    END
  END chanx_left_out[24]
  PIN chanx_left_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 12.43 0.8 12.73 ;
    END
  END chanx_left_out[25]
  PIN chanx_left_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 20.16 0.595 20.3 ;
    END
  END chanx_left_out[26]
  PIN chanx_left_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 63.68 0.595 63.82 ;
    END
  END chanx_left_out[27]
  PIN chanx_left_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 20.84 0.595 20.98 ;
    END
  END chanx_left_out[28]
  PIN chanx_left_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 31.38 0.595 31.52 ;
    END
  END chanx_left_out[29]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 45.32 0.595 45.46 ;
    END
  END ccff_tail[0]
  PIN Test_en_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.5 0 82.64 0.485 ;
    END
  END Test_en_S_in
  PIN Test_en_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.34 130.075 84.48 130.56 ;
    END
  END Test_en_N_out
  PIN pReset_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.56 0 41.7 0.485 ;
    END
  END pReset_S_in
  PIN pReset_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 80.34 134.32 80.48 ;
    END
  END pReset_E_in
  PIN pReset_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 79.66 0.595 79.8 ;
    END
  END pReset_W_in
  PIN pReset_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.72 130.075 39.86 130.56 ;
    END
  END pReset_N_out
  PIN pReset_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 53.14 0.595 53.28 ;
    END
  END pReset_W_out
  PIN pReset_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 102.1 134.32 102.24 ;
    END
  END pReset_E_out
  PIN Reset_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.42 0 83.56 0.485 ;
    END
  END Reset_S_in
  PIN Reset_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.26 130.075 85.4 130.56 ;
    END
  END Reset_N_out
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 36.5 130.075 36.64 130.56 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_1_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.76 130.075 73.9 130.56 ;
    END
  END prog_clk_1_N_in
  PIN prog_clk_1_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.76 0 73.9 0.485 ;
    END
  END prog_clk_1_S_in
  PIN prog_clk_1_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 79.66 134.32 79.8 ;
    END
  END prog_clk_1_E_out
  PIN prog_clk_1_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 34.44 0.595 34.58 ;
    END
  END prog_clk_1_W_out
  PIN prog_clk_2_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.06 130.075 99.2 130.56 ;
    END
  END prog_clk_2_N_in
  PIN prog_clk_2_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 115.7 134.32 115.84 ;
    END
  END prog_clk_2_E_in
  PIN prog_clk_2_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.34 0 84.48 0.485 ;
    END
  END prog_clk_2_S_in
  PIN prog_clk_2_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 115.02 0.595 115.16 ;
    END
  END prog_clk_2_W_in
  PIN prog_clk_2_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 121.48 0.595 121.62 ;
    END
  END prog_clk_2_W_out
  PIN prog_clk_2_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.14 0 98.28 0.485 ;
    END
  END prog_clk_2_S_out
  PIN prog_clk_2_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.22 130.075 97.36 130.56 ;
    END
  END prog_clk_2_N_out
  PIN prog_clk_2_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 117.74 134.32 117.88 ;
    END
  END prog_clk_2_E_out
  PIN prog_clk_3_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 109.92 0.595 110.06 ;
    END
  END prog_clk_3_W_in
  PIN prog_clk_3_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 109.92 134.32 110.06 ;
    END
  END prog_clk_3_E_in
  PIN prog_clk_3_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.11 0 83.41 0.8 ;
    END
  END prog_clk_3_S_in
  PIN prog_clk_3_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.75 129.76 99.05 130.56 ;
    END
  END prog_clk_3_N_in
  PIN prog_clk_3_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 107.2 134.32 107.34 ;
    END
  END prog_clk_3_E_out
  PIN prog_clk_3_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 118.42 0.595 118.56 ;
    END
  END prog_clk_3_W_out
  PIN prog_clk_3_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.14 130.075 98.28 130.56 ;
    END
  END prog_clk_3_N_out
  PIN prog_clk_3_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.06 0 99.2 0.485 ;
    END
  END prog_clk_3_S_out
  PIN clk_1_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.84 130.075 72.98 130.56 ;
    END
  END clk_1_N_in
  PIN clk_1_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.84 0 72.98 0.485 ;
    END
  END clk_1_S_in
  PIN clk_1_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 101.42 134.32 101.56 ;
    END
  END clk_1_E_out
  PIN clk_1_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 33.76 0.595 33.9 ;
    END
  END clk_1_W_out
  PIN clk_2_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.47 129.76 90.77 130.56 ;
    END
  END clk_2_N_in
  PIN clk_2_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 113.32 134.32 113.46 ;
    END
  END clk_2_E_in
  PIN clk_2_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.26 0 85.4 0.485 ;
    END
  END clk_2_S_in
  PIN clk_2_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 110.6 0.595 110.74 ;
    END
  END clk_2_W_in
  PIN clk_2_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 112.98 0.595 113.12 ;
    END
  END clk_2_W_out
  PIN clk_2_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.98 0 100.12 0.485 ;
    END
  END clk_2_S_out
  PIN clk_2_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.98 130.075 100.12 130.56 ;
    END
  END clk_2_N_out
  PIN clk_2_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 110.6 134.32 110.74 ;
    END
  END clk_2_E_out
  PIN clk_3_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 112.3 0.595 112.44 ;
    END
  END clk_3_W_in
  PIN clk_3_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 112.3 134.32 112.44 ;
    END
  END clk_3_E_in
  PIN clk_3_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.95 0 85.25 0.8 ;
    END
  END clk_3_S_in
  PIN clk_3_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.78 130.075 90.92 130.56 ;
    END
  END clk_3_N_in
  PIN clk_3_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 133.725 107.88 134.32 108.02 ;
    END
  END clk_3_E_out
  PIN clk_3_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 120.46 0.595 120.6 ;
    END
  END clk_3_W_out
  PIN clk_3_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.36 130.075 101.5 130.56 ;
    END
  END clk_3_N_out
  PIN clk_3_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.36 0 101.5 0.485 ;
    END
  END clk_3_S_out
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 22.88 3.2 26.08 ;
        RECT 131.12 22.88 134.32 26.08 ;
        RECT 0 63.68 3.2 66.88 ;
        RECT 131.12 63.68 134.32 66.88 ;
        RECT 0 104.48 3.2 107.68 ;
        RECT 131.12 104.48 134.32 107.68 ;
      LAYER met4 ;
        RECT 44.78 0 45.38 0.6 ;
        RECT 74.22 0 74.82 0.6 ;
        RECT 13.5 5.44 14.1 6.04 ;
        RECT 120.22 5.44 120.82 6.04 ;
        RECT 13.5 124.52 14.1 125.12 ;
        RECT 120.22 124.52 120.82 125.12 ;
        RECT 44.78 129.96 45.38 130.56 ;
        RECT 74.22 129.96 74.82 130.56 ;
      LAYER met1 ;
        RECT 30.36 2.48 30.84 2.96 ;
        RECT 103.48 2.48 103.96 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 133.84 7.92 134.32 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 133.84 13.36 134.32 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 133.84 18.8 134.32 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 133.84 24.24 134.32 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 133.84 29.68 134.32 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 133.84 35.12 134.32 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 133.84 40.56 134.32 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 133.84 46 134.32 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 133.84 51.44 134.32 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 133.84 56.88 134.32 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 133.84 62.32 134.32 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 133.84 67.76 134.32 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 133.84 73.2 134.32 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 133.84 78.64 134.32 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 133.84 84.08 134.32 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 133.84 89.52 134.32 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 133.84 94.96 134.32 95.44 ;
        RECT 0 100.4 0.48 100.88 ;
        RECT 133.84 100.4 134.32 100.88 ;
        RECT 0 105.84 0.48 106.32 ;
        RECT 133.84 105.84 134.32 106.32 ;
        RECT 0 111.28 0.48 111.76 ;
        RECT 133.84 111.28 134.32 111.76 ;
        RECT 0 116.72 0.48 117.2 ;
        RECT 133.84 116.72 134.32 117.2 ;
        RECT 0 122.16 0.48 122.64 ;
        RECT 133.84 122.16 134.32 122.64 ;
        RECT 30.36 127.6 30.84 128.08 ;
        RECT 103.48 127.6 103.96 128.08 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 43.28 3.2 46.48 ;
        RECT 131.12 43.28 134.32 46.48 ;
        RECT 0 84.08 3.2 87.28 ;
        RECT 131.12 84.08 134.32 87.28 ;
      LAYER met4 ;
        RECT 59.5 0 60.1 0.6 ;
        RECT 88.94 0 89.54 0.6 ;
        RECT 59.5 129.96 60.1 130.56 ;
        RECT 88.94 129.96 89.54 130.56 ;
      LAYER met1 ;
        RECT 30.36 -0.24 30.84 0.24 ;
        RECT 103.48 -0.24 103.96 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 133.84 5.2 134.32 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 133.84 10.64 134.32 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 133.84 16.08 134.32 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 133.84 21.52 134.32 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 133.84 26.96 134.32 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 133.84 32.4 134.32 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 133.84 37.84 134.32 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 133.84 43.28 134.32 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 133.84 48.72 134.32 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 133.84 54.16 134.32 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 133.84 59.6 134.32 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 133.84 65.04 134.32 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 133.84 70.48 134.32 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 133.84 75.92 134.32 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 133.84 81.36 134.32 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 133.84 86.8 134.32 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 133.84 92.24 134.32 92.72 ;
        RECT 0 97.68 0.48 98.16 ;
        RECT 133.84 97.68 134.32 98.16 ;
        RECT 0 103.12 0.48 103.6 ;
        RECT 133.84 103.12 134.32 103.6 ;
        RECT 0 108.56 0.48 109.04 ;
        RECT 133.84 108.56 134.32 109.04 ;
        RECT 0 114 0.48 114.48 ;
        RECT 133.84 114 134.32 114.48 ;
        RECT 0 119.44 0.48 119.92 ;
        RECT 133.84 119.44 134.32 119.92 ;
        RECT 0 124.88 0.48 125.36 ;
        RECT 133.84 124.88 134.32 125.36 ;
        RECT 30.36 130.32 30.84 130.8 ;
        RECT 103.48 130.32 103.96 130.8 ;
    END
  END VSS
  OBS
    LAYER met2 ;
      RECT 89.1 130.255 89.38 130.625 ;
      RECT 59.66 130.255 59.94 130.625 ;
      POLYGON 75.28 130.46 75.28 121.31 75.14 121.31 75.14 130.32 75.1 130.32 75.1 130.46 ;
      POLYGON 84.09 130.405 84.09 130.035 84.02 130.035 84.02 129.87 84.08 129.87 84.08 129.55 83.82 129.55 83.82 129.87 83.88 129.87 83.88 130.035 83.81 130.035 83.81 130.405 ;
      POLYGON 70.75 130.405 70.75 130.035 70.68 130.035 70.68 126.24 70.54 126.24 70.54 130.035 70.47 130.035 70.47 130.405 ;
      RECT 34.14 129.55 34.4 129.87 ;
      RECT 17.58 124.45 17.84 124.77 ;
      POLYGON 1.22 80.14 1.22 80 0.3 80 0.3 50.05 2.14 50.05 2.14 49.91 0.16 49.91 0.16 80.14 ;
      POLYGON 86.78 11.46 86.78 0.525 86.85 0.525 86.85 0.155 86.57 0.155 86.57 0.525 86.64 0.525 86.64 11.46 ;
      POLYGON 109.32 9.76 109.32 5.965 109.39 5.965 109.39 5.595 109.11 5.595 109.11 5.965 109.18 5.965 109.18 9.76 ;
      POLYGON 67 8.74 67 0.24 67.04 0.24 67.04 0.1 66.86 0.1 66.86 8.74 ;
      RECT 127.52 6.13 127.78 6.45 ;
      RECT 18.96 6.13 19.22 6.45 ;
      RECT 10.68 6.13 10.94 6.45 ;
      RECT 124.76 5.79 125.02 6.11 ;
      RECT 122 5.79 122.26 6.11 ;
      RECT 12.52 5.79 12.78 6.11 ;
      POLYGON 95.98 1.26 95.98 0.525 96.05 0.525 96.05 0.155 95.77 0.155 95.77 0.525 95.84 0.525 95.84 1.26 ;
      POLYGON 64.24 1.26 64.24 0.525 64.31 0.525 64.31 0.155 64.03 0.155 64.03 0.525 64.1 0.525 64.1 1.26 ;
      RECT 94.86 0.69 95.12 1.01 ;
      RECT 91.18 0.69 91.44 1.01 ;
      RECT 41.96 0.69 42.22 1.01 ;
      RECT 89.1 -0.065 89.38 0.305 ;
      RECT 59.66 -0.065 59.94 0.305 ;
      POLYGON 103.68 130.28 103.68 124.84 134.04 124.84 134.04 5.72 127.54 5.72 127.54 6.205 126.84 6.205 126.84 5.72 126.62 5.72 126.62 6.205 125.92 6.205 125.92 5.72 125.7 5.72 125.7 6.205 125 6.205 125 5.72 124.78 5.72 124.78 6.205 124.08 6.205 124.08 5.72 123.86 5.72 123.86 6.205 123.16 6.205 123.16 5.72 122.02 5.72 122.02 6.205 121.32 6.205 121.32 5.72 121.1 5.72 121.1 6.205 120.4 6.205 120.4 5.72 120.18 5.72 120.18 6.205 119.48 6.205 119.48 5.72 103.68 5.72 103.68 0.28 101.78 0.28 101.78 0.765 101.08 0.765 101.08 0.28 100.4 0.28 100.4 0.765 99.7 0.765 99.7 0.28 99.48 0.28 99.48 0.765 98.78 0.765 98.78 0.28 98.56 0.28 98.56 0.765 97.86 0.765 97.86 0.28 97.64 0.28 97.64 0.765 96.94 0.765 96.94 0.28 96.72 0.28 96.72 0.765 96.02 0.765 96.02 0.28 95.8 0.28 95.8 0.765 95.1 0.765 95.1 0.28 94.88 0.28 94.88 0.765 94.18 0.765 94.18 0.28 93.96 0.28 93.96 0.765 93.26 0.765 93.26 0.28 93.04 0.28 93.04 0.765 92.34 0.765 92.34 0.28 92.12 0.28 92.12 0.765 91.42 0.765 91.42 0.28 91.2 0.28 91.2 0.765 90.5 0.765 90.5 0.28 90.28 0.28 90.28 0.765 89.58 0.765 89.58 0.28 88.44 0.28 88.44 0.765 87.74 0.765 87.74 0.28 87.52 0.28 87.52 0.765 86.82 0.765 86.82 0.28 86.6 0.28 86.6 0.765 85.9 0.765 85.9 0.28 85.68 0.28 85.68 0.765 84.98 0.765 84.98 0.28 84.76 0.28 84.76 0.765 84.06 0.765 84.06 0.28 83.84 0.28 83.84 0.765 83.14 0.765 83.14 0.28 82.92 0.28 82.92 0.765 82.22 0.765 82.22 0.28 81.54 0.28 81.54 0.765 80.84 0.765 80.84 0.28 80.62 0.28 80.62 0.765 79.92 0.765 79.92 0.28 79.7 0.28 79.7 0.765 79 0.765 79 0.28 78.78 0.28 78.78 0.765 78.08 0.765 78.08 0.28 77.86 0.28 77.86 0.765 77.16 0.765 77.16 0.28 76.94 0.28 76.94 0.765 76.24 0.765 76.24 0.28 76.02 0.28 76.02 0.765 75.32 0.765 75.32 0.28 75.1 0.28 75.1 0.765 74.4 0.765 74.4 0.28 74.18 0.28 74.18 0.765 73.48 0.765 73.48 0.28 73.26 0.28 73.26 0.765 72.56 0.765 72.56 0.28 71.88 0.28 71.88 0.765 71.18 0.765 71.18 0.28 70.96 0.28 70.96 0.765 70.26 0.765 70.26 0.28 70.04 0.28 70.04 0.765 69.34 0.765 69.34 0.28 69.12 0.28 69.12 0.765 68.42 0.765 68.42 0.28 67.74 0.28 67.74 0.765 67.04 0.765 67.04 0.28 66.82 0.28 66.82 0.765 66.12 0.765 66.12 0.28 65.9 0.28 65.9 0.765 65.2 0.765 65.2 0.28 64.98 0.28 64.98 0.765 64.28 0.765 64.28 0.28 64.06 0.28 64.06 0.765 63.36 0.765 63.36 0.28 63.14 0.28 63.14 0.765 62.44 0.765 62.44 0.28 62.22 0.28 62.22 0.765 61.52 0.765 61.52 0.28 61.3 0.28 61.3 0.765 60.6 0.765 60.6 0.28 59.46 0.28 59.46 0.765 58.76 0.765 58.76 0.28 49.34 0.28 49.34 0.765 48.64 0.765 48.64 0.28 48.42 0.28 48.42 0.765 47.72 0.765 47.72 0.28 47.5 0.28 47.5 0.765 46.8 0.765 46.8 0.28 46.58 0.28 46.58 0.765 45.88 0.765 45.88 0.28 45.66 0.28 45.66 0.765 44.96 0.765 44.96 0.28 44.74 0.28 44.74 0.765 44.04 0.765 44.04 0.28 43.82 0.28 43.82 0.765 43.12 0.765 43.12 0.28 42.9 0.28 42.9 0.765 42.2 0.765 42.2 0.28 41.98 0.28 41.98 0.765 41.28 0.765 41.28 0.28 41.06 0.28 41.06 0.765 40.36 0.765 40.36 0.28 40.14 0.28 40.14 0.765 39.44 0.765 39.44 0.28 30.64 0.28 30.64 5.72 18.98 5.72 18.98 6.205 18.28 6.205 18.28 5.72 18.06 5.72 18.06 6.205 17.36 6.205 17.36 5.72 17.14 5.72 17.14 6.205 16.44 6.205 16.44 5.72 15.76 5.72 15.76 6.205 15.06 6.205 15.06 5.72 14.84 5.72 14.84 6.205 14.14 6.205 14.14 5.72 13.92 5.72 13.92 6.205 13.22 6.205 13.22 5.72 12.54 5.72 12.54 6.205 11.84 6.205 11.84 5.72 11.62 5.72 11.62 6.205 10.92 6.205 10.92 5.72 10.7 5.72 10.7 6.205 10 6.205 10 5.72 9.78 5.72 9.78 6.205 9.08 6.205 9.08 5.72 8.86 5.72 8.86 6.205 8.16 6.205 8.16 5.72 7.94 5.72 7.94 6.205 7.24 6.205 7.24 5.72 4.26 5.72 4.26 6.205 3.56 6.205 3.56 5.72 3.34 5.72 3.34 6.205 2.64 6.205 2.64 5.72 0.28 5.72 0.28 124.84 3.56 124.84 3.56 124.355 4.26 124.355 4.26 124.84 10.92 124.84 10.92 124.355 11.62 124.355 11.62 124.84 11.84 124.84 11.84 124.355 12.54 124.355 12.54 124.84 14.14 124.84 14.14 124.355 14.84 124.355 14.84 124.84 16.9 124.84 16.9 124.355 17.6 124.355 17.6 124.84 17.82 124.84 17.82 124.355 18.52 124.355 18.52 124.84 18.74 124.84 18.74 124.355 19.44 124.355 19.44 124.84 20.12 124.84 20.12 124.355 20.82 124.355 20.82 124.84 30.64 124.84 30.64 130.28 34.38 130.28 34.38 129.795 35.08 129.795 35.08 130.28 35.3 130.28 35.3 129.795 36 129.795 36 130.28 36.22 130.28 36.22 129.795 36.92 129.795 36.92 130.28 37.14 130.28 37.14 129.795 37.84 129.795 37.84 130.28 38.52 130.28 38.52 129.795 39.22 129.795 39.22 130.28 39.44 130.28 39.44 129.795 40.14 129.795 40.14 130.28 40.82 130.28 40.82 129.795 41.52 129.795 41.52 130.28 41.74 130.28 41.74 129.795 42.44 129.795 42.44 130.28 43.12 130.28 43.12 129.795 43.82 129.795 43.82 130.28 44.04 130.28 44.04 129.795 44.74 129.795 44.74 130.28 44.96 130.28 44.96 129.795 45.66 129.795 45.66 130.28 45.88 130.28 45.88 129.795 46.58 129.795 46.58 130.28 46.8 130.28 46.8 129.795 47.5 129.795 47.5 130.28 47.72 130.28 47.72 129.795 48.42 129.795 48.42 130.28 48.64 130.28 48.64 129.795 49.34 129.795 49.34 130.28 49.56 130.28 49.56 129.795 50.26 129.795 50.26 130.28 58.76 130.28 58.76 129.795 59.46 129.795 59.46 130.28 60.6 130.28 60.6 129.795 61.3 129.795 61.3 130.28 61.52 130.28 61.52 129.795 62.22 129.795 62.22 130.28 62.44 130.28 62.44 129.795 63.14 129.795 63.14 130.28 63.36 130.28 63.36 129.795 64.06 129.795 64.06 130.28 64.28 130.28 64.28 129.795 64.98 129.795 64.98 130.28 65.2 130.28 65.2 129.795 65.9 129.795 65.9 130.28 66.12 130.28 66.12 129.795 66.82 129.795 66.82 130.28 67.04 130.28 67.04 129.795 67.74 129.795 67.74 130.28 67.96 130.28 67.96 129.795 68.66 129.795 68.66 130.28 68.88 130.28 68.88 129.795 69.58 129.795 69.58 130.28 69.8 130.28 69.8 129.795 70.5 129.795 70.5 130.28 70.72 130.28 70.72 129.795 71.42 129.795 71.42 130.28 71.64 130.28 71.64 129.795 72.34 129.795 72.34 130.28 72.56 130.28 72.56 129.795 73.26 129.795 73.26 130.28 73.48 130.28 73.48 129.795 74.18 129.795 74.18 130.28 74.4 130.28 74.4 129.795 75.1 129.795 75.1 130.28 75.32 130.28 75.32 129.795 76.02 129.795 76.02 130.28 76.24 130.28 76.24 129.795 76.94 129.795 76.94 130.28 77.16 130.28 77.16 129.795 77.86 129.795 77.86 130.28 78.08 130.28 78.08 129.795 78.78 129.795 78.78 130.28 79 130.28 79 129.795 79.7 129.795 79.7 130.28 79.92 130.28 79.92 129.795 80.62 129.795 80.62 130.28 81.3 130.28 81.3 129.795 82 129.795 82 130.28 82.22 130.28 82.22 129.795 82.92 129.795 82.92 130.28 83.14 130.28 83.14 129.795 83.84 129.795 83.84 130.28 84.06 130.28 84.06 129.795 84.76 129.795 84.76 130.28 84.98 130.28 84.98 129.795 85.68 129.795 85.68 130.28 85.9 130.28 85.9 129.795 86.6 129.795 86.6 130.28 86.82 130.28 86.82 129.795 87.52 129.795 87.52 130.28 87.74 130.28 87.74 129.795 88.44 129.795 88.44 130.28 89.58 130.28 89.58 129.795 90.28 129.795 90.28 130.28 90.5 130.28 90.5 129.795 91.2 129.795 91.2 130.28 91.42 130.28 91.42 129.795 92.12 129.795 92.12 130.28 92.34 130.28 92.34 129.795 93.04 129.795 93.04 130.28 93.72 130.28 93.72 129.795 94.42 129.795 94.42 130.28 94.64 130.28 94.64 129.795 95.34 129.795 95.34 130.28 95.56 130.28 95.56 129.795 96.26 129.795 96.26 130.28 96.94 130.28 96.94 129.795 97.64 129.795 97.64 130.28 97.86 130.28 97.86 129.795 98.56 129.795 98.56 130.28 98.78 130.28 98.78 129.795 99.48 129.795 99.48 130.28 99.7 130.28 99.7 129.795 100.4 129.795 100.4 130.28 101.08 130.28 101.08 129.795 101.78 129.795 101.78 130.28 ;
    LAYER met4 ;
      POLYGON 102.745 130.385 102.745 130.055 102.73 130.055 102.73 112.39 102.43 112.39 102.43 130.055 102.415 130.055 102.415 130.385 ;
      POLYGON 71.465 130.385 71.465 130.055 71.45 130.055 71.45 128.03 71.15 128.03 71.15 130.055 71.135 130.055 71.135 130.385 ;
      POLYGON 69.61 130.37 69.61 121.91 69.31 121.91 69.31 130.07 69.09 130.07 69.09 130.37 ;
      POLYGON 66.85 130.37 66.85 119.19 66.55 119.19 66.55 130.07 66.33 130.07 66.33 130.37 ;
      POLYGON 53.05 95.01 53.05 0.505 53.065 0.505 53.065 0.175 52.735 0.175 52.735 0.505 52.75 0.505 52.75 95.01 ;
      POLYGON 103.65 16.81 103.65 5.945 103.665 5.945 103.665 5.615 103.335 5.615 103.335 5.945 103.35 5.945 103.35 16.81 ;
      POLYGON 12.57 14.09 12.57 5.945 12.585 5.945 12.585 5.615 12.255 5.615 12.255 5.945 12.27 5.945 12.27 14.09 ;
      POLYGON 103.56 130.16 103.56 124.72 119.82 124.72 119.82 124.12 121.22 124.12 121.22 124.72 133.92 124.72 133.92 5.84 121.22 5.84 121.22 6.44 119.82 6.44 119.82 5.84 103.56 5.84 103.56 0.4 98.53 0.4 98.53 1.2 97.43 1.2 97.43 0.4 96.69 0.4 96.69 1.2 95.59 1.2 95.59 0.4 94.85 0.4 94.85 1.2 93.75 1.2 93.75 0.4 93.01 0.4 93.01 1.2 91.91 1.2 91.91 0.4 91.17 0.4 91.17 1.2 90.07 1.2 90.07 0.4 89.94 0.4 89.94 1 88.54 1 88.54 0.4 87.49 0.4 87.49 1.2 86.39 1.2 86.39 0.4 85.65 0.4 85.65 1.2 84.55 1.2 84.55 0.4 83.81 0.4 83.81 1.2 82.71 1.2 82.71 0.4 81.97 0.4 81.97 1.2 80.87 1.2 80.87 0.4 80.13 0.4 80.13 1.2 79.03 1.2 79.03 0.4 78.29 0.4 78.29 1.2 77.19 1.2 77.19 0.4 76.45 0.4 76.45 1.2 75.35 1.2 75.35 0.4 75.22 0.4 75.22 1 73.82 1 73.82 0.4 72.77 0.4 72.77 1.2 71.67 1.2 71.67 0.4 70.93 0.4 70.93 1.2 69.83 1.2 69.83 0.4 69.09 0.4 69.09 1.2 67.99 1.2 67.99 0.4 67.25 0.4 67.25 1.2 66.15 1.2 66.15 0.4 65.41 0.4 65.41 1.2 64.31 1.2 64.31 0.4 63.57 0.4 63.57 1.2 62.47 1.2 62.47 0.4 61.73 0.4 61.73 1.2 60.63 1.2 60.63 0.4 60.5 0.4 60.5 1 59.1 1 59.1 0.4 45.78 0.4 45.78 1 44.38 1 44.38 0.4 30.76 0.4 30.76 5.84 14.5 5.84 14.5 6.44 13.1 6.44 13.1 5.84 0.4 5.84 0.4 124.72 13.1 124.72 13.1 124.12 14.5 124.12 14.5 124.72 30.76 124.72 30.76 130.16 44.38 130.16 44.38 129.56 45.78 129.56 45.78 130.16 59.1 130.16 59.1 129.56 60.5 129.56 60.5 130.16 61.55 130.16 61.55 129.36 62.65 129.36 62.65 130.16 63.39 130.16 63.39 129.36 64.49 129.36 64.49 130.16 65.23 130.16 65.23 129.36 66.33 129.36 66.33 130.16 67.99 130.16 67.99 129.36 69.09 129.36 69.09 130.16 69.83 130.16 69.83 129.36 70.93 129.36 70.93 130.16 71.67 130.16 71.67 129.36 72.77 129.36 72.77 130.16 73.82 130.16 73.82 129.56 75.22 129.56 75.22 130.16 75.35 130.16 75.35 129.36 76.45 129.36 76.45 130.16 77.19 130.16 77.19 129.36 78.29 129.36 78.29 130.16 79.03 130.16 79.03 129.36 80.13 129.36 80.13 130.16 80.87 130.16 80.87 129.36 81.97 129.36 81.97 130.16 82.71 130.16 82.71 129.36 83.81 129.36 83.81 130.16 84.55 130.16 84.55 129.36 85.65 129.36 85.65 130.16 86.39 130.16 86.39 129.36 87.49 129.36 87.49 130.16 88.54 130.16 88.54 129.56 89.94 129.56 89.94 130.16 90.07 130.16 90.07 129.36 91.17 129.36 91.17 130.16 91.91 130.16 91.91 129.36 93.01 129.36 93.01 130.16 98.35 130.16 98.35 129.36 99.45 129.36 99.45 130.16 ;
    LAYER met3 ;
      POLYGON 89.405 130.605 89.405 130.6 89.62 130.6 89.62 130.28 89.405 130.28 89.405 130.275 89.075 130.275 89.075 130.28 88.86 130.28 88.86 130.6 89.075 130.6 89.075 130.605 ;
      POLYGON 59.965 130.605 59.965 130.6 60.18 130.6 60.18 130.28 59.965 130.28 59.965 130.275 59.635 130.275 59.635 130.28 59.42 130.28 59.42 130.6 59.635 130.6 59.635 130.605 ;
      POLYGON 101.595 130.385 101.595 130.37 102.39 130.37 102.39 130.38 102.77 130.38 102.77 130.06 102.39 130.06 102.39 130.07 101.595 130.07 101.595 130.055 101.265 130.055 101.265 130.07 91.015 130.07 91.015 130.055 90.685 130.055 90.685 130.385 91.015 130.385 91.015 130.37 101.265 130.37 101.265 130.385 ;
      POLYGON 84.115 130.385 84.115 130.055 83.785 130.055 83.785 130.07 83.45 130.07 83.45 130.06 83.07 130.06 83.07 130.38 83.45 130.38 83.45 130.37 83.785 130.37 83.785 130.385 ;
      POLYGON 70.775 130.385 70.775 130.055 70.445 130.055 70.445 130.06 70.035 130.06 70.035 130.38 70.445 130.38 70.445 130.385 ;
      POLYGON 76.09 130.38 76.09 130.06 75.71 130.06 75.71 130.07 71.49 130.07 71.49 130.06 71.11 130.06 71.11 130.38 71.49 130.38 71.49 130.37 75.71 130.37 75.71 130.38 ;
      POLYGON 123.66 124.93 123.66 123.95 123.36 123.95 123.36 124.63 101.74 124.63 101.74 124.93 ;
      POLYGON 20.16 124.93 20.16 123.95 19.86 123.95 19.86 124.63 17.86 124.63 17.86 123.95 17.56 123.95 17.56 124.93 ;
      RECT 1.19 58.66 1.57 58.98 ;
      RECT 1.19 47.78 1.57 48.1 ;
      POLYGON 133.335 26.345 133.335 26.015 133.005 26.015 133.005 26.03 125.43 26.03 125.43 26.33 133.005 26.33 133.005 26.345 ;
      RECT 1.035 13.1 1.57 13.42 ;
      POLYGON 120.915 5.945 120.915 5.615 120.585 5.615 120.585 5.63 109.415 5.63 109.415 5.615 109.085 5.615 109.085 5.945 109.415 5.945 109.415 5.93 120.585 5.93 120.585 5.945 ;
      POLYGON 12.355 5.945 12.355 5.94 12.61 5.94 12.61 5.62 12.355 5.62 12.355 5.615 12.025 5.615 12.025 5.62 11.655 5.62 11.655 5.94 12.025 5.94 12.025 5.945 ;
      POLYGON 103.69 5.94 103.69 5.62 103.31 5.62 103.31 5.63 102.66 5.63 102.66 5.93 103.31 5.93 103.31 5.94 ;
      POLYGON 76.05 1.85 76.05 0.5 76.09 0.5 76.09 0.18 75.71 0.18 75.71 0.5 75.75 0.5 75.75 1.85 ;
      POLYGON 72.385 0.675 72.385 0.67 72.41 0.67 72.41 0.35 72.385 0.35 72.385 0.345 71.655 0.345 71.655 0.675 ;
      POLYGON 96.075 0.505 96.075 0.175 95.745 0.175 95.745 0.19 94.49 0.19 94.49 0.18 94.11 0.18 94.11 0.5 94.49 0.5 94.49 0.49 95.745 0.49 95.745 0.505 ;
      POLYGON 86.875 0.505 86.875 0.175 86.545 0.175 86.545 0.19 85.29 0.19 85.29 0.18 84.91 0.18 84.91 0.5 85.29 0.5 85.29 0.49 86.545 0.49 86.545 0.505 ;
      POLYGON 64.335 0.505 64.335 0.49 68.35 0.49 68.35 0.5 68.73 0.5 68.73 0.18 68.35 0.18 68.35 0.19 64.335 0.19 64.335 0.175 64.005 0.175 64.005 0.505 ;
      POLYGON 49.155 0.505 49.155 0.49 52.71 0.49 52.71 0.5 53.09 0.5 53.09 0.18 52.71 0.18 52.71 0.19 49.155 0.19 49.155 0.175 48.825 0.175 48.825 0.505 ;
      POLYGON 89.405 0.285 89.405 0.28 89.62 0.28 89.62 -0.04 89.405 -0.04 89.405 -0.045 89.075 -0.045 89.075 -0.04 88.86 -0.04 88.86 0.28 89.075 0.28 89.075 0.285 ;
      POLYGON 59.965 0.285 59.965 0.28 60.18 0.28 60.18 -0.04 59.965 -0.04 59.965 -0.045 59.635 -0.045 59.635 -0.04 59.42 -0.04 59.42 0.28 59.635 0.28 59.635 0.285 ;
      POLYGON 103.56 130.16 103.56 124.72 133.92 124.72 133.92 68.21 133.12 68.21 133.12 67.11 133.92 67.11 133.92 66.85 133.12 66.85 133.12 65.75 133.92 65.75 133.92 65.49 133.12 65.49 133.12 64.39 133.92 64.39 133.92 64.13 133.12 64.13 133.12 63.03 133.92 63.03 133.92 62.77 133.12 62.77 133.12 61.67 133.92 61.67 133.92 61.41 133.12 61.41 133.12 60.31 133.92 60.31 133.92 60.05 133.12 60.05 133.12 58.95 133.92 58.95 133.92 47.81 133.12 47.81 133.12 46.71 133.92 46.71 133.92 46.45 133.12 46.45 133.12 45.35 133.92 45.35 133.92 45.09 133.12 45.09 133.12 43.99 133.92 43.99 133.92 27.41 133.12 27.41 133.12 26.31 133.92 26.31 133.92 26.05 133.12 26.05 133.12 24.95 133.92 24.95 133.92 24.69 133.12 24.69 133.12 23.59 133.92 23.59 133.92 23.33 133.12 23.33 133.12 22.23 133.92 22.23 133.92 21.97 133.12 21.97 133.12 20.87 133.92 20.87 133.92 14.49 133.12 14.49 133.12 13.39 133.92 13.39 133.92 13.13 133.12 13.13 133.12 12.03 133.92 12.03 133.92 11.77 133.12 11.77 133.12 10.67 133.92 10.67 133.92 5.84 103.56 5.84 103.56 0.4 30.76 0.4 30.76 5.84 0.4 5.84 0.4 10.67 1.2 10.67 1.2 11.77 0.4 11.77 0.4 12.03 1.2 12.03 1.2 13.13 0.4 13.13 0.4 13.39 1.2 13.39 1.2 14.49 0.4 14.49 0.4 23.59 1.2 23.59 1.2 24.69 0.4 24.69 0.4 42.63 1.2 42.63 1.2 43.73 0.4 43.73 0.4 43.99 1.2 43.99 1.2 45.09 0.4 45.09 0.4 45.35 1.2 45.35 1.2 46.45 0.4 46.45 0.4 46.71 1.2 46.71 1.2 47.81 0.4 47.81 0.4 48.07 1.2 48.07 1.2 49.17 0.4 49.17 0.4 49.43 1.2 49.43 1.2 50.53 0.4 50.53 0.4 53.51 1.2 53.51 1.2 54.61 0.4 54.61 0.4 54.87 1.2 54.87 1.2 55.97 0.4 55.97 0.4 56.23 1.2 56.23 1.2 57.33 0.4 57.33 0.4 57.59 1.2 57.59 1.2 58.69 0.4 58.69 0.4 58.95 1.2 58.95 1.2 60.05 0.4 60.05 0.4 60.31 1.2 60.31 1.2 61.41 0.4 61.41 0.4 61.67 1.2 61.67 1.2 62.77 0.4 62.77 0.4 63.03 1.2 63.03 1.2 64.13 0.4 64.13 0.4 64.39 1.2 64.39 1.2 65.49 0.4 65.49 0.4 65.75 1.2 65.75 1.2 66.85 0.4 66.85 0.4 67.11 1.2 67.11 1.2 68.21 0.4 68.21 0.4 124.72 30.76 124.72 30.76 130.16 ;
    LAYER met1 ;
      POLYGON 103.2 130.8 103.2 130.32 89.4 130.32 89.4 130.31 89.08 130.31 89.08 130.32 59.96 130.32 59.96 130.31 59.64 130.31 59.64 130.32 31.12 130.32 31.12 130.8 ;
      RECT 53.96 124.88 133.56 125.36 ;
      RECT 0.76 124.88 52.76 125.36 ;
      POLYGON 133.795 66.88 133.795 66.82 133.445 66.82 133.445 66.74 130.34 66.74 130.34 66.88 ;
      POLYGON 133.795 62.12 133.795 62.06 133.445 62.06 133.445 61.98 123.44 61.98 123.44 62.12 ;
      RECT 53.96 5.2 133.56 5.68 ;
      RECT 0.76 5.2 52.76 5.68 ;
      POLYGON 89.4 0.25 89.4 0.24 103.2 0.24 103.2 -0.24 31.12 -0.24 31.12 0.24 59.64 0.24 59.64 0.25 59.96 0.25 59.96 0.24 89.08 0.24 89.08 0.25 ;
      POLYGON 103.2 130.28 103.2 130.04 103.68 130.04 103.68 128.36 103.2 128.36 103.2 127.32 103.68 127.32 103.68 124.84 133.56 124.84 133.56 124.6 134.04 124.6 134.04 122.92 133.56 122.92 133.56 121.88 134.04 121.88 134.04 120.2 133.56 120.2 133.56 119.16 134.04 119.16 134.04 118.16 133.445 118.16 133.445 117.46 133.56 117.46 133.56 116.44 134.04 116.44 134.04 116.12 133.445 116.12 133.445 115.42 134.04 115.42 134.04 114.76 133.56 114.76 133.56 113.74 133.445 113.74 133.445 113.04 134.04 113.04 134.04 112.72 133.445 112.72 133.445 112.02 133.56 112.02 133.56 111.02 133.445 111.02 133.445 109.64 134.04 109.64 134.04 109.32 133.56 109.32 133.56 108.3 133.445 108.3 133.445 106.92 134.04 106.92 134.04 106.6 133.56 106.6 133.56 105.56 134.04 105.56 134.04 103.88 133.56 103.88 133.56 102.84 134.04 102.84 134.04 102.52 133.445 102.52 133.445 101.14 133.56 101.14 133.56 100.12 134.04 100.12 134.04 98.44 133.56 98.44 133.56 97.4 134.04 97.4 134.04 95.72 133.56 95.72 133.56 94.68 134.04 94.68 134.04 93 133.56 93 133.56 91.96 134.04 91.96 134.04 90.28 133.56 90.28 133.56 89.26 133.445 89.26 133.445 88.56 134.04 88.56 134.04 87.56 133.56 87.56 133.56 86.52 134.04 86.52 134.04 84.84 133.56 84.84 133.56 83.8 134.04 83.8 134.04 82.12 133.56 82.12 133.56 81.08 134.04 81.08 134.04 80.76 133.445 80.76 133.445 79.38 133.56 79.38 133.56 78.36 134.04 78.36 134.04 76.68 133.56 76.68 133.56 75.64 134.04 75.64 134.04 73.96 133.56 73.96 133.56 72.92 134.04 72.92 134.04 71.24 133.56 71.24 133.56 70.2 134.04 70.2 134.04 68.52 133.56 68.52 133.56 67.5 133.445 67.5 133.445 66.12 134.04 66.12 134.04 65.8 133.56 65.8 133.56 64.78 133.445 64.78 133.445 63.4 134.04 63.4 134.04 63.08 133.56 63.08 133.56 62.06 133.445 62.06 133.445 60.68 134.04 60.68 134.04 60.36 133.56 60.36 133.56 59.34 133.445 59.34 133.445 57.96 134.04 57.96 134.04 57.64 133.56 57.64 133.56 56.62 133.445 56.62 133.445 55.24 134.04 55.24 134.04 54.92 133.56 54.92 133.56 53.9 133.445 53.9 133.445 53.2 134.04 53.2 134.04 52.88 133.445 52.88 133.445 52.18 133.56 52.18 133.56 51.16 134.04 51.16 134.04 50.84 133.445 50.84 133.445 49.46 133.56 49.46 133.56 48.44 134.04 48.44 134.04 48.12 133.445 48.12 133.445 46.74 133.56 46.74 133.56 45.74 133.445 45.74 133.445 44.36 134.04 44.36 134.04 44.04 133.56 44.04 133.56 43.02 133.445 43.02 133.445 41.64 134.04 41.64 134.04 41.32 133.56 41.32 133.56 40.3 133.445 40.3 133.445 38.92 134.04 38.92 134.04 38.6 133.56 38.6 133.56 37.58 133.445 37.58 133.445 36.2 134.04 36.2 134.04 35.88 133.56 35.88 133.56 34.84 134.04 34.84 134.04 34.52 133.445 34.52 133.445 33.14 133.56 33.14 133.56 32.12 134.04 32.12 134.04 31.8 133.445 31.8 133.445 30.42 133.56 30.42 133.56 29.4 134.04 29.4 134.04 29.08 133.445 29.08 133.445 27.7 133.56 27.7 133.56 26.68 134.04 26.68 134.04 26.36 133.445 26.36 133.445 24.98 133.56 24.98 133.56 23.98 133.445 23.98 133.445 22.6 134.04 22.6 134.04 22.28 133.56 22.28 133.56 21.26 133.445 21.26 133.445 19.88 134.04 19.88 134.04 19.56 133.56 19.56 133.56 18.54 133.445 18.54 133.445 17.16 134.04 17.16 134.04 16.84 133.56 16.84 133.56 15.82 133.445 15.82 133.445 14.44 134.04 14.44 134.04 14.12 133.56 14.12 133.56 13.08 134.04 13.08 134.04 12.76 133.445 12.76 133.445 11.38 133.56 11.38 133.56 10.36 134.04 10.36 134.04 8.68 133.56 8.68 133.56 7.64 134.04 7.64 134.04 5.96 133.56 5.96 133.56 5.72 103.68 5.72 103.68 3.24 103.2 3.24 103.2 2.2 103.68 2.2 103.68 0.52 103.2 0.52 103.2 0.28 31.12 0.28 31.12 0.52 30.64 0.52 30.64 2.2 31.12 2.2 31.12 3.24 30.64 3.24 30.64 5.72 0.76 5.72 0.76 5.96 0.28 5.96 0.28 6.96 0.875 6.96 0.875 7.66 0.76 7.66 0.76 8.66 0.875 8.66 0.875 9.36 0.28 9.36 0.28 10.36 0.76 10.36 0.76 11.38 0.875 11.38 0.875 12.08 0.28 12.08 0.28 12.4 0.875 12.4 0.875 13.1 0.76 13.1 0.76 14.12 0.28 14.12 0.28 14.44 0.875 14.44 0.875 15.82 0.76 15.82 0.76 16.84 0.28 16.84 0.28 17.16 0.875 17.16 0.875 18.54 0.76 18.54 0.76 19.56 0.28 19.56 0.28 19.88 0.875 19.88 0.875 21.26 0.76 21.26 0.76 22.28 0.28 22.28 0.28 22.6 0.875 22.6 0.875 23.98 0.76 23.98 0.76 24.98 0.875 24.98 0.875 26.36 0.28 26.36 0.28 26.68 0.76 26.68 0.76 27.7 0.875 27.7 0.875 29.08 0.28 29.08 0.28 29.4 0.76 29.4 0.76 30.42 0.875 30.42 0.875 31.8 0.28 31.8 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 33.48 0.875 33.48 0.875 34.86 0.76 34.86 0.76 35.86 0.875 35.86 0.875 36.56 0.28 36.56 0.28 36.88 0.875 36.88 0.875 37.58 0.76 37.58 0.76 38.6 0.28 38.6 0.28 38.92 0.875 38.92 0.875 40.3 0.76 40.3 0.76 41.32 0.28 41.32 0.28 41.64 0.875 41.64 0.875 43.02 0.76 43.02 0.76 44.04 0.28 44.04 0.28 44.36 0.875 44.36 0.875 45.74 0.76 45.74 0.76 46.74 0.875 46.74 0.875 48.12 0.28 48.12 0.28 48.44 0.76 48.44 0.76 49.46 0.875 49.46 0.875 50.84 0.28 50.84 0.28 51.16 0.76 51.16 0.76 52.18 0.875 52.18 0.875 53.56 0.28 53.56 0.28 53.88 0.76 53.88 0.76 54.9 0.875 54.9 0.875 56.28 0.28 56.28 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 57.96 0.875 57.96 0.875 59.34 0.76 59.34 0.76 60.36 0.28 60.36 0.28 60.68 0.875 60.68 0.875 62.06 0.76 62.06 0.76 63.08 0.28 63.08 0.28 63.4 0.875 63.4 0.875 64.78 0.76 64.78 0.76 65.8 0.28 65.8 0.28 66.12 0.875 66.12 0.875 67.5 0.76 67.5 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.38 0.875 79.38 0.875 80.08 0.28 80.08 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 88.56 0.875 88.56 0.875 89.26 0.76 89.26 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 0.76 97.4 0.76 98.44 0.28 98.44 0.28 100.12 0.76 100.12 0.76 101.16 0.28 101.16 0.28 102.84 0.76 102.84 0.76 103.88 0.28 103.88 0.28 105.56 0.76 105.56 0.76 106.6 0.28 106.6 0.28 108.28 0.76 108.28 0.76 109.32 0.28 109.32 0.28 109.64 0.875 109.64 0.875 111.02 0.76 111.02 0.76 112.02 0.875 112.02 0.875 113.4 0.28 113.4 0.28 113.72 0.76 113.72 0.76 114.74 0.875 114.74 0.875 115.44 0.28 115.44 0.28 116.44 0.76 116.44 0.76 117.48 0.28 117.48 0.28 118.14 0.875 118.14 0.875 118.84 0.28 118.84 0.28 119.16 0.76 119.16 0.76 120.18 0.875 120.18 0.875 120.88 0.28 120.88 0.28 121.2 0.875 121.2 0.875 121.9 0.76 121.9 0.76 122.92 0.28 122.92 0.28 124.6 0.76 124.6 0.76 124.84 30.64 124.84 30.64 127.32 31.12 127.32 31.12 128.36 30.64 128.36 30.64 130.04 31.12 130.04 31.12 130.28 ;
    LAYER met5 ;
      POLYGON 102.36 128.96 102.36 123.52 132.72 123.52 132.72 109.28 129.52 109.28 129.52 102.88 132.72 102.88 132.72 88.88 129.52 88.88 129.52 82.48 132.72 82.48 132.72 68.48 129.52 68.48 129.52 62.08 132.72 62.08 132.72 48.08 129.52 48.08 129.52 41.68 132.72 41.68 132.72 27.68 129.52 27.68 129.52 21.28 132.72 21.28 132.72 7.04 102.36 7.04 102.36 1.6 31.96 1.6 31.96 7.04 1.6 7.04 1.6 21.28 4.8 21.28 4.8 27.68 1.6 27.68 1.6 41.68 4.8 41.68 4.8 48.08 1.6 48.08 1.6 62.08 4.8 62.08 4.8 68.48 1.6 68.48 1.6 82.48 4.8 82.48 4.8 88.88 1.6 88.88 1.6 102.88 4.8 102.88 4.8 109.28 1.6 109.28 1.6 123.52 31.96 123.52 31.96 128.96 ;
    LAYER li1 ;
      POLYGON 103.96 130.645 103.96 130.475 100.725 130.475 100.725 129.675 100.395 129.675 100.395 130.475 99.885 130.475 99.885 129.995 99.555 129.995 99.555 130.475 99.045 130.475 99.045 129.995 98.715 129.995 98.715 130.475 98.205 130.475 98.205 129.995 97.875 129.995 97.875 130.475 97.365 130.475 97.365 129.995 97.035 129.995 97.035 130.475 96.525 130.475 96.525 129.995 96.195 129.995 96.195 130.475 95.165 130.475 95.165 129.995 94.835 129.995 94.835 130.475 94.325 130.475 94.325 129.995 93.995 129.995 93.995 130.475 93.485 130.475 93.485 129.995 93.155 129.995 93.155 130.475 92.645 130.475 92.645 129.995 92.315 129.995 92.315 130.475 91.805 130.475 91.805 129.995 91.475 129.995 91.475 130.475 90.965 130.475 90.965 129.675 90.635 129.675 90.635 130.475 89.685 130.475 89.685 129.675 89.355 129.675 89.355 130.475 88.845 130.475 88.845 129.995 88.515 129.995 88.515 130.475 88.005 130.475 88.005 129.995 87.675 129.995 87.675 130.475 87.165 130.475 87.165 129.995 86.835 129.995 86.835 130.475 86.325 130.475 86.325 129.995 85.995 129.995 85.995 130.475 85.485 130.475 85.485 129.995 85.155 129.995 85.155 130.475 84.165 130.475 84.165 129.675 83.835 129.675 83.835 130.475 83.325 130.475 83.325 129.995 82.995 129.995 82.995 130.475 82.485 130.475 82.485 129.995 82.155 129.995 82.155 130.475 81.645 130.475 81.645 129.995 81.315 129.995 81.315 130.475 80.805 130.475 80.805 129.995 80.475 129.995 80.475 130.475 79.965 130.475 79.965 129.995 79.635 129.995 79.635 130.475 78.605 130.475 78.605 129.995 78.275 129.995 78.275 130.475 77.765 130.475 77.765 129.995 77.435 129.995 77.435 130.475 76.925 130.475 76.925 129.995 76.595 129.995 76.595 130.475 76.085 130.475 76.085 129.995 75.755 129.995 75.755 130.475 75.245 130.475 75.245 129.995 74.915 129.995 74.915 130.475 74.405 130.475 74.405 129.675 74.075 129.675 74.075 130.475 71.625 130.475 71.625 130.015 71.32 130.015 71.32 130.475 70.65 130.475 70.65 130.015 70.48 130.015 70.48 130.475 69.81 130.475 69.81 130.015 69.64 130.015 69.64 130.475 68.97 130.475 68.97 130.015 68.8 130.015 68.8 130.475 68.13 130.475 68.13 130.015 67.875 130.015 67.875 130.475 67.485 130.475 67.485 130.015 67.18 130.015 67.18 130.475 66.51 130.475 66.51 130.015 66.34 130.015 66.34 130.475 65.67 130.475 65.67 130.015 65.5 130.015 65.5 130.475 64.83 130.475 64.83 130.015 64.66 130.015 64.66 130.475 63.99 130.475 63.99 130.015 63.735 130.015 63.735 130.475 63.225 130.475 63.225 130.015 62.97 130.015 62.97 130.475 62.3 130.475 62.3 130.015 62.13 130.015 62.13 130.475 61.46 130.475 61.46 130.015 61.29 130.015 61.29 130.475 60.62 130.475 60.62 130.015 60.45 130.015 60.45 130.475 59.78 130.475 59.78 130.015 59.475 130.015 59.475 130.475 59.125 130.475 59.125 129.74 58.785 129.74 58.785 130.475 54.365 130.475 54.365 129.74 54.035 129.74 54.035 130.475 53.565 130.475 53.565 130.015 53.31 130.015 53.31 130.475 52.64 130.475 52.64 130.015 52.47 130.015 52.47 130.475 51.8 130.475 51.8 130.015 51.63 130.015 51.63 130.475 50.96 130.475 50.96 130.015 50.79 130.015 50.79 130.475 50.12 130.475 50.12 130.015 49.815 130.015 49.815 130.475 49.585 130.475 49.585 129.675 49.255 129.675 49.255 130.475 48.745 130.475 48.745 129.995 48.415 129.995 48.415 130.475 47.905 130.475 47.905 129.995 47.575 129.995 47.575 130.475 46.985 130.475 46.985 129.995 46.815 129.995 46.815 130.475 46.145 130.475 46.145 129.995 45.975 129.995 45.975 130.475 45.285 130.475 45.285 130.015 45.03 130.015 45.03 130.475 44.36 130.475 44.36 130.015 44.19 130.015 44.19 130.475 43.52 130.475 43.52 130.015 43.35 130.015 43.35 130.475 42.68 130.475 42.68 130.015 42.51 130.015 42.51 130.475 41.84 130.475 41.84 130.015 41.535 130.015 41.535 130.475 41.145 130.475 41.145 130.015 40.89 130.015 40.89 130.475 40.22 130.475 40.22 130.015 40.05 130.015 40.05 130.475 39.38 130.475 39.38 130.015 39.21 130.015 39.21 130.475 38.54 130.475 38.54 130.015 38.37 130.015 38.37 130.475 37.7 130.475 37.7 130.015 37.395 130.015 37.395 130.475 37.005 130.475 37.005 130.015 36.75 130.015 36.75 130.475 36.08 130.475 36.08 130.015 35.91 130.015 35.91 130.475 35.24 130.475 35.24 130.015 35.07 130.015 35.07 130.475 34.4 130.475 34.4 130.015 34.23 130.015 34.23 130.475 33.56 130.475 33.56 130.015 33.255 130.015 33.255 130.475 30.36 130.475 30.36 130.645 ;
      RECT 103.04 127.755 103.96 127.925 ;
      RECT 30.36 127.755 32.2 127.925 ;
      POLYGON 134.32 125.205 134.32 125.035 131.045 125.035 131.045 124.575 130.74 124.575 130.74 125.035 129.255 125.035 129.255 124.595 129.065 124.595 129.065 125.035 127.165 125.035 127.165 124.575 126.835 124.575 126.835 125.035 124.235 125.035 124.235 124.675 123.905 124.675 123.905 125.035 123.205 125.035 123.205 124.655 122.875 124.655 122.875 125.035 121.375 125.035 121.375 124.655 121.045 124.655 121.045 125.035 119.085 125.035 119.085 124.575 118.78 124.575 118.78 125.035 117.295 125.035 117.295 124.595 117.105 124.595 117.105 125.035 115.205 125.035 115.205 124.575 114.875 124.575 114.875 125.035 112.275 125.035 112.275 124.675 111.945 124.675 111.945 125.035 111.245 125.035 111.245 124.655 110.915 124.655 110.915 125.035 110.08 125.035 110.08 124.215 109.85 124.215 109.85 125.035 107.625 125.035 107.625 124.235 107.295 124.235 107.295 125.035 106.785 125.035 106.785 124.555 106.455 124.555 106.455 125.035 105.945 125.035 105.945 124.555 105.615 124.555 105.615 125.035 105.105 125.035 105.105 124.555 104.775 124.555 104.775 125.035 104.265 125.035 104.265 124.555 103.935 124.555 103.935 125.035 103.425 125.035 103.425 124.555 103.095 124.555 103.095 125.035 102.58 125.035 102.58 125.205 ;
      POLYGON 32.2 125.205 32.2 125.035 30.295 125.035 30.295 124.655 29.965 124.655 29.965 125.035 27.69 125.035 27.69 124.215 27.46 124.215 27.46 125.035 26.31 125.035 26.31 124.215 26.08 124.215 26.08 125.035 25.675 125.035 25.675 124.53 25.39 124.53 25.39 125.035 23.55 125.035 23.55 124.215 23.32 124.215 23.32 125.035 22.915 125.035 22.915 124.235 22.605 124.235 22.605 125.035 21.105 125.035 21.105 124.575 20.8 124.575 20.8 125.035 19.315 125.035 19.315 124.595 19.125 124.595 19.125 125.035 17.225 125.035 17.225 124.575 16.895 124.575 16.895 125.035 14.295 125.035 14.295 124.675 13.965 124.675 13.965 125.035 13.265 125.035 13.265 124.655 12.935 124.655 12.935 125.035 11.445 125.035 11.445 124.575 11.14 124.575 11.14 125.035 9.655 125.035 9.655 124.595 9.465 124.595 9.465 125.035 7.565 125.035 7.565 124.575 7.235 124.575 7.235 125.035 4.635 125.035 4.635 124.675 4.305 124.675 4.305 125.035 3.605 125.035 3.605 124.655 3.275 124.655 3.275 125.035 0 125.035 0 125.205 ;
      RECT 133.4 122.315 134.32 122.485 ;
      RECT 0 122.315 1.84 122.485 ;
      RECT 133.4 119.595 134.32 119.765 ;
      RECT 0 119.595 1.84 119.765 ;
      RECT 133.4 116.875 134.32 117.045 ;
      RECT 0 116.875 1.84 117.045 ;
      RECT 133.4 114.155 134.32 114.325 ;
      RECT 0 114.155 1.84 114.325 ;
      RECT 133.4 111.435 134.32 111.605 ;
      RECT 0 111.435 1.84 111.605 ;
      RECT 133.4 108.715 134.32 108.885 ;
      RECT 0 108.715 1.84 108.885 ;
      RECT 133.4 105.995 134.32 106.165 ;
      RECT 0 105.995 1.84 106.165 ;
      RECT 133.4 103.275 134.32 103.445 ;
      RECT 0 103.275 3.68 103.445 ;
      RECT 133.4 100.555 134.32 100.725 ;
      RECT 0 100.555 3.68 100.725 ;
      RECT 133.4 97.835 134.32 98.005 ;
      RECT 0 97.835 1.84 98.005 ;
      RECT 133.4 95.115 134.32 95.285 ;
      RECT 0 95.115 1.84 95.285 ;
      RECT 133.4 92.395 134.32 92.565 ;
      RECT 0 92.395 1.84 92.565 ;
      RECT 133.4 89.675 134.32 89.845 ;
      RECT 0 89.675 1.84 89.845 ;
      RECT 132.48 86.955 134.32 87.125 ;
      RECT 0 86.955 1.84 87.125 ;
      RECT 132.48 84.235 134.32 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 133.4 81.515 134.32 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 133.4 78.795 134.32 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 133.4 76.075 134.32 76.245 ;
      RECT 0 76.075 1.84 76.245 ;
      RECT 133.4 73.355 134.32 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 133.4 70.635 134.32 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 133.86 67.915 134.32 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 133.4 65.195 134.32 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 133.4 62.475 134.32 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 133.4 59.755 134.32 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 133.4 57.035 134.32 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 133.4 54.315 134.32 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 133.4 51.595 134.32 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 133.4 48.875 134.32 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 133.4 46.155 134.32 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 133.4 43.435 134.32 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 133.4 40.715 134.32 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 133.4 37.995 134.32 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 133.4 35.275 134.32 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 133.4 32.555 134.32 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 130.64 29.835 134.32 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 130.64 27.115 134.32 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 133.4 24.395 134.32 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 133.4 21.675 134.32 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 133.4 18.955 134.32 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 133.4 16.235 134.32 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 133.4 13.515 134.32 13.685 ;
      RECT 0 13.515 1.84 13.685 ;
      RECT 133.4 10.795 134.32 10.965 ;
      RECT 0 10.795 1.84 10.965 ;
      RECT 133.4 8.075 134.32 8.245 ;
      RECT 0 8.075 1.84 8.245 ;
      POLYGON 130.73 6.345 130.73 5.525 134.32 5.525 134.32 5.355 101.66 5.355 101.66 5.525 102.175 5.525 102.175 6.005 102.505 6.005 102.505 5.525 103.015 5.525 103.015 6.005 103.345 6.005 103.345 5.525 103.855 5.525 103.855 6.005 104.185 6.005 104.185 5.525 104.695 5.525 104.695 6.005 105.025 6.005 105.025 5.525 105.535 5.525 105.535 6.005 105.865 6.005 105.865 5.525 106.375 5.525 106.375 6.325 106.705 6.325 106.705 5.525 108.155 5.525 108.155 5.905 108.485 5.905 108.485 5.525 109.185 5.525 109.185 5.885 109.515 5.885 109.515 5.525 112.115 5.525 112.115 5.985 112.445 5.985 112.445 5.525 114.345 5.525 114.345 5.965 114.535 5.965 114.535 5.525 116.02 5.525 116.02 5.985 116.325 5.985 116.325 5.525 117.85 5.525 117.85 6.03 118.135 6.03 118.135 5.525 118.435 5.525 118.435 6.26 118.765 6.26 118.765 5.525 126.865 5.525 126.865 6.26 127.205 6.26 127.205 5.525 127.96 5.525 127.96 6.26 128.3 6.26 128.3 5.525 129.81 5.525 129.81 6.03 130.095 6.03 130.095 5.525 130.5 5.525 130.5 6.345 ;
      POLYGON 29.53 6.345 29.53 5.525 30.885 5.525 30.885 5.905 31.215 5.905 31.215 5.525 34.04 5.525 34.04 5.355 0 5.355 0 5.525 3.275 5.525 3.275 5.905 3.605 5.905 3.605 5.525 4.305 5.525 4.305 5.885 4.635 5.885 4.635 5.525 7.235 5.525 7.235 5.985 7.565 5.985 7.565 5.525 9.465 5.525 9.465 5.965 9.655 5.965 9.655 5.525 11.14 5.525 11.14 5.985 11.445 5.985 11.445 5.525 12.475 5.525 12.475 5.905 12.805 5.905 12.805 5.525 13.505 5.525 13.505 5.885 13.835 5.885 13.835 5.525 16.435 5.525 16.435 5.985 16.765 5.985 16.765 5.525 18.665 5.525 18.665 5.965 18.855 5.965 18.855 5.525 20.34 5.525 20.34 5.985 20.645 5.985 20.645 5.525 25.365 5.525 25.365 5.905 25.695 5.905 25.695 5.525 26.54 5.525 26.54 6.345 26.77 6.345 26.77 5.525 27.92 5.525 27.92 6.345 28.15 6.345 28.15 5.525 29.3 5.525 29.3 6.345 ;
      RECT 103.04 2.635 103.96 2.805 ;
      RECT 30.36 2.635 34.04 2.805 ;
      POLYGON 100.725 0.885 100.725 0.085 103.96 0.085 103.96 -0.085 30.36 -0.085 30.36 0.085 33.555 0.085 33.555 0.565 33.725 0.565 33.725 0.085 34.395 0.085 34.395 0.565 34.565 0.565 34.565 0.085 35.155 0.085 35.155 0.565 35.485 0.565 35.485 0.085 35.995 0.085 35.995 0.565 36.325 0.565 36.325 0.085 36.835 0.085 36.835 0.885 37.165 0.885 37.165 0.085 40.455 0.085 40.455 0.565 40.625 0.565 40.625 0.085 41.295 0.085 41.295 0.565 41.465 0.565 41.465 0.085 42.055 0.085 42.055 0.565 42.385 0.565 42.385 0.085 42.895 0.085 42.895 0.565 43.225 0.565 43.225 0.085 43.735 0.085 43.735 0.885 44.065 0.885 44.065 0.085 44.675 0.085 44.675 0.565 45.005 0.565 45.005 0.085 45.515 0.085 45.515 0.565 45.845 0.565 45.845 0.085 46.355 0.085 46.355 0.565 46.685 0.565 46.685 0.085 47.195 0.085 47.195 0.565 47.525 0.565 47.525 0.085 48.035 0.085 48.035 0.565 48.365 0.565 48.365 0.085 48.875 0.085 48.875 0.885 49.205 0.885 49.205 0.085 49.815 0.085 49.815 0.545 50.12 0.545 50.12 0.085 50.79 0.085 50.79 0.545 50.96 0.545 50.96 0.085 51.63 0.085 51.63 0.545 51.8 0.545 51.8 0.085 52.47 0.085 52.47 0.545 52.64 0.545 52.64 0.085 53.31 0.085 53.31 0.545 53.565 0.545 53.565 0.085 54.295 0.085 54.295 0.885 54.625 0.885 54.625 0.085 55.135 0.085 55.135 0.565 55.465 0.565 55.465 0.085 55.975 0.085 55.975 0.565 56.305 0.565 56.305 0.085 56.815 0.085 56.815 0.565 57.145 0.565 57.145 0.085 57.655 0.085 57.655 0.565 57.985 0.565 57.985 0.085 58.495 0.085 58.495 0.565 58.825 0.565 58.825 0.085 59.815 0.085 59.815 0.885 60.145 0.885 60.145 0.085 60.655 0.085 60.655 0.565 60.985 0.565 60.985 0.085 61.495 0.085 61.495 0.565 61.825 0.565 61.825 0.085 62.335 0.085 62.335 0.565 62.665 0.565 62.665 0.085 63.175 0.085 63.175 0.565 63.505 0.565 63.505 0.085 64.015 0.085 64.015 0.565 64.345 0.565 64.345 0.085 65.375 0.085 65.375 0.565 65.705 0.565 65.705 0.085 66.215 0.085 66.215 0.565 66.545 0.565 66.545 0.085 67.055 0.085 67.055 0.565 67.385 0.565 67.385 0.085 67.895 0.085 67.895 0.565 68.225 0.565 68.225 0.085 68.735 0.085 68.735 0.565 69.065 0.565 69.065 0.085 69.575 0.085 69.575 0.885 69.905 0.885 69.905 0.085 70.895 0.085 70.895 0.565 71.225 0.565 71.225 0.085 71.735 0.085 71.735 0.565 72.065 0.565 72.065 0.085 72.575 0.085 72.575 0.565 72.905 0.565 72.905 0.085 73.415 0.085 73.415 0.565 73.745 0.565 73.745 0.085 74.255 0.085 74.255 0.565 74.585 0.565 74.585 0.085 75.095 0.085 75.095 0.885 75.425 0.885 75.425 0.085 76.415 0.085 76.415 0.565 76.745 0.565 76.745 0.085 77.255 0.085 77.255 0.565 77.585 0.565 77.585 0.085 78.095 0.085 78.095 0.565 78.425 0.565 78.425 0.085 78.935 0.085 78.935 0.565 79.265 0.565 79.265 0.085 79.775 0.085 79.775 0.565 80.105 0.565 80.105 0.085 80.615 0.085 80.615 0.885 80.945 0.885 80.945 0.085 82.315 0.085 82.315 0.565 82.485 0.565 82.485 0.085 83.155 0.085 83.155 0.565 83.325 0.565 83.325 0.085 83.915 0.085 83.915 0.565 84.245 0.565 84.245 0.085 84.755 0.085 84.755 0.565 85.085 0.565 85.085 0.085 85.595 0.085 85.595 0.885 85.925 0.885 85.925 0.085 86.455 0.085 86.455 0.565 86.625 0.565 86.625 0.085 87.295 0.085 87.295 0.565 87.465 0.565 87.465 0.085 88.055 0.085 88.055 0.565 88.385 0.565 88.385 0.085 88.895 0.085 88.895 0.565 89.225 0.565 89.225 0.085 89.735 0.085 89.735 0.885 90.065 0.885 90.065 0.085 90.635 0.085 90.635 0.885 90.965 0.885 90.965 0.085 91.475 0.085 91.475 0.565 91.805 0.565 91.805 0.085 92.315 0.085 92.315 0.565 92.645 0.565 92.645 0.085 93.155 0.085 93.155 0.565 93.485 0.565 93.485 0.085 93.995 0.085 93.995 0.565 94.325 0.565 94.325 0.085 94.835 0.085 94.835 0.565 95.165 0.565 95.165 0.085 96.195 0.085 96.195 0.565 96.525 0.565 96.525 0.085 97.035 0.085 97.035 0.565 97.365 0.565 97.365 0.085 97.875 0.085 97.875 0.565 98.205 0.565 98.205 0.085 98.715 0.085 98.715 0.565 99.045 0.565 99.045 0.085 99.555 0.085 99.555 0.565 99.885 0.565 99.885 0.085 100.395 0.085 100.395 0.885 ;
      POLYGON 103.79 130.39 103.79 124.95 134.15 124.95 134.15 5.61 103.79 5.61 103.79 0.17 30.53 0.17 30.53 5.61 0.17 5.61 0.17 124.95 30.53 124.95 30.53 130.39 ;
    LAYER mcon ;
      RECT 59.025 130.475 59.195 130.645 ;
      RECT 58.565 130.475 58.735 130.645 ;
      RECT 58.105 130.475 58.275 130.645 ;
      RECT 57.645 130.475 57.815 130.645 ;
      RECT 57.185 130.475 57.355 130.645 ;
      RECT 56.725 130.475 56.895 130.645 ;
      RECT 56.265 130.475 56.435 130.645 ;
      RECT 55.805 130.475 55.975 130.645 ;
      RECT 55.345 130.475 55.515 130.645 ;
      RECT 54.885 130.475 55.055 130.645 ;
      RECT 54.425 130.475 54.595 130.645 ;
      RECT 53.965 130.475 54.135 130.645 ;
      RECT 128.485 5.355 128.655 5.525 ;
      RECT 128.025 5.355 128.195 5.525 ;
      RECT 127.565 5.355 127.735 5.525 ;
      RECT 127.105 5.355 127.275 5.525 ;
      RECT 126.645 5.355 126.815 5.525 ;
      RECT 126.185 5.355 126.355 5.525 ;
      RECT 125.725 5.355 125.895 5.525 ;
      RECT 125.265 5.355 125.435 5.525 ;
      RECT 124.805 5.355 124.975 5.525 ;
      RECT 124.345 5.355 124.515 5.525 ;
      RECT 123.885 5.355 124.055 5.525 ;
      RECT 123.425 5.355 123.595 5.525 ;
      RECT 122.965 5.355 123.135 5.525 ;
      RECT 122.505 5.355 122.675 5.525 ;
      RECT 122.045 5.355 122.215 5.525 ;
      RECT 121.585 5.355 121.755 5.525 ;
      RECT 121.125 5.355 121.295 5.525 ;
      RECT 120.665 5.355 120.835 5.525 ;
      RECT 120.205 5.355 120.375 5.525 ;
      RECT 119.745 5.355 119.915 5.525 ;
      RECT 119.285 5.355 119.455 5.525 ;
      RECT 118.825 5.355 118.995 5.525 ;
      RECT 118.365 5.355 118.535 5.525 ;
    LAYER via ;
      RECT 89.165 130.365 89.315 130.515 ;
      RECT 59.725 130.365 59.875 130.515 ;
      RECT 68.235 129.975 68.385 130.125 ;
      RECT 65.475 129.975 65.625 130.125 ;
      RECT 47.075 129.975 47.225 130.125 ;
      RECT 35.575 129.975 35.725 130.125 ;
      RECT 17.635 124.535 17.785 124.685 ;
      RECT 124.815 5.875 124.965 6.025 ;
      RECT 14.415 5.875 14.565 6.025 ;
      RECT 12.575 5.875 12.725 6.025 ;
      RECT 93.535 0.435 93.685 0.585 ;
      RECT 86.175 0.435 86.325 0.585 ;
      RECT 72.145 0.435 72.295 0.585 ;
      RECT 40.635 0.435 40.785 0.585 ;
      RECT 89.165 0.045 89.315 0.195 ;
      RECT 59.725 0.045 59.875 0.195 ;
    LAYER via2 ;
      RECT 89.14 130.34 89.34 130.54 ;
      RECT 59.7 130.34 59.9 130.54 ;
      RECT 101.33 130.12 101.53 130.32 ;
      RECT 90.75 130.12 90.95 130.32 ;
      RECT 83.85 130.12 84.05 130.32 ;
      RECT 70.51 130.12 70.71 130.32 ;
      RECT 1.05 24.04 1.25 24.24 ;
      RECT 120.65 5.68 120.85 5.88 ;
      RECT 109.15 5.68 109.35 5.88 ;
      RECT 12.09 5.68 12.29 5.88 ;
      RECT 95.81 0.24 96.01 0.44 ;
      RECT 86.61 0.24 86.81 0.44 ;
      RECT 64.07 0.24 64.27 0.44 ;
      RECT 48.89 0.24 49.09 0.44 ;
      RECT 89.14 0.02 89.34 0.22 ;
      RECT 59.7 0.02 59.9 0.22 ;
    LAYER via3 ;
      RECT 89.14 130.34 89.34 130.54 ;
      RECT 59.7 130.34 59.9 130.54 ;
      RECT 102.48 130.12 102.68 130.32 ;
      RECT 83.16 130.12 83.36 130.32 ;
      RECT 75.8 130.12 76 130.32 ;
      RECT 71.2 130.12 71.4 130.32 ;
      RECT 70.28 130.12 70.48 130.32 ;
      RECT 103.4 5.68 103.6 5.88 ;
      RECT 12.32 5.68 12.52 5.88 ;
      RECT 83.16 0.92 83.36 1.12 ;
      RECT 77.64 0.92 77.84 1.12 ;
      RECT 64.76 0.92 64.96 1.12 ;
      RECT 72.12 0.41 72.32 0.61 ;
      RECT 94.2 0.24 94.4 0.44 ;
      RECT 85 0.24 85.2 0.44 ;
      RECT 75.8 0.24 76 0.44 ;
      RECT 68.44 0.24 68.64 0.44 ;
      RECT 52.8 0.24 53 0.44 ;
      RECT 89.14 0.02 89.34 0.22 ;
      RECT 59.7 0.02 59.9 0.22 ;
    LAYER OVERLAP ;
      POLYGON 30.36 0 30.36 5.44 0 5.44 0 125.12 30.36 125.12 30.36 130.56 103.96 130.56 103.96 125.12 134.32 125.12 134.32 5.44 103.96 5.44 103.96 0 ;
  END
END sb_1__1_

END LIBRARY
