//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module sb_8__1_
(
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
    bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
    bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
    bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
    ccff_head,
    chanx_left_in,
    chany_bottom_in,
    chany_top_in,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_,
    pReset,
    prog_clk,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
    ccff_tail,
    chanx_left_out,
    chany_bottom_out,
    chany_top_out
);

    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
    input bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
    input bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
    input bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
    input bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
    input ccff_head;
    input [0:29]chanx_left_in;
    input [0:29]chany_bottom_in;
    input [0:29]chany_top_in;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_;
    input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_;
    input pReset;
    input prog_clk;
    input top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_;
    input top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_;
    input top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_;
    input top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_;
    input top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_;
    input top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_;
    input top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
    input top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
    input top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
    input top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
    input top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
    input top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
    output ccff_tail;
    output [0:29]chanx_left_out;
    output [0:29]chany_bottom_out;
    output [0:29]chany_top_out;

    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
    wire bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
    wire bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
    wire bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
    wire bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
    wire ccff_head;
    wire ccff_tail;
    wire [0:29]chanx_left_in;
    wire [0:29]chanx_left_out;
    wire [0:29]chany_bottom_in;
    wire [0:29]chany_bottom_out;
    wire [0:29]chany_top_in;
    wire [0:29]chany_top_out;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_;
    wire left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_;
    wire [0:3]mux_bottom_track_11_undriven_sram_inv;
    wire [0:2]mux_bottom_track_13_undriven_sram_inv;
    wire [0:3]mux_bottom_track_1_undriven_sram_inv;
    wire [0:2]mux_bottom_track_21_undriven_sram_inv;
    wire [0:2]mux_bottom_track_29_undriven_sram_inv;
    wire [0:2]mux_bottom_track_37_undriven_sram_inv;
    wire [0:3]mux_bottom_track_3_undriven_sram_inv;
    wire [0:2]mux_bottom_track_45_undriven_sram_inv;
    wire [0:2]mux_bottom_track_53_undriven_sram_inv;
    wire [0:3]mux_bottom_track_5_undriven_sram_inv;
    wire [0:3]mux_bottom_track_7_undriven_sram_inv;
    wire [0:2]mux_left_track_11_undriven_sram_inv;
    wire [0:2]mux_left_track_13_undriven_sram_inv;
    wire [0:2]mux_left_track_15_undriven_sram_inv;
    wire [0:2]mux_left_track_17_undriven_sram_inv;
    wire [0:2]mux_left_track_19_undriven_sram_inv;
    wire [0:2]mux_left_track_1_undriven_sram_inv;
    wire [0:2]mux_left_track_21_undriven_sram_inv;
    wire [0:2]mux_left_track_23_undriven_sram_inv;
    wire [0:1]mux_left_track_25_undriven_sram_inv;
    wire [0:1]mux_left_track_27_undriven_sram_inv;
    wire [0:1]mux_left_track_29_undriven_sram_inv;
    wire [0:1]mux_left_track_31_undriven_sram_inv;
    wire [0:1]mux_left_track_33_undriven_sram_inv;
    wire [0:1]mux_left_track_35_undriven_sram_inv;
    wire [0:1]mux_left_track_37_undriven_sram_inv;
    wire [0:2]mux_left_track_3_undriven_sram_inv;
    wire [0:1]mux_left_track_41_undriven_sram_inv;
    wire [0:1]mux_left_track_45_undriven_sram_inv;
    wire [0:1]mux_left_track_47_undriven_sram_inv;
    wire [0:1]mux_left_track_49_undriven_sram_inv;
    wire [0:1]mux_left_track_51_undriven_sram_inv;
    wire [0:1]mux_left_track_53_undriven_sram_inv;
    wire [0:1]mux_left_track_55_undriven_sram_inv;
    wire [0:1]mux_left_track_57_undriven_sram_inv;
    wire [0:2]mux_left_track_5_undriven_sram_inv;
    wire [0:2]mux_left_track_7_undriven_sram_inv;
    wire [0:2]mux_left_track_9_undriven_sram_inv;
    wire [0:3]mux_top_track_0_undriven_sram_inv;
    wire [0:3]mux_top_track_10_undriven_sram_inv;
    wire [0:2]mux_top_track_12_undriven_sram_inv;
    wire [0:2]mux_top_track_20_undriven_sram_inv;
    wire [0:2]mux_top_track_28_undriven_sram_inv;
    wire [0:3]mux_top_track_2_undriven_sram_inv;
    wire [0:2]mux_top_track_36_undriven_sram_inv;
    wire [0:2]mux_top_track_44_undriven_sram_inv;
    wire [0:3]mux_top_track_4_undriven_sram_inv;
    wire [0:2]mux_top_track_52_undriven_sram_inv;
    wire [0:3]mux_top_track_6_undriven_sram_inv;
    wire [0:3]mux_tree_tapbuf_size10_0_sram;
    wire mux_tree_tapbuf_size10_mem_0_ccff_tail;
    wire [0:3]mux_tree_tapbuf_size11_0_sram;
    wire [0:3]mux_tree_tapbuf_size11_1_sram;
    wire [0:3]mux_tree_tapbuf_size11_2_sram;
    wire mux_tree_tapbuf_size11_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size11_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size11_mem_2_ccff_tail;
    wire [0:1]mux_tree_tapbuf_size2_0_sram;
    wire [0:1]mux_tree_tapbuf_size2_1_sram;
    wire [0:1]mux_tree_tapbuf_size2_2_sram;
    wire [0:1]mux_tree_tapbuf_size2_3_sram;
    wire [0:1]mux_tree_tapbuf_size2_4_sram;
    wire [0:1]mux_tree_tapbuf_size2_5_sram;
    wire [0:1]mux_tree_tapbuf_size2_6_sram;
    wire mux_tree_tapbuf_size2_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_2_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_3_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_4_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_5_ccff_tail;
    wire [0:1]mux_tree_tapbuf_size3_0_sram;
    wire [0:1]mux_tree_tapbuf_size3_1_sram;
    wire [0:1]mux_tree_tapbuf_size3_2_sram;
    wire [0:1]mux_tree_tapbuf_size3_3_sram;
    wire [0:1]mux_tree_tapbuf_size3_4_sram;
    wire [0:1]mux_tree_tapbuf_size3_5_sram;
    wire [0:1]mux_tree_tapbuf_size3_6_sram;
    wire [0:1]mux_tree_tapbuf_size3_7_sram;
    wire mux_tree_tapbuf_size3_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_2_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_3_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_4_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_5_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_6_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_7_ccff_tail;
    wire [0:2]mux_tree_tapbuf_size4_0_sram;
    wire [0:2]mux_tree_tapbuf_size4_1_sram;
    wire [0:2]mux_tree_tapbuf_size4_2_sram;
    wire [0:2]mux_tree_tapbuf_size4_3_sram;
    wire [0:2]mux_tree_tapbuf_size4_4_sram;
    wire [0:2]mux_tree_tapbuf_size4_5_sram;
    wire mux_tree_tapbuf_size4_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size4_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size4_mem_2_ccff_tail;
    wire mux_tree_tapbuf_size4_mem_3_ccff_tail;
    wire mux_tree_tapbuf_size4_mem_4_ccff_tail;
    wire mux_tree_tapbuf_size4_mem_5_ccff_tail;
    wire [0:2]mux_tree_tapbuf_size5_0_sram;
    wire [0:2]mux_tree_tapbuf_size5_1_sram;
    wire [0:2]mux_tree_tapbuf_size5_2_sram;
    wire [0:2]mux_tree_tapbuf_size5_3_sram;
    wire mux_tree_tapbuf_size5_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_2_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_3_ccff_tail;
    wire [0:2]mux_tree_tapbuf_size6_0_sram;
    wire [0:2]mux_tree_tapbuf_size6_1_sram;
    wire [0:2]mux_tree_tapbuf_size6_2_sram;
    wire [0:2]mux_tree_tapbuf_size6_3_sram;
    wire [0:2]mux_tree_tapbuf_size6_4_sram;
    wire [0:2]mux_tree_tapbuf_size6_5_sram;
    wire [0:2]mux_tree_tapbuf_size6_6_sram;
    wire [0:2]mux_tree_tapbuf_size6_7_sram;
    wire [0:2]mux_tree_tapbuf_size6_8_sram;
    wire mux_tree_tapbuf_size6_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size6_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size6_mem_2_ccff_tail;
    wire mux_tree_tapbuf_size6_mem_3_ccff_tail;
    wire mux_tree_tapbuf_size6_mem_4_ccff_tail;
    wire mux_tree_tapbuf_size6_mem_5_ccff_tail;
    wire mux_tree_tapbuf_size6_mem_6_ccff_tail;
    wire mux_tree_tapbuf_size6_mem_7_ccff_tail;
    wire mux_tree_tapbuf_size6_mem_8_ccff_tail;
    wire [0:2]mux_tree_tapbuf_size7_0_sram;
    wire [0:2]mux_tree_tapbuf_size7_1_sram;
    wire [0:2]mux_tree_tapbuf_size7_2_sram;
    wire [0:2]mux_tree_tapbuf_size7_3_sram;
    wire [0:2]mux_tree_tapbuf_size7_4_sram;
    wire mux_tree_tapbuf_size7_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size7_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size7_mem_2_ccff_tail;
    wire mux_tree_tapbuf_size7_mem_3_ccff_tail;
    wire mux_tree_tapbuf_size7_mem_4_ccff_tail;
    wire [0:3]mux_tree_tapbuf_size8_0_sram;
    wire [0:3]mux_tree_tapbuf_size8_1_sram;
    wire mux_tree_tapbuf_size8_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size8_mem_1_ccff_tail;
    wire [0:3]mux_tree_tapbuf_size9_0_sram;
    wire [0:3]mux_tree_tapbuf_size9_1_sram;
    wire [0:3]mux_tree_tapbuf_size9_2_sram;
    wire [0:3]mux_tree_tapbuf_size9_3_sram;
    wire mux_tree_tapbuf_size9_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size9_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size9_mem_2_ccff_tail;
    wire mux_tree_tapbuf_size9_mem_3_ccff_tail;
    wire pReset;
    wire prog_clk;
    wire top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_;
    wire top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_;
    wire top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_;
    wire top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_;
    wire top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_;
    wire top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_;
    wire top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
    wire top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
    wire top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
    wire top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
    wire top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
    wire top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;

assign chanx_left_out[29] = chany_top_in[1];
assign chany_bottom_out[4] = chany_top_in[3];
assign chany_bottom_out[17] = chany_top_in[16];
assign chany_bottom_out[19] = chany_top_in[18];
assign chany_bottom_out[20] = chany_top_in[19];
assign chany_bottom_out[21] = chany_top_in[20];
assign chany_bottom_out[23] = chany_top_in[22];
assign chany_bottom_out[24] = chany_top_in[23];
assign chany_bottom_out[25] = chany_top_in[24];
assign chanx_left_out[21] = chany_top_in[25];
assign chany_bottom_out[27] = chany_top_in[26];
assign chany_bottom_out[28] = chany_top_in[27];
assign chany_bottom_out[7] = chany_top_in[6];
assign chany_bottom_out[29] = chany_top_in[28];
assign chany_top_out[4] = chany_bottom_in[3];
assign chany_top_out[7] = chany_bottom_in[6];
assign chany_top_out[8] = chany_bottom_in[7];
assign chany_top_out[9] = chany_bottom_in[8];
assign chany_top_out[11] = chany_bottom_in[10];
assign chany_top_out[12] = chany_bottom_in[11];
assign chany_top_out[13] = chany_bottom_in[12];
assign chany_top_out[15] = chany_bottom_in[14];
assign chany_top_out[16] = chany_bottom_in[15];
assign chany_bottom_out[8] = chany_top_in[7];
assign chany_top_out[17] = chany_bottom_in[16];
assign chany_top_out[19] = chany_bottom_in[18];
assign chany_top_out[20] = chany_bottom_in[19];
assign chany_top_out[21] = chany_bottom_in[20];
assign chany_top_out[23] = chany_bottom_in[22];
assign chany_top_out[24] = chany_bottom_in[23];
assign chany_top_out[25] = chany_bottom_in[24];
assign chany_top_out[27] = chany_bottom_in[26];
assign chany_top_out[28] = chany_bottom_in[27];
assign chany_top_out[29] = chany_bottom_in[28];
assign chany_bottom_out[9] = chany_top_in[8];
assign chanx_left_out[19] = left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
assign chany_bottom_out[11] = chany_top_in[10];
assign chany_bottom_out[12] = chany_top_in[11];
assign chany_bottom_out[13] = chany_top_in[12];
assign chany_bottom_out[15] = chany_top_in[14];
assign chany_bottom_out[16] = chany_top_in[15];
    mux_tree_tapbuf_size9_mem mem_bottom_track_1
    (
        .ccff_head(mux_tree_tapbuf_size6_mem_2_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size9_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size9_1_sram)
    );
    mux_tree_tapbuf_size11_mem mem_bottom_track_11
    (
        .ccff_head(mux_tree_tapbuf_size11_mem_1_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size11_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size11_2_sram)
    );
    mux_tree_tapbuf_size7_mem mem_bottom_track_13
    (
        .ccff_head(mux_tree_tapbuf_size11_mem_2_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size7_mem_3_ccff_tail),
        .mem_out(mux_tree_tapbuf_size7_3_sram)
    );
    mux_tree_tapbuf_size7_mem mem_bottom_track_21
    (
        .ccff_head(mux_tree_tapbuf_size7_mem_3_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size7_mem_4_ccff_tail),
        .mem_out(mux_tree_tapbuf_size7_4_sram)
    );
    mux_tree_tapbuf_size6_mem mem_bottom_track_29
    (
        .ccff_head(mux_tree_tapbuf_size7_mem_4_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size6_mem_3_ccff_tail),
        .mem_out(mux_tree_tapbuf_size6_3_sram)
    );
    mux_tree_tapbuf_size9_mem mem_bottom_track_3
    (
        .ccff_head(mux_tree_tapbuf_size9_mem_1_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size9_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size9_2_sram)
    );
    mux_tree_tapbuf_size5_mem mem_bottom_track_37
    (
        .ccff_head(mux_tree_tapbuf_size6_mem_3_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_0_sram)
    );
    mux_tree_tapbuf_size5_mem mem_bottom_track_45
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_1_sram)
    );
    mux_tree_tapbuf_size9_mem mem_bottom_track_5
    (
        .ccff_head(mux_tree_tapbuf_size9_mem_2_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size9_mem_3_ccff_tail),
        .mem_out(mux_tree_tapbuf_size9_3_sram)
    );
    mux_tree_tapbuf_size6_mem mem_bottom_track_53
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size6_mem_4_ccff_tail),
        .mem_out(mux_tree_tapbuf_size6_4_sram)
    );
    mux_tree_tapbuf_size11_mem mem_bottom_track_7
    (
        .ccff_head(mux_tree_tapbuf_size9_mem_3_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size11_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size11_1_sram)
    );
    mux_tree_tapbuf_size6_mem mem_left_track_1
    (
        .ccff_head(mux_tree_tapbuf_size6_mem_4_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size6_mem_5_ccff_tail),
        .mem_out(mux_tree_tapbuf_size6_5_sram)
    );
    mux_tree_tapbuf_size5_mem mem_left_track_11
    (
        .ccff_head(mux_tree_tapbuf_size6_mem_8_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_3_sram)
    );
    mux_tree_tapbuf_size4_mem mem_left_track_13
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size4_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size4_0_sram)
    );
    mux_tree_tapbuf_size4_mem mem_left_track_15
    (
        .ccff_head(mux_tree_tapbuf_size4_mem_0_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size4_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size4_1_sram)
    );
    mux_tree_tapbuf_size4_mem mem_left_track_17
    (
        .ccff_head(mux_tree_tapbuf_size4_mem_1_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size4_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size4_2_sram)
    );
    mux_tree_tapbuf_size4_mem mem_left_track_19
    (
        .ccff_head(mux_tree_tapbuf_size4_mem_2_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size4_mem_3_ccff_tail),
        .mem_out(mux_tree_tapbuf_size4_3_sram)
    );
    mux_tree_tapbuf_size4_mem mem_left_track_21
    (
        .ccff_head(mux_tree_tapbuf_size4_mem_3_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size4_mem_4_ccff_tail),
        .mem_out(mux_tree_tapbuf_size4_4_sram)
    );
    mux_tree_tapbuf_size4_mem mem_left_track_23
    (
        .ccff_head(mux_tree_tapbuf_size4_mem_4_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size4_mem_5_ccff_tail),
        .mem_out(mux_tree_tapbuf_size4_5_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_25
    (
        .ccff_head(mux_tree_tapbuf_size4_mem_5_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_0_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_27
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_0_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_1_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_29
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_1_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_2_sram)
    );
    mux_tree_tapbuf_size6_mem mem_left_track_3
    (
        .ccff_head(mux_tree_tapbuf_size6_mem_5_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size6_mem_6_ccff_tail),
        .mem_out(mux_tree_tapbuf_size6_6_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_31
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_2_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_3_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_3_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_33
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_3_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_4_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_4_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_35
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_4_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_5_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_5_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_37
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_5_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_6_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_6_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_41
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_6_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_0_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_45
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_0_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_1_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_47
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_1_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_2_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_49
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_2_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_3_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_3_sram)
    );
    mux_tree_tapbuf_size5_mem mem_left_track_5
    (
        .ccff_head(mux_tree_tapbuf_size6_mem_6_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_2_sram)
    );
    mux_tree_tapbuf_size3_mem mem_left_track_51
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_3_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size3_mem_7_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_7_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_53
    (
        .ccff_head(mux_tree_tapbuf_size3_mem_7_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_4_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_4_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_55
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_4_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size2_mem_5_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_5_sram)
    );
    mux_tree_tapbuf_size2_mem mem_left_track_57
    (
        .ccff_head(mux_tree_tapbuf_size2_mem_5_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_6_sram)
    );
    mux_tree_tapbuf_size6_mem mem_left_track_7
    (
        .ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size6_mem_7_ccff_tail),
        .mem_out(mux_tree_tapbuf_size6_7_sram)
    );
    mux_tree_tapbuf_size6_mem mem_left_track_9
    (
        .ccff_head(mux_tree_tapbuf_size6_mem_7_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size6_mem_8_ccff_tail),
        .mem_out(mux_tree_tapbuf_size6_8_sram)
    );
    mux_tree_tapbuf_size9_mem mem_top_track_0
    (
        .ccff_head(ccff_head),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size9_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size9_0_sram)
    );
    mux_tree_tapbuf_size11_mem mem_top_track_10
    (
        .ccff_head(mux_tree_tapbuf_size10_mem_0_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size11_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size11_0_sram)
    );
    mux_tree_tapbuf_size7_mem mem_top_track_12
    (
        .ccff_head(mux_tree_tapbuf_size11_mem_0_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size7_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size7_0_sram)
    );
    mux_tree_tapbuf_size8_mem mem_top_track_2
    (
        .ccff_head(mux_tree_tapbuf_size9_mem_0_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size8_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size8_0_sram)
    );
    mux_tree_tapbuf_size7_mem mem_top_track_20
    (
        .ccff_head(mux_tree_tapbuf_size7_mem_0_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size7_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size7_1_sram)
    );
    mux_tree_tapbuf_size7_mem mem_top_track_28
    (
        .ccff_head(mux_tree_tapbuf_size7_mem_1_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size7_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size7_2_sram)
    );
    mux_tree_tapbuf_size6_mem mem_top_track_36
    (
        .ccff_head(mux_tree_tapbuf_size7_mem_2_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size6_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size6_0_sram)
    );
    mux_tree_tapbuf_size8_mem mem_top_track_4
    (
        .ccff_head(mux_tree_tapbuf_size8_mem_0_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size8_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size8_1_sram)
    );
    mux_tree_tapbuf_size6_mem mem_top_track_44
    (
        .ccff_head(mux_tree_tapbuf_size6_mem_0_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size6_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size6_1_sram)
    );
    mux_tree_tapbuf_size6_mem mem_top_track_52
    (
        .ccff_head(mux_tree_tapbuf_size6_mem_1_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size6_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size6_2_sram)
    );
    mux_tree_tapbuf_size10_mem mem_top_track_6
    (
        .ccff_head(mux_tree_tapbuf_size8_mem_1_ccff_tail),
        .pReset(pReset),
        .prog_clk(prog_clk),
        .ccff_tail(mux_tree_tapbuf_size10_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size10_0_sram)
    );
    mux_tree_tapbuf_size9 mux_bottom_track_1
    (
        .in({chany_top_in[3], chany_top_in[19], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[1], chanx_left_in[12], chanx_left_in[23]}),
        .sram(mux_tree_tapbuf_size9_1_sram),
        .sram_inv(mux_bottom_track_1_undriven_sram_inv),
        .out(chany_bottom_out[0])
    );
    mux_tree_tapbuf_size11 mux_bottom_track_11
    (
        .in({chany_top_in[10], chany_top_in[24], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[5], chanx_left_in[16], chanx_left_in[27]}),
        .sram(mux_tree_tapbuf_size11_2_sram),
        .sram_inv(mux_bottom_track_11_undriven_sram_inv),
        .out(chany_bottom_out[5])
    );
    mux_tree_tapbuf_size7 mux_bottom_track_13
    (
        .in({chany_top_in[11], chany_top_in[26], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, chanx_left_in[6], chanx_left_in[17], chanx_left_in[28]}),
        .sram(mux_tree_tapbuf_size7_3_sram),
        .sram_inv(mux_bottom_track_13_undriven_sram_inv),
        .out(chany_bottom_out[6])
    );
    mux_tree_tapbuf_size7 mux_bottom_track_21
    (
        .in({chany_top_in[12], chany_top_in[27], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, chanx_left_in[7], chanx_left_in[18], chanx_left_in[29]}),
        .sram(mux_tree_tapbuf_size7_4_sram),
        .sram_inv(mux_bottom_track_21_undriven_sram_inv),
        .out(chany_bottom_out[10])
    );
    mux_tree_tapbuf_size6 mux_bottom_track_29
    (
        .in({chany_top_in[14], chany_top_in[28], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, chanx_left_in[8], chanx_left_in[19]}),
        .sram(mux_tree_tapbuf_size6_3_sram),
        .sram_inv(mux_bottom_track_29_undriven_sram_inv),
        .out(chany_bottom_out[14])
    );
    mux_tree_tapbuf_size9 mux_bottom_track_3
    (
        .in({chany_top_in[6], chany_top_in[20], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, chanx_left_in[2], chanx_left_in[13], chanx_left_in[24]}),
        .sram(mux_tree_tapbuf_size9_2_sram),
        .sram_inv(mux_bottom_track_3_undriven_sram_inv),
        .out(chany_bottom_out[1])
    );
    mux_tree_tapbuf_size5 mux_bottom_track_37
    (
        .in({chany_top_in[15], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[9], chanx_left_in[20]}),
        .sram(mux_tree_tapbuf_size5_0_sram),
        .sram_inv(mux_bottom_track_37_undriven_sram_inv),
        .out(chany_bottom_out[18])
    );
    mux_tree_tapbuf_size5 mux_bottom_track_45
    (
        .in({chany_top_in[16], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, chanx_left_in[10], chanx_left_in[21]}),
        .sram(mux_tree_tapbuf_size5_1_sram),
        .sram_inv(mux_bottom_track_45_undriven_sram_inv),
        .out(chany_bottom_out[22])
    );
    mux_tree_tapbuf_size9 mux_bottom_track_5
    (
        .in({chany_top_in[7], chany_top_in[22], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[3], chanx_left_in[14], chanx_left_in[25]}),
        .sram(mux_tree_tapbuf_size9_3_sram),
        .sram_inv(mux_bottom_track_5_undriven_sram_inv),
        .out(chany_bottom_out[2])
    );
    mux_tree_tapbuf_size6 mux_bottom_track_53
    (
        .in({chany_top_in[18], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[0], chanx_left_in[11], chanx_left_in[22]}),
        .sram(mux_tree_tapbuf_size6_4_sram),
        .sram_inv(mux_bottom_track_53_undriven_sram_inv),
        .out(chany_bottom_out[26])
    );
    mux_tree_tapbuf_size11 mux_bottom_track_7
    (
        .in({chany_top_in[8], chany_top_in[23], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, chanx_left_in[4], chanx_left_in[15], chanx_left_in[26]}),
        .sram(mux_tree_tapbuf_size11_1_sram),
        .sram_inv(mux_bottom_track_7_undriven_sram_inv),
        .out(chany_bottom_out[3])
    );
    mux_tree_tapbuf_size6 mux_left_track_1
    (
        .in({chany_top_in[0], chany_top_in[3], chany_bottom_in[3], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
        .sram(mux_tree_tapbuf_size6_5_sram),
        .sram_inv(mux_left_track_1_undriven_sram_inv),
        .out(chanx_left_out[0])
    );
    mux_tree_tapbuf_size5 mux_left_track_11
    (
        .in({chany_top_in[11], chany_bottom_in[5], chany_bottom_in[11], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
        .sram(mux_tree_tapbuf_size5_3_sram),
        .sram_inv(mux_left_track_11_undriven_sram_inv),
        .out(chanx_left_out[5])
    );
    mux_tree_tapbuf_size4 mux_left_track_13
    (
        .in({chany_top_in[12], chany_bottom_in[9], chany_bottom_in[12], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
        .sram(mux_tree_tapbuf_size4_0_sram),
        .sram_inv(mux_left_track_13_undriven_sram_inv),
        .out(chanx_left_out[6])
    );
    mux_tree_tapbuf_size4 mux_left_track_15
    (
        .in({chany_top_in[14], chany_bottom_in[13], chany_bottom_in[14], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_}),
        .sram(mux_tree_tapbuf_size4_1_sram),
        .sram_inv(mux_left_track_15_undriven_sram_inv),
        .out(chanx_left_out[7])
    );
    mux_tree_tapbuf_size4 mux_left_track_17
    (
        .in({chany_top_in[15], chany_bottom_in[15], chany_bottom_in[17], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
        .sram(mux_tree_tapbuf_size4_2_sram),
        .sram_inv(mux_left_track_17_undriven_sram_inv),
        .out(chanx_left_out[8])
    );
    mux_tree_tapbuf_size4 mux_left_track_19
    (
        .in({chany_top_in[16], chany_bottom_in[16], chany_bottom_in[21], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_}),
        .sram(mux_tree_tapbuf_size4_3_sram),
        .sram_inv(mux_left_track_19_undriven_sram_inv),
        .out(chanx_left_out[9])
    );
    mux_tree_tapbuf_size4 mux_left_track_21
    (
        .in({chany_top_in[18], chany_bottom_in[18], chany_bottom_in[25], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
        .sram(mux_tree_tapbuf_size4_4_sram),
        .sram_inv(mux_left_track_21_undriven_sram_inv),
        .out(chanx_left_out[10])
    );
    mux_tree_tapbuf_size4 mux_left_track_23
    (
        .in({chany_top_in[19], chany_bottom_in[19], chany_bottom_in[29], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
        .sram(mux_tree_tapbuf_size4_5_sram),
        .sram_inv(mux_left_track_23_undriven_sram_inv),
        .out(chanx_left_out[11])
    );
    mux_tree_tapbuf_size3 mux_left_track_25
    (
        .in({chany_top_in[20], chany_bottom_in[20], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
        .sram(mux_tree_tapbuf_size3_0_sram),
        .sram_inv(mux_left_track_25_undriven_sram_inv),
        .out(chanx_left_out[12])
    );
    mux_tree_tapbuf_size3 mux_left_track_27
    (
        .in({chany_top_in[22], chany_bottom_in[22], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_}),
        .sram(mux_tree_tapbuf_size3_1_sram),
        .sram_inv(mux_left_track_27_undriven_sram_inv),
        .out(chanx_left_out[13])
    );
    mux_tree_tapbuf_size3 mux_left_track_29
    (
        .in({chany_top_in[23], chany_bottom_in[23], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
        .sram(mux_tree_tapbuf_size3_2_sram),
        .sram_inv(mux_left_track_29_undriven_sram_inv),
        .out(chanx_left_out[14])
    );
    mux_tree_tapbuf_size6 mux_left_track_3
    (
        .in({chany_top_in[6], chany_bottom_in[0], chany_bottom_in[6], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_}),
        .sram(mux_tree_tapbuf_size6_6_sram),
        .sram_inv(mux_left_track_3_undriven_sram_inv),
        .out(chanx_left_out[1])
    );
    mux_tree_tapbuf_size3 mux_left_track_31
    (
        .in({chany_top_in[24], chany_bottom_in[24], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_}),
        .sram(mux_tree_tapbuf_size3_3_sram),
        .sram_inv(mux_left_track_31_undriven_sram_inv),
        .out(chanx_left_out[15])
    );
    mux_tree_tapbuf_size3 mux_left_track_33
    (
        .in({chany_top_in[26], chany_bottom_in[26], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
        .sram(mux_tree_tapbuf_size3_4_sram),
        .sram_inv(mux_left_track_33_undriven_sram_inv),
        .out(chanx_left_out[16])
    );
    mux_tree_tapbuf_size3 mux_left_track_35
    (
        .in({chany_top_in[27], chany_bottom_in[27], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_}),
        .sram(mux_tree_tapbuf_size3_5_sram),
        .sram_inv(mux_left_track_35_undriven_sram_inv),
        .out(chanx_left_out[17])
    );
    mux_tree_tapbuf_size3 mux_left_track_37
    (
        .in({chany_top_in[28], chany_bottom_in[28], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
        .sram(mux_tree_tapbuf_size3_6_sram),
        .sram_inv(mux_left_track_37_undriven_sram_inv),
        .out(chanx_left_out[18])
    );
    mux_tree_tapbuf_size2 mux_left_track_41
    (
        .in({chany_top_in[29], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
        .sram(mux_tree_tapbuf_size2_0_sram),
        .sram_inv(mux_left_track_41_undriven_sram_inv),
        .out(chanx_left_out[20])
    );
    mux_tree_tapbuf_size2 mux_left_track_45
    (
        .in({chany_top_in[21], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
        .sram(mux_tree_tapbuf_size2_1_sram),
        .sram_inv(mux_left_track_45_undriven_sram_inv),
        .out(chanx_left_out[22])
    );
    mux_tree_tapbuf_size2 mux_left_track_47
    (
        .in({chany_top_in[17], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_}),
        .sram(mux_tree_tapbuf_size2_2_sram),
        .sram_inv(mux_left_track_47_undriven_sram_inv),
        .out(chanx_left_out[23])
    );
    mux_tree_tapbuf_size2 mux_left_track_49
    (
        .in({chany_top_in[13], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
        .sram(mux_tree_tapbuf_size2_3_sram),
        .sram_inv(mux_left_track_49_undriven_sram_inv),
        .out(chanx_left_out[24])
    );
    mux_tree_tapbuf_size5 mux_left_track_5
    (
        .in({chany_top_in[7], chany_bottom_in[1], chany_bottom_in[7], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
        .sram(mux_tree_tapbuf_size5_2_sram),
        .sram_inv(mux_left_track_5_undriven_sram_inv),
        .out(chanx_left_out[2])
    );
    mux_tree_tapbuf_size3 mux_left_track_51
    (
        .in({chany_top_in[9], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_}),
        .sram(mux_tree_tapbuf_size3_7_sram),
        .sram_inv(mux_left_track_51_undriven_sram_inv),
        .out(chanx_left_out[25])
    );
    mux_tree_tapbuf_size2 mux_left_track_53
    (
        .in({chany_top_in[5], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
        .sram(mux_tree_tapbuf_size2_4_sram),
        .sram_inv(mux_left_track_53_undriven_sram_inv),
        .out(chanx_left_out[26])
    );
    mux_tree_tapbuf_size2 mux_left_track_55
    (
        .in({chany_top_in[4], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
        .sram(mux_tree_tapbuf_size2_5_sram),
        .sram_inv(mux_left_track_55_undriven_sram_inv),
        .out(chanx_left_out[27])
    );
    mux_tree_tapbuf_size2 mux_left_track_57
    (
        .in({chany_top_in[2], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
        .sram(mux_tree_tapbuf_size2_6_sram),
        .sram_inv(mux_left_track_57_undriven_sram_inv),
        .out(chanx_left_out[28])
    );
    mux_tree_tapbuf_size6 mux_left_track_7
    (
        .in({chany_top_in[8], chany_bottom_in[2], chany_bottom_in[8], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
        .sram(mux_tree_tapbuf_size6_7_sram),
        .sram_inv(mux_left_track_7_undriven_sram_inv),
        .out(chanx_left_out[3])
    );
    mux_tree_tapbuf_size6 mux_left_track_9
    (
        .in({chany_top_in[10], chany_bottom_in[4], chany_bottom_in[10], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_}),
        .sram(mux_tree_tapbuf_size6_8_sram),
        .sram_inv(mux_left_track_9_undriven_sram_inv),
        .out(chanx_left_out[4])
    );
    mux_tree_tapbuf_size9 mux_top_track_0
    (
        .in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[3], chany_bottom_in[19], chanx_left_in[0], chanx_left_in[11], chanx_left_in[22]}),
        .sram(mux_tree_tapbuf_size9_0_sram),
        .sram_inv(mux_top_track_0_undriven_sram_inv),
        .out(chany_top_out[0])
    );
    mux_tree_tapbuf_size11 mux_top_track_10
    (
        .in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[10], chany_bottom_in[24], chanx_left_in[7], chanx_left_in[18], chanx_left_in[29]}),
        .sram(mux_tree_tapbuf_size11_0_sram),
        .sram_inv(mux_top_track_10_undriven_sram_inv),
        .out(chany_top_out[5])
    );
    mux_tree_tapbuf_size7 mux_top_track_12
    (
        .in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, chany_bottom_in[11], chany_bottom_in[26], chanx_left_in[6], chanx_left_in[17], chanx_left_in[28]}),
        .sram(mux_tree_tapbuf_size7_0_sram),
        .sram_inv(mux_top_track_12_undriven_sram_inv),
        .out(chany_top_out[6])
    );
    mux_tree_tapbuf_size8 mux_top_track_2
    (
        .in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[6], chany_bottom_in[20], chanx_left_in[10], chanx_left_in[21]}),
        .sram(mux_tree_tapbuf_size8_0_sram),
        .sram_inv(mux_top_track_2_undriven_sram_inv),
        .out(chany_top_out[1])
    );
    mux_tree_tapbuf_size7 mux_top_track_20
    (
        .in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, chany_bottom_in[12], chany_bottom_in[27], chanx_left_in[5], chanx_left_in[16], chanx_left_in[27]}),
        .sram(mux_tree_tapbuf_size7_1_sram),
        .sram_inv(mux_top_track_20_undriven_sram_inv),
        .out(chany_top_out[10])
    );
    mux_tree_tapbuf_size7 mux_top_track_28
    (
        .in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[14], chany_bottom_in[28], chanx_left_in[4], chanx_left_in[15], chanx_left_in[26]}),
        .sram(mux_tree_tapbuf_size7_2_sram),
        .sram_inv(mux_top_track_28_undriven_sram_inv),
        .out(chany_top_out[14])
    );
    mux_tree_tapbuf_size6 mux_top_track_36
    (
        .in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[15], chanx_left_in[3], chanx_left_in[14], chanx_left_in[25]}),
        .sram(mux_tree_tapbuf_size6_0_sram),
        .sram_inv(mux_top_track_36_undriven_sram_inv),
        .out(chany_top_out[18])
    );
    mux_tree_tapbuf_size8 mux_top_track_4
    (
        .in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[7], chany_bottom_in[22], chanx_left_in[9], chanx_left_in[20]}),
        .sram(mux_tree_tapbuf_size8_1_sram),
        .sram_inv(mux_top_track_4_undriven_sram_inv),
        .out(chany_top_out[2])
    );
    mux_tree_tapbuf_size6 mux_top_track_44
    (
        .in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[16], chanx_left_in[2], chanx_left_in[13], chanx_left_in[24]}),
        .sram(mux_tree_tapbuf_size6_1_sram),
        .sram_inv(mux_top_track_44_undriven_sram_inv),
        .out(chany_top_out[22])
    );
    mux_tree_tapbuf_size6 mux_top_track_52
    (
        .in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[18], chanx_left_in[1], chanx_left_in[12], chanx_left_in[23]}),
        .sram(mux_tree_tapbuf_size6_2_sram),
        .sram_inv(mux_top_track_52_undriven_sram_inv),
        .out(chany_top_out[26])
    );
    mux_tree_tapbuf_size10 mux_top_track_6
    (
        .in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[8], chany_bottom_in[23], chanx_left_in[8], chanx_left_in[19]}),
        .sram(mux_tree_tapbuf_size10_0_sram),
        .sram_inv(mux_top_track_6_undriven_sram_inv),
        .out(chany_top_out[3])
    );
endmodule

