//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module sb_0__8_
(
    prog_reset,
    prog_clk,
    chanx_right_in,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_,
    chany_bottom_in,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
    ccff_head,
    chanx_right_out,
    chany_bottom_out,
    ccff_tail
);

    input prog_reset;
    input prog_clk;
    input [0:29]chanx_right_in;
    input right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
    input right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
    input right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
    input right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
    input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
    input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
    input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
    input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
    input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
    input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
    input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_;
    input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_;
    input [0:29]chany_bottom_in;
    input bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
    input bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
    input bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
    input bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
    input ccff_head;
    output [0:29]chanx_right_out;
    output [0:29]chany_bottom_out;
    output ccff_tail;

    wire prog_reset;
    wire prog_clk;
    wire [0:29]chanx_right_in;
    wire right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
    wire right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
    wire right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
    wire right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
    wire right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
    wire right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
    wire right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
    wire right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
    wire right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
    wire right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
    wire right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_;
    wire right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_;
    wire [0:29]chany_bottom_in;
    wire bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
    wire bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
    wire bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
    wire bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
    wire ccff_head;
    wire [0:29]chanx_right_out;
    wire [0:29]chany_bottom_out;
    wire ccff_tail;
    wire [0:1]mux_bottom_track_11_undriven_sram_inv;
    wire [0:1]mux_bottom_track_13_undriven_sram_inv;
    wire [0:1]mux_bottom_track_15_undriven_sram_inv;
    wire [0:1]mux_bottom_track_17_undriven_sram_inv;
    wire [0:1]mux_bottom_track_19_undriven_sram_inv;
    wire [0:1]mux_bottom_track_1_undriven_sram_inv;
    wire [0:1]mux_bottom_track_29_undriven_sram_inv;
    wire [0:1]mux_bottom_track_31_undriven_sram_inv;
    wire [0:1]mux_bottom_track_33_undriven_sram_inv;
    wire [0:1]mux_bottom_track_35_undriven_sram_inv;
    wire [0:1]mux_bottom_track_3_undriven_sram_inv;
    wire [0:1]mux_bottom_track_45_undriven_sram_inv;
    wire [0:1]mux_bottom_track_47_undriven_sram_inv;
    wire [0:1]mux_bottom_track_49_undriven_sram_inv;
    wire [0:1]mux_bottom_track_51_undriven_sram_inv;
    wire [0:1]mux_bottom_track_5_undriven_sram_inv;
    wire [0:1]mux_bottom_track_7_undriven_sram_inv;
    wire [0:1]mux_bottom_track_9_undriven_sram_inv;
    wire [0:2]mux_right_track_0_undriven_sram_inv;
    wire [0:2]mux_right_track_10_undriven_sram_inv;
    wire [0:1]mux_right_track_12_undriven_sram_inv;
    wire [0:1]mux_right_track_14_undriven_sram_inv;
    wire [0:1]mux_right_track_16_undriven_sram_inv;
    wire [0:1]mux_right_track_18_undriven_sram_inv;
    wire [0:1]mux_right_track_20_undriven_sram_inv;
    wire [0:1]mux_right_track_22_undriven_sram_inv;
    wire [0:1]mux_right_track_24_undriven_sram_inv;
    wire [0:1]mux_right_track_26_undriven_sram_inv;
    wire [0:1]mux_right_track_28_undriven_sram_inv;
    wire [0:2]mux_right_track_2_undriven_sram_inv;
    wire [0:1]mux_right_track_30_undriven_sram_inv;
    wire [0:1]mux_right_track_32_undriven_sram_inv;
    wire [0:1]mux_right_track_34_undriven_sram_inv;
    wire [0:1]mux_right_track_36_undriven_sram_inv;
    wire [0:1]mux_right_track_38_undriven_sram_inv;
    wire [0:1]mux_right_track_40_undriven_sram_inv;
    wire [0:1]mux_right_track_42_undriven_sram_inv;
    wire [0:1]mux_right_track_44_undriven_sram_inv;
    wire [0:1]mux_right_track_46_undriven_sram_inv;
    wire [0:1]mux_right_track_48_undriven_sram_inv;
    wire [0:2]mux_right_track_4_undriven_sram_inv;
    wire [0:1]mux_right_track_50_undriven_sram_inv;
    wire [0:1]mux_right_track_52_undriven_sram_inv;
    wire [0:1]mux_right_track_54_undriven_sram_inv;
    wire [0:1]mux_right_track_56_undriven_sram_inv;
    wire [0:1]mux_right_track_58_undriven_sram_inv;
    wire [0:2]mux_right_track_6_undriven_sram_inv;
    wire [0:2]mux_right_track_8_undriven_sram_inv;
    wire [0:1]mux_tree_tapbuf_size2_0_sram;
    wire [0:1]mux_tree_tapbuf_size2_10_sram;
    wire [0:1]mux_tree_tapbuf_size2_11_sram;
    wire [0:1]mux_tree_tapbuf_size2_12_sram;
    wire [0:1]mux_tree_tapbuf_size2_13_sram;
    wire [0:1]mux_tree_tapbuf_size2_14_sram;
    wire [0:1]mux_tree_tapbuf_size2_15_sram;
    wire [0:1]mux_tree_tapbuf_size2_16_sram;
    wire [0:1]mux_tree_tapbuf_size2_17_sram;
    wire [0:1]mux_tree_tapbuf_size2_18_sram;
    wire [0:1]mux_tree_tapbuf_size2_19_sram;
    wire [0:1]mux_tree_tapbuf_size2_1_sram;
    wire [0:1]mux_tree_tapbuf_size2_20_sram;
    wire [0:1]mux_tree_tapbuf_size2_21_sram;
    wire [0:1]mux_tree_tapbuf_size2_22_sram;
    wire [0:1]mux_tree_tapbuf_size2_23_sram;
    wire [0:1]mux_tree_tapbuf_size2_24_sram;
    wire [0:1]mux_tree_tapbuf_size2_25_sram;
    wire [0:1]mux_tree_tapbuf_size2_26_sram;
    wire [0:1]mux_tree_tapbuf_size2_27_sram;
    wire [0:1]mux_tree_tapbuf_size2_28_sram;
    wire [0:1]mux_tree_tapbuf_size2_2_sram;
    wire [0:1]mux_tree_tapbuf_size2_3_sram;
    wire [0:1]mux_tree_tapbuf_size2_4_sram;
    wire [0:1]mux_tree_tapbuf_size2_5_sram;
    wire [0:1]mux_tree_tapbuf_size2_6_sram;
    wire [0:1]mux_tree_tapbuf_size2_7_sram;
    wire [0:1]mux_tree_tapbuf_size2_8_sram;
    wire [0:1]mux_tree_tapbuf_size2_9_sram;
    wire mux_tree_tapbuf_size2_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_10_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_11_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_12_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_13_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_14_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_15_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_16_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_17_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_18_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_19_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_20_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_21_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_22_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_23_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_24_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_25_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_26_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_27_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_2_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_3_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_4_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_5_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_6_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_7_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_8_ccff_tail;
    wire mux_tree_tapbuf_size2_mem_9_ccff_tail;
    wire [0:1]mux_tree_tapbuf_size3_0_sram;
    wire [0:1]mux_tree_tapbuf_size3_10_sram;
    wire [0:1]mux_tree_tapbuf_size3_11_sram;
    wire [0:1]mux_tree_tapbuf_size3_12_sram;
    wire [0:1]mux_tree_tapbuf_size3_1_sram;
    wire [0:1]mux_tree_tapbuf_size3_2_sram;
    wire [0:1]mux_tree_tapbuf_size3_3_sram;
    wire [0:1]mux_tree_tapbuf_size3_4_sram;
    wire [0:1]mux_tree_tapbuf_size3_5_sram;
    wire [0:1]mux_tree_tapbuf_size3_6_sram;
    wire [0:1]mux_tree_tapbuf_size3_7_sram;
    wire [0:1]mux_tree_tapbuf_size3_8_sram;
    wire [0:1]mux_tree_tapbuf_size3_9_sram;
    wire mux_tree_tapbuf_size3_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_10_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_11_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_12_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_2_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_3_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_4_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_5_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_6_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_7_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_8_ccff_tail;
    wire mux_tree_tapbuf_size3_mem_9_ccff_tail;
    wire [0:2]mux_tree_tapbuf_size5_0_sram;
    wire [0:2]mux_tree_tapbuf_size5_1_sram;
    wire [0:2]mux_tree_tapbuf_size5_2_sram;
    wire [0:2]mux_tree_tapbuf_size5_3_sram;
    wire [0:2]mux_tree_tapbuf_size5_4_sram;
    wire [0:2]mux_tree_tapbuf_size5_5_sram;
    wire mux_tree_tapbuf_size5_mem_0_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_1_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_2_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_3_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_4_ccff_tail;
    wire mux_tree_tapbuf_size5_mem_5_ccff_tail;

assign chany_bottom_out[28] = chanx_right_in[0];
assign chany_bottom_out[27] = chanx_right_in[1];
assign chany_bottom_out[26] = chanx_right_in[2];
assign chany_bottom_out[21] = chanx_right_in[7];
assign chany_bottom_out[20] = chanx_right_in[8];
assign chany_bottom_out[19] = chanx_right_in[9];
assign chany_bottom_out[18] = chanx_right_in[10];
assign chany_bottom_out[13] = chanx_right_in[15];
assign chany_bottom_out[12] = chanx_right_in[16];
assign chany_bottom_out[11] = chanx_right_in[17];
assign chany_bottom_out[10] = chanx_right_in[18];
assign chany_bottom_out[29] = chanx_right_in[29];
    mux_tree_tapbuf_size5 mux_right_track_0
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_, chany_bottom_in[28]}),
        .sram(mux_tree_tapbuf_size5_0_sram),
        .sram_inv(mux_right_track_0_undriven_sram_inv),
        .out(chanx_right_out[0])
    );
    mux_tree_tapbuf_size5 mux_right_track_2
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[27]}),
        .sram(mux_tree_tapbuf_size5_1_sram),
        .sram_inv(mux_right_track_2_undriven_sram_inv),
        .out(chanx_right_out[1])
    );
    mux_tree_tapbuf_size5 mux_right_track_4
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_, chany_bottom_in[26]}),
        .sram(mux_tree_tapbuf_size5_2_sram),
        .sram_inv(mux_right_track_4_undriven_sram_inv),
        .out(chanx_right_out[2])
    );
    mux_tree_tapbuf_size5 mux_right_track_6
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_, chany_bottom_in[25]}),
        .sram(mux_tree_tapbuf_size5_3_sram),
        .sram_inv(mux_right_track_6_undriven_sram_inv),
        .out(chanx_right_out[3])
    );
    mux_tree_tapbuf_size5 mux_right_track_8
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[24]}),
        .sram(mux_tree_tapbuf_size5_4_sram),
        .sram_inv(mux_right_track_8_undriven_sram_inv),
        .out(chanx_right_out[4])
    );
    mux_tree_tapbuf_size5 mux_right_track_10
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_, chany_bottom_in[23]}),
        .sram(mux_tree_tapbuf_size5_5_sram),
        .sram_inv(mux_right_track_10_undriven_sram_inv),
        .out(chanx_right_out[5])
    );
    mux_tree_tapbuf_size5_mem mem_right_track_0
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(ccff_head),
        .ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_0_sram)
    );
    mux_tree_tapbuf_size5_mem mem_right_track_2
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_1_sram)
    );
    mux_tree_tapbuf_size5_mem mem_right_track_4
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_2_sram)
    );
    mux_tree_tapbuf_size5_mem mem_right_track_6
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_3_sram)
    );
    mux_tree_tapbuf_size5_mem mem_right_track_8
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_4_sram)
    );
    mux_tree_tapbuf_size5_mem mem_right_track_10
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
        .mem_out(mux_tree_tapbuf_size5_5_sram)
    );
    mux_tree_tapbuf_size3 mux_right_track_12
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[22]}),
        .sram(mux_tree_tapbuf_size3_0_sram),
        .sram_inv(mux_right_track_12_undriven_sram_inv),
        .out(chanx_right_out[6])
    );
    mux_tree_tapbuf_size3 mux_right_track_14
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_, chany_bottom_in[21]}),
        .sram(mux_tree_tapbuf_size3_1_sram),
        .sram_inv(mux_right_track_14_undriven_sram_inv),
        .out(chanx_right_out[7])
    );
    mux_tree_tapbuf_size3 mux_right_track_16
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[20]}),
        .sram(mux_tree_tapbuf_size3_2_sram),
        .sram_inv(mux_right_track_16_undriven_sram_inv),
        .out(chanx_right_out[8])
    );
    mux_tree_tapbuf_size3 mux_right_track_28
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[14]}),
        .sram(mux_tree_tapbuf_size3_3_sram),
        .sram_inv(mux_right_track_28_undriven_sram_inv),
        .out(chanx_right_out[14])
    );
    mux_tree_tapbuf_size3 mux_right_track_30
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_, chany_bottom_in[13]}),
        .sram(mux_tree_tapbuf_size3_4_sram),
        .sram_inv(mux_right_track_30_undriven_sram_inv),
        .out(chanx_right_out[15])
    );
    mux_tree_tapbuf_size3 mux_right_track_32
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[12]}),
        .sram(mux_tree_tapbuf_size3_5_sram),
        .sram_inv(mux_right_track_32_undriven_sram_inv),
        .out(chanx_right_out[16])
    );
    mux_tree_tapbuf_size3 mux_right_track_34
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_, chany_bottom_in[11]}),
        .sram(mux_tree_tapbuf_size3_6_sram),
        .sram_inv(mux_right_track_34_undriven_sram_inv),
        .out(chanx_right_out[17])
    );
    mux_tree_tapbuf_size3 mux_right_track_44
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[6]}),
        .sram(mux_tree_tapbuf_size3_7_sram),
        .sram_inv(mux_right_track_44_undriven_sram_inv),
        .out(chanx_right_out[22])
    );
    mux_tree_tapbuf_size3 mux_right_track_46
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_, chany_bottom_in[5]}),
        .sram(mux_tree_tapbuf_size3_8_sram),
        .sram_inv(mux_right_track_46_undriven_sram_inv),
        .out(chanx_right_out[23])
    );
    mux_tree_tapbuf_size3 mux_right_track_48
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_, chany_bottom_in[4]}),
        .sram(mux_tree_tapbuf_size3_9_sram),
        .sram_inv(mux_right_track_48_undriven_sram_inv),
        .out(chanx_right_out[24])
    );
    mux_tree_tapbuf_size3 mux_right_track_58
    (
        .in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_, chany_bottom_in[29]}),
        .sram(mux_tree_tapbuf_size3_10_sram),
        .sram_inv(mux_right_track_58_undriven_sram_inv),
        .out(chanx_right_out[29])
    );
    mux_tree_tapbuf_size3 mux_bottom_track_1
    (
        .in({chanx_right_in[28], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size3_11_sram),
        .sram_inv(mux_bottom_track_1_undriven_sram_inv),
        .out(chany_bottom_out[0])
    );
    mux_tree_tapbuf_size3 mux_bottom_track_7
    (
        .in({chanx_right_in[25], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size3_12_sram),
        .sram_inv(mux_bottom_track_7_undriven_sram_inv),
        .out(chany_bottom_out[3])
    );
    mux_tree_tapbuf_size3_mem mem_right_track_12
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size3_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_0_sram)
    );
    mux_tree_tapbuf_size3_mem mem_right_track_14
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size3_mem_0_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size3_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_1_sram)
    );
    mux_tree_tapbuf_size3_mem mem_right_track_16
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size3_mem_1_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size3_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_2_sram)
    );
    mux_tree_tapbuf_size3_mem mem_right_track_28
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_4_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size3_mem_3_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_3_sram)
    );
    mux_tree_tapbuf_size3_mem mem_right_track_30
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size3_mem_3_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size3_mem_4_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_4_sram)
    );
    mux_tree_tapbuf_size3_mem mem_right_track_32
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size3_mem_4_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size3_mem_5_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_5_sram)
    );
    mux_tree_tapbuf_size3_mem mem_right_track_34
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size3_mem_5_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size3_mem_6_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_6_sram)
    );
    mux_tree_tapbuf_size3_mem mem_right_track_44
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_8_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size3_mem_7_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_7_sram)
    );
    mux_tree_tapbuf_size3_mem mem_right_track_46
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size3_mem_7_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size3_mem_8_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_8_sram)
    );
    mux_tree_tapbuf_size3_mem mem_right_track_48
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size3_mem_8_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size3_mem_9_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_9_sram)
    );
    mux_tree_tapbuf_size3_mem mem_right_track_58
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_12_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size3_mem_10_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_10_sram)
    );
    mux_tree_tapbuf_size3_mem mem_bottom_track_1
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size3_mem_10_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size3_mem_11_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_11_sram)
    );
    mux_tree_tapbuf_size3_mem mem_bottom_track_7
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_14_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size3_mem_12_ccff_tail),
        .mem_out(mux_tree_tapbuf_size3_12_sram)
    );
    mux_tree_tapbuf_size2 mux_right_track_18
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[19]}),
        .sram(mux_tree_tapbuf_size2_0_sram),
        .sram_inv(mux_right_track_18_undriven_sram_inv),
        .out(chanx_right_out[9])
    );
    mux_tree_tapbuf_size2 mux_right_track_20
    (
        .in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[18]}),
        .sram(mux_tree_tapbuf_size2_1_sram),
        .sram_inv(mux_right_track_20_undriven_sram_inv),
        .out(chanx_right_out[10])
    );
    mux_tree_tapbuf_size2 mux_right_track_22
    (
        .in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, chany_bottom_in[17]}),
        .sram(mux_tree_tapbuf_size2_2_sram),
        .sram_inv(mux_right_track_22_undriven_sram_inv),
        .out(chanx_right_out[11])
    );
    mux_tree_tapbuf_size2 mux_right_track_24
    (
        .in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[16]}),
        .sram(mux_tree_tapbuf_size2_3_sram),
        .sram_inv(mux_right_track_24_undriven_sram_inv),
        .out(chanx_right_out[12])
    );
    mux_tree_tapbuf_size2 mux_right_track_26
    (
        .in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, chany_bottom_in[15]}),
        .sram(mux_tree_tapbuf_size2_4_sram),
        .sram_inv(mux_right_track_26_undriven_sram_inv),
        .out(chanx_right_out[13])
    );
    mux_tree_tapbuf_size2 mux_right_track_36
    (
        .in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[10]}),
        .sram(mux_tree_tapbuf_size2_5_sram),
        .sram_inv(mux_right_track_36_undriven_sram_inv),
        .out(chanx_right_out[18])
    );
    mux_tree_tapbuf_size2 mux_right_track_38
    (
        .in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, chany_bottom_in[9]}),
        .sram(mux_tree_tapbuf_size2_6_sram),
        .sram_inv(mux_right_track_38_undriven_sram_inv),
        .out(chanx_right_out[19])
    );
    mux_tree_tapbuf_size2 mux_right_track_40
    (
        .in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[8]}),
        .sram(mux_tree_tapbuf_size2_7_sram),
        .sram_inv(mux_right_track_40_undriven_sram_inv),
        .out(chanx_right_out[20])
    );
    mux_tree_tapbuf_size2 mux_right_track_42
    (
        .in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, chany_bottom_in[7]}),
        .sram(mux_tree_tapbuf_size2_8_sram),
        .sram_inv(mux_right_track_42_undriven_sram_inv),
        .out(chanx_right_out[21])
    );
    mux_tree_tapbuf_size2 mux_right_track_50
    (
        .in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[3]}),
        .sram(mux_tree_tapbuf_size2_9_sram),
        .sram_inv(mux_right_track_50_undriven_sram_inv),
        .out(chanx_right_out[25])
    );
    mux_tree_tapbuf_size2 mux_right_track_52
    (
        .in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[2]}),
        .sram(mux_tree_tapbuf_size2_10_sram),
        .sram_inv(mux_right_track_52_undriven_sram_inv),
        .out(chanx_right_out[26])
    );
    mux_tree_tapbuf_size2 mux_right_track_54
    (
        .in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, chany_bottom_in[1]}),
        .sram(mux_tree_tapbuf_size2_11_sram),
        .sram_inv(mux_right_track_54_undriven_sram_inv),
        .out(chanx_right_out[27])
    );
    mux_tree_tapbuf_size2 mux_right_track_56
    (
        .in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[0]}),
        .sram(mux_tree_tapbuf_size2_12_sram),
        .sram_inv(mux_right_track_56_undriven_sram_inv),
        .out(chanx_right_out[28])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_3
    (
        .in({chanx_right_in[27], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_13_sram),
        .sram_inv(mux_bottom_track_3_undriven_sram_inv),
        .out(chany_bottom_out[1])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_5
    (
        .in({chanx_right_in[26], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_14_sram),
        .sram_inv(mux_bottom_track_5_undriven_sram_inv),
        .out(chany_bottom_out[2])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_9
    (
        .in({chanx_right_in[24], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_15_sram),
        .sram_inv(mux_bottom_track_9_undriven_sram_inv),
        .out(chany_bottom_out[4])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_11
    (
        .in({chanx_right_in[23], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_16_sram),
        .sram_inv(mux_bottom_track_11_undriven_sram_inv),
        .out(chany_bottom_out[5])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_13
    (
        .in({chanx_right_in[22], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_17_sram),
        .sram_inv(mux_bottom_track_13_undriven_sram_inv),
        .out(chany_bottom_out[6])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_15
    (
        .in({chanx_right_in[21], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_18_sram),
        .sram_inv(mux_bottom_track_15_undriven_sram_inv),
        .out(chany_bottom_out[7])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_17
    (
        .in({chanx_right_in[20], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_19_sram),
        .sram_inv(mux_bottom_track_17_undriven_sram_inv),
        .out(chany_bottom_out[8])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_19
    (
        .in({chanx_right_in[19], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_20_sram),
        .sram_inv(mux_bottom_track_19_undriven_sram_inv),
        .out(chany_bottom_out[9])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_29
    (
        .in({chanx_right_in[14], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_21_sram),
        .sram_inv(mux_bottom_track_29_undriven_sram_inv),
        .out(chany_bottom_out[14])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_31
    (
        .in({chanx_right_in[13], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_22_sram),
        .sram_inv(mux_bottom_track_31_undriven_sram_inv),
        .out(chany_bottom_out[15])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_33
    (
        .in({chanx_right_in[12], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_23_sram),
        .sram_inv(mux_bottom_track_33_undriven_sram_inv),
        .out(chany_bottom_out[16])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_35
    (
        .in({chanx_right_in[11], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_24_sram),
        .sram_inv(mux_bottom_track_35_undriven_sram_inv),
        .out(chany_bottom_out[17])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_45
    (
        .in({chanx_right_in[6], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_25_sram),
        .sram_inv(mux_bottom_track_45_undriven_sram_inv),
        .out(chany_bottom_out[22])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_47
    (
        .in({chanx_right_in[5], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_26_sram),
        .sram_inv(mux_bottom_track_47_undriven_sram_inv),
        .out(chany_bottom_out[23])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_49
    (
        .in({chanx_right_in[4], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_27_sram),
        .sram_inv(mux_bottom_track_49_undriven_sram_inv),
        .out(chany_bottom_out[24])
    );
    mux_tree_tapbuf_size2 mux_bottom_track_51
    (
        .in({chanx_right_in[3], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
        .sram(mux_tree_tapbuf_size2_28_sram),
        .sram_inv(mux_bottom_track_51_undriven_sram_inv),
        .out(chany_bottom_out[25])
    );
    mux_tree_tapbuf_size2_mem mem_right_track_18
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size3_mem_2_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_0_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_0_sram)
    );
    mux_tree_tapbuf_size2_mem mem_right_track_20
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_0_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_1_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_1_sram)
    );
    mux_tree_tapbuf_size2_mem mem_right_track_22
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_1_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_2_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_2_sram)
    );
    mux_tree_tapbuf_size2_mem mem_right_track_24
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_2_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_3_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_3_sram)
    );
    mux_tree_tapbuf_size2_mem mem_right_track_26
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_3_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_4_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_4_sram)
    );
    mux_tree_tapbuf_size2_mem mem_right_track_36
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size3_mem_6_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_5_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_5_sram)
    );
    mux_tree_tapbuf_size2_mem mem_right_track_38
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_5_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_6_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_6_sram)
    );
    mux_tree_tapbuf_size2_mem mem_right_track_40
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_6_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_7_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_7_sram)
    );
    mux_tree_tapbuf_size2_mem mem_right_track_42
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_7_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_8_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_8_sram)
    );
    mux_tree_tapbuf_size2_mem mem_right_track_50
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size3_mem_9_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_9_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_9_sram)
    );
    mux_tree_tapbuf_size2_mem mem_right_track_52
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_9_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_10_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_10_sram)
    );
    mux_tree_tapbuf_size2_mem mem_right_track_54
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_10_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_11_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_11_sram)
    );
    mux_tree_tapbuf_size2_mem mem_right_track_56
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_11_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_12_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_12_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_3
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size3_mem_11_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_13_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_13_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_5
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_13_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_14_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_14_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_9
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size3_mem_12_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_15_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_15_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_11
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_15_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_16_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_16_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_13
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_16_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_17_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_17_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_15
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_17_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_18_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_18_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_17
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_18_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_19_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_19_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_19
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_19_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_20_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_20_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_29
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_20_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_21_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_21_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_31
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_21_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_22_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_22_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_33
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_22_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_23_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_23_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_35
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_23_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_24_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_24_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_45
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_24_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_25_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_25_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_47
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_25_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_26_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_26_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_49
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_26_ccff_tail),
        .ccff_tail(mux_tree_tapbuf_size2_mem_27_ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_27_sram)
    );
    mux_tree_tapbuf_size2_mem mem_bottom_track_51
    (
        .prog_reset(prog_reset),
        .prog_clk(prog_clk),
        .ccff_head(mux_tree_tapbuf_size2_mem_27_ccff_tail),
        .ccff_tail(ccff_tail),
        .mem_out(mux_tree_tapbuf_size2_28_sram)
    );
endmodule

