VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER fieldpoly
  TYPE MASTERSLICE ;
END fieldpoly

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER diff
  TYPE MASTERSLICE ;
END diff

LAYER licon1
  TYPE MASTERSLICE ;
END licon1

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_0__0_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 113.16 BY 103.36 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 14.65 102 14.79 103.36 ;
    END
  END prog_clk[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.55 102 67.69 103.36 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.03 102 62.17 103.36 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.31 102 70.45 103.36 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 102 45.61 103.36 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.63 102 43.77 103.36 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.91 102 29.05 103.36 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.39 102 69.53 103.36 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.47 102 68.61 103.36 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.95 102 63.09 103.36 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 102 52.05 103.36 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 102 50.21 103.36 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.79 102 41.93 103.36 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.15 102 72.29 103.36 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.09 102 20.39 103.36 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.29 102 29.59 103.36 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.53 102 49.83 103.36 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.73 102 59.03 103.36 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 14.57 102 14.87 103.36 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.01 102 44.31 103.36 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 102 47.45 103.36 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.23 102 2.37 103.36 ;
    END
  END top_left_grid_pin_1_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 46.09 113.16 46.39 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 16.17 113.16 16.47 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 12.09 113.16 12.39 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 8.01 113.16 8.31 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 13.45 113.16 13.75 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 9.37 113.16 9.67 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 31.13 113.16 31.43 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 47.45 113.16 47.75 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 14.81 113.16 15.11 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 71.93 113.16 72.23 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 25.69 113.16 25.99 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 29.77 113.16 30.07 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 18.89 113.16 19.19 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 44.73 113.16 45.03 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 17.53 113.16 17.83 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 42.01 113.16 42.31 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 3.93 113.16 4.23 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 63.77 113.16 64.07 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 50.17 113.16 50.47 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 58.33 113.16 58.63 ;
    END
  END chanx_right_in[19]
  PIN right_top_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.87 74.8 110.01 76.16 ;
    END
  END right_top_grid_pin_42_[0]
  PIN right_top_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 99.13 84.64 99.43 ;
    END
  END right_top_grid_pin_43_[0]
  PIN right_top_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.79 74.8 110.93 76.16 ;
    END
  END right_top_grid_pin_44_[0]
  PIN right_top_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.95 74.8 109.09 76.16 ;
    END
  END right_top_grid_pin_45_[0]
  PIN right_top_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 91.65 84.64 91.95 ;
    END
  END right_top_grid_pin_46_[0]
  PIN right_top_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 90.29 84.64 90.59 ;
    END
  END right_top_grid_pin_47_[0]
  PIN right_top_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.11 74.8 107.25 76.16 ;
    END
  END right_top_grid_pin_48_[0]
  PIN right_top_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.03 74.8 108.17 76.16 ;
    END
  END right_top_grid_pin_49_[0]
  PIN right_bottom_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.87 0 110.01 1.36 ;
    END
  END right_bottom_grid_pin_1_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.79 0 110.93 1.36 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.71 102 42.85 103.36 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.69 102 25.83 103.36 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.23 102 71.37 103.36 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.15 102 49.29 103.36 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.27 102 36.41 103.36 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.55 102 44.69 103.36 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 5.37 102 5.67 103.36 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.85 102 69.15 103.36 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.93 102 22.23 103.36 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 9.05 102 9.35 103.36 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 102 46.53 103.36 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 102 51.13 103.36 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.29 102 7.43 103.36 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.77 102 24.07 103.36 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.21 102 7.51 103.36 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.85 102 46.15 103.36 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 102 48.37 103.36 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 102 52.97 103.36 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.69 102 47.99 103.36 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 25.61 102 25.91 103.36 ;
    END
  END chany_top_out[19]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 59.69 113.16 59.99 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 66.49 113.16 66.79 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 6.65 113.16 6.95 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 67.85 113.16 68.15 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 35.21 113.16 35.51 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 56.97 113.16 57.27 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 28.41 113.16 28.71 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 51.53 113.16 51.83 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 33.85 113.16 34.15 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 40.65 113.16 40.95 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 24.33 113.16 24.63 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 55.61 113.16 55.91 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 69.21 113.16 69.51 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 61.05 113.16 61.35 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 22.97 113.16 23.27 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 39.29 113.16 39.59 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 36.57 113.16 36.87 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 62.41 113.16 62.71 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 20.25 113.16 20.55 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 52.89 113.16 53.19 ;
    END
  END chanx_right_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 68.53 1.38 68.83 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 112.68 2.48 113.16 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 112.68 7.92 113.16 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 112.68 13.36 113.16 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 112.68 18.8 113.16 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 112.68 24.24 113.16 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 112.68 29.68 113.16 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 112.68 35.12 113.16 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 112.68 40.56 113.16 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 112.68 46 113.16 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 112.68 51.44 113.16 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 112.68 56.88 113.16 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 112.68 62.32 113.16 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 112.68 67.76 113.16 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 112.68 73.2 113.16 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 84.16 78.64 84.64 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 84.16 84.08 84.64 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 84.16 89.52 84.64 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 84.16 94.96 84.64 95.44 ;
        RECT 0 100.4 0.48 100.88 ;
        RECT 84.16 100.4 84.64 100.88 ;
      LAYER met4 ;
        RECT 12.58 0 13.18 0.6 ;
        RECT 42.02 0 42.62 0.6 ;
        RECT 71.46 0 72.06 0.6 ;
        RECT 106.42 0 107.02 0.6 ;
        RECT 106.42 75.56 107.02 76.16 ;
        RECT 12.58 102.76 13.18 103.36 ;
        RECT 42.02 102.76 42.62 103.36 ;
        RECT 71.46 102.76 72.06 103.36 ;
      LAYER met5 ;
        RECT 0 16.08 3.2 19.28 ;
        RECT 109.96 16.08 113.16 19.28 ;
        RECT 0 56.88 3.2 60.08 ;
        RECT 109.96 56.88 113.16 60.08 ;
        RECT 0 95.64 3.2 98.84 ;
        RECT 81.44 95.64 84.64 98.84 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 0 113.16 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 112.68 5.2 113.16 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 112.68 10.64 113.16 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 112.68 16.08 113.16 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 112.68 21.52 113.16 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 112.68 26.96 113.16 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 112.68 32.4 113.16 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 112.68 37.84 113.16 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 112.68 43.28 113.16 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 112.68 48.72 113.16 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 112.68 54.16 113.16 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 112.68 59.6 113.16 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 112.68 65.04 113.16 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 112.68 70.48 113.16 70.96 ;
        RECT 0 75.92 113.16 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 84.16 81.36 84.64 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 84.16 86.8 84.64 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 84.16 92.24 84.64 92.72 ;
        RECT 0 97.68 0.48 98.16 ;
        RECT 84.16 97.68 84.64 98.16 ;
        RECT 0 103.12 84.64 103.36 ;
      LAYER met4 ;
        RECT 27.3 0 27.9 0.6 ;
        RECT 56.74 0 57.34 0.6 ;
        RECT 27.3 102.76 27.9 103.36 ;
        RECT 56.74 102.76 57.34 103.36 ;
      LAYER met5 ;
        RECT 0 36.48 3.2 39.68 ;
        RECT 109.96 36.48 113.16 39.68 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 0 103.275 84.64 103.445 ;
      RECT 80.96 100.555 84.64 100.725 ;
      RECT 0 100.555 3.68 100.725 ;
      RECT 83.72 97.835 84.64 98.005 ;
      RECT 0 97.835 3.68 98.005 ;
      RECT 80.96 95.115 84.64 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 80.96 92.395 84.64 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 84.18 89.675 84.64 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 84.18 86.955 84.64 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 84.18 84.235 84.64 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 83.72 81.515 84.64 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 80.96 78.795 84.64 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 80.96 76.075 113.16 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 111.32 73.355 113.16 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 112.24 70.635 113.16 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 112.24 67.915 113.16 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 112.24 65.195 113.16 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 112.24 62.475 113.16 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 112.24 59.755 113.16 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 112.24 57.035 113.16 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 112.24 54.315 113.16 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 112.24 51.595 113.16 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 111.32 48.875 113.16 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 111.32 46.155 113.16 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 112.24 43.435 113.16 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 112.24 40.715 113.16 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 112.24 37.995 113.16 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 111.32 35.275 113.16 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 111.32 32.555 113.16 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 112.24 29.835 113.16 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 112.24 27.115 113.16 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 112.24 24.395 113.16 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 112.24 21.675 113.16 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 112.24 18.955 113.16 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 112.24 16.235 113.16 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 112.24 13.515 113.16 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 112.24 10.795 113.16 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 112.24 8.075 113.16 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 112.24 5.355 113.16 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 112.24 2.635 113.16 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 113.16 0.085 ;
    LAYER met2 ;
      RECT 56.9 103.175 57.18 103.545 ;
      RECT 27.46 103.175 27.74 103.545 ;
      RECT 45.87 101.5 46.13 101.82 ;
      RECT 56.9 -0.185 57.18 0.185 ;
      RECT 27.46 -0.185 27.74 0.185 ;
      POLYGON 84.36 103.08 84.36 75.88 106.83 75.88 106.83 74.52 107.53 74.52 107.53 75.88 107.75 75.88 107.75 74.52 108.45 74.52 108.45 75.88 108.67 75.88 108.67 74.52 109.37 74.52 109.37 75.88 109.59 75.88 109.59 74.52 110.29 74.52 110.29 75.88 110.51 75.88 110.51 74.52 111.21 74.52 111.21 75.88 112.88 75.88 112.88 0.28 111.21 0.28 111.21 1.64 110.51 1.64 110.51 0.28 110.29 0.28 110.29 1.64 109.59 1.64 109.59 0.28 0.28 0.28 0.28 103.08 1.95 103.08 1.95 101.72 2.65 101.72 2.65 103.08 7.01 103.08 7.01 101.72 7.71 101.72 7.71 103.08 14.37 103.08 14.37 101.72 15.07 101.72 15.07 103.08 25.41 103.08 25.41 101.72 26.11 101.72 26.11 103.08 28.63 103.08 28.63 101.72 29.33 101.72 29.33 103.08 35.99 103.08 35.99 101.72 36.69 101.72 36.69 103.08 41.51 103.08 41.51 101.72 42.21 101.72 42.21 103.08 42.43 103.08 42.43 101.72 43.13 101.72 43.13 103.08 43.35 103.08 43.35 101.72 44.05 101.72 44.05 103.08 44.27 103.08 44.27 101.72 44.97 101.72 44.97 103.08 45.19 103.08 45.19 101.72 45.89 101.72 45.89 103.08 46.11 103.08 46.11 101.72 46.81 101.72 46.81 103.08 47.03 103.08 47.03 101.72 47.73 101.72 47.73 103.08 47.95 103.08 47.95 101.72 48.65 101.72 48.65 103.08 48.87 103.08 48.87 101.72 49.57 101.72 49.57 103.08 49.79 103.08 49.79 101.72 50.49 101.72 50.49 103.08 50.71 103.08 50.71 101.72 51.41 101.72 51.41 103.08 51.63 103.08 51.63 101.72 52.33 101.72 52.33 103.08 52.55 103.08 52.55 101.72 53.25 101.72 53.25 103.08 61.75 103.08 61.75 101.72 62.45 101.72 62.45 103.08 62.67 103.08 62.67 101.72 63.37 101.72 63.37 103.08 67.27 103.08 67.27 101.72 67.97 101.72 67.97 103.08 68.19 103.08 68.19 101.72 68.89 101.72 68.89 103.08 69.11 103.08 69.11 101.72 69.81 101.72 69.81 103.08 70.03 103.08 70.03 101.72 70.73 101.72 70.73 103.08 70.95 103.08 70.95 101.72 71.65 101.72 71.65 103.08 71.87 103.08 71.87 101.72 72.57 101.72 72.57 103.08 ;
    LAYER met4 ;
      POLYGON 84.24 102.96 84.24 75.76 106.02 75.76 106.02 75.16 107.42 75.16 107.42 75.76 112.76 75.76 112.76 0.4 107.42 0.4 107.42 1 106.02 1 106.02 0.4 72.46 0.4 72.46 1 71.06 1 71.06 0.4 57.74 0.4 57.74 1 56.34 1 56.34 0.4 43.02 0.4 43.02 1 41.62 1 41.62 0.4 28.3 0.4 28.3 1 26.9 1 26.9 0.4 13.58 0.4 13.58 1 12.18 1 12.18 0.4 0.4 0.4 0.4 102.96 4.97 102.96 4.97 101.6 6.07 101.6 6.07 102.96 6.81 102.96 6.81 101.6 7.91 101.6 7.91 102.96 8.65 102.96 8.65 101.6 9.75 101.6 9.75 102.96 12.18 102.96 12.18 102.36 13.58 102.36 13.58 102.96 14.17 102.96 14.17 101.6 15.27 101.6 15.27 102.96 19.69 102.96 19.69 101.6 20.79 101.6 20.79 102.96 21.53 102.96 21.53 101.6 22.63 101.6 22.63 102.96 23.37 102.96 23.37 101.6 24.47 101.6 24.47 102.96 25.21 102.96 25.21 101.6 26.31 101.6 26.31 102.96 26.9 102.96 26.9 102.36 28.3 102.36 28.3 102.96 28.89 102.96 28.89 101.6 29.99 101.6 29.99 102.96 41.62 102.96 41.62 102.36 43.02 102.36 43.02 102.96 43.61 102.96 43.61 101.6 44.71 101.6 44.71 102.96 45.45 102.96 45.45 101.6 46.55 101.6 46.55 102.96 47.29 102.96 47.29 101.6 48.39 101.6 48.39 102.96 49.13 102.96 49.13 101.6 50.23 101.6 50.23 102.96 56.34 102.96 56.34 102.36 57.74 102.36 57.74 102.96 58.33 102.96 58.33 101.6 59.43 101.6 59.43 102.96 68.45 102.96 68.45 101.6 69.55 101.6 69.55 102.96 71.06 102.96 71.06 102.36 72.46 102.36 72.46 102.96 ;
    LAYER met3 ;
      POLYGON 57.205 103.525 57.205 103.52 57.42 103.52 57.42 103.2 57.205 103.2 57.205 103.195 56.875 103.195 56.875 103.2 56.66 103.2 56.66 103.52 56.875 103.52 56.875 103.525 ;
      POLYGON 27.765 103.525 27.765 103.52 27.98 103.52 27.98 103.2 27.765 103.2 27.765 103.195 27.435 103.195 27.435 103.2 27.22 103.2 27.22 103.52 27.435 103.52 27.435 103.525 ;
      POLYGON 111.485 37.565 111.485 37.235 111.155 37.235 111.155 37.25 106.11 37.25 106.11 37.55 111.155 37.55 111.155 37.565 ;
      POLYGON 57.205 0.165 57.205 0.16 57.42 0.16 57.42 -0.16 57.205 -0.16 57.205 -0.165 56.875 -0.165 56.875 -0.16 56.66 -0.16 56.66 0.16 56.875 0.16 56.875 0.165 ;
      POLYGON 27.765 0.165 27.765 0.16 27.98 0.16 27.98 -0.16 27.765 -0.16 27.765 -0.165 27.435 -0.165 27.435 -0.16 27.22 -0.16 27.22 0.16 27.435 0.16 27.435 0.165 ;
      POLYGON 84.24 102.96 84.24 99.83 82.86 99.83 82.86 98.73 84.24 98.73 84.24 92.35 82.86 92.35 82.86 91.25 84.24 91.25 84.24 90.99 82.86 90.99 82.86 89.89 84.24 89.89 84.24 75.76 112.76 75.76 112.76 72.63 111.38 72.63 111.38 71.53 112.76 71.53 112.76 69.91 111.38 69.91 111.38 68.81 112.76 68.81 112.76 68.55 111.38 68.55 111.38 67.45 112.76 67.45 112.76 67.19 111.38 67.19 111.38 66.09 112.76 66.09 112.76 64.47 111.38 64.47 111.38 63.37 112.76 63.37 112.76 63.11 111.38 63.11 111.38 62.01 112.76 62.01 112.76 61.75 111.38 61.75 111.38 60.65 112.76 60.65 112.76 60.39 111.38 60.39 111.38 59.29 112.76 59.29 112.76 59.03 111.38 59.03 111.38 57.93 112.76 57.93 112.76 57.67 111.38 57.67 111.38 56.57 112.76 56.57 112.76 56.31 111.38 56.31 111.38 55.21 112.76 55.21 112.76 53.59 111.38 53.59 111.38 52.49 112.76 52.49 112.76 52.23 111.38 52.23 111.38 51.13 112.76 51.13 112.76 50.87 111.38 50.87 111.38 49.77 112.76 49.77 112.76 48.15 111.38 48.15 111.38 47.05 112.76 47.05 112.76 46.79 111.38 46.79 111.38 45.69 112.76 45.69 112.76 45.43 111.38 45.43 111.38 44.33 112.76 44.33 112.76 42.71 111.38 42.71 111.38 41.61 112.76 41.61 112.76 41.35 111.38 41.35 111.38 40.25 112.76 40.25 112.76 39.99 111.38 39.99 111.38 38.89 112.76 38.89 112.76 37.27 111.38 37.27 111.38 36.17 112.76 36.17 112.76 35.91 111.38 35.91 111.38 34.81 112.76 34.81 112.76 34.55 111.38 34.55 111.38 33.45 112.76 33.45 112.76 31.83 111.38 31.83 111.38 30.73 112.76 30.73 112.76 30.47 111.38 30.47 111.38 29.37 112.76 29.37 112.76 29.11 111.38 29.11 111.38 28.01 112.76 28.01 112.76 26.39 111.38 26.39 111.38 25.29 112.76 25.29 112.76 25.03 111.38 25.03 111.38 23.93 112.76 23.93 112.76 23.67 111.38 23.67 111.38 22.57 112.76 22.57 112.76 20.95 111.38 20.95 111.38 19.85 112.76 19.85 112.76 19.59 111.38 19.59 111.38 18.49 112.76 18.49 112.76 18.23 111.38 18.23 111.38 17.13 112.76 17.13 112.76 16.87 111.38 16.87 111.38 15.77 112.76 15.77 112.76 15.51 111.38 15.51 111.38 14.41 112.76 14.41 112.76 14.15 111.38 14.15 111.38 13.05 112.76 13.05 112.76 12.79 111.38 12.79 111.38 11.69 112.76 11.69 112.76 10.07 111.38 10.07 111.38 8.97 112.76 8.97 112.76 8.71 111.38 8.71 111.38 7.61 112.76 7.61 112.76 7.35 111.38 7.35 111.38 6.25 112.76 6.25 112.76 4.63 111.38 4.63 111.38 3.53 112.76 3.53 112.76 0.4 0.4 0.4 0.4 68.13 1.78 68.13 1.78 69.23 0.4 69.23 0.4 102.96 ;
    LAYER met5 ;
      POLYGON 78.24 100.16 78.24 92.44 81.44 92.44 81.44 72.96 109.96 72.96 109.96 63.28 106.76 63.28 106.76 53.68 109.96 53.68 109.96 42.88 106.76 42.88 106.76 33.28 109.96 33.28 109.96 22.48 106.76 22.48 106.76 12.88 109.96 12.88 109.96 3.2 3.2 3.2 3.2 12.88 6.4 12.88 6.4 22.48 3.2 22.48 3.2 33.28 6.4 33.28 6.4 42.88 3.2 42.88 3.2 53.68 6.4 53.68 6.4 63.28 3.2 63.28 3.2 92.44 6.4 92.44 6.4 100.16 ;
    LAYER met1 ;
      POLYGON 84.36 102.84 84.36 101.16 83.88 101.16 83.88 100.12 84.36 100.12 84.36 98.44 83.88 98.44 83.88 97.4 84.36 97.4 84.36 95.72 83.88 95.72 83.88 94.68 84.36 94.68 84.36 93 83.88 93 83.88 91.96 84.36 91.96 84.36 90.28 83.88 90.28 83.88 89.24 84.36 89.24 84.36 87.56 83.88 87.56 83.88 86.52 84.36 86.52 84.36 84.84 83.88 84.84 83.88 83.8 84.36 83.8 84.36 82.12 83.88 82.12 83.88 81.08 84.36 81.08 84.36 79.4 83.88 79.4 83.88 78.36 84.36 78.36 84.36 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 0.76 97.4 0.76 98.44 0.28 98.44 0.28 100.12 0.76 100.12 0.76 101.16 0.28 101.16 0.28 102.84 ;
      POLYGON 112.88 75.64 112.88 73.96 112.4 73.96 112.4 72.92 112.88 72.92 112.88 71.24 112.4 71.24 112.4 70.2 112.88 70.2 112.88 68.52 112.4 68.52 112.4 67.48 112.88 67.48 112.88 65.8 112.4 65.8 112.4 64.76 112.88 64.76 112.88 63.08 112.4 63.08 112.4 62.04 112.88 62.04 112.88 60.36 112.4 60.36 112.4 59.32 112.88 59.32 112.88 57.64 112.4 57.64 112.4 56.6 112.88 56.6 112.88 54.92 112.4 54.92 112.4 53.88 112.88 53.88 112.88 52.2 112.4 52.2 112.4 51.16 112.88 51.16 112.88 49.48 112.4 49.48 112.4 48.44 112.88 48.44 112.88 46.76 112.4 46.76 112.4 45.72 112.88 45.72 112.88 44.04 112.4 44.04 112.4 43 112.88 43 112.88 41.32 112.4 41.32 112.4 40.28 112.88 40.28 112.88 38.6 112.4 38.6 112.4 37.56 112.88 37.56 112.88 35.88 112.4 35.88 112.4 34.84 112.88 34.84 112.88 33.16 112.4 33.16 112.4 32.12 112.88 32.12 112.88 30.44 112.4 30.44 112.4 29.4 112.88 29.4 112.88 27.72 112.4 27.72 112.4 26.68 112.88 26.68 112.88 25 112.4 25 112.4 23.96 112.88 23.96 112.88 22.28 112.4 22.28 112.4 21.24 112.88 21.24 112.88 19.56 112.4 19.56 112.4 18.52 112.88 18.52 112.88 16.84 112.4 16.84 112.4 15.8 112.88 15.8 112.88 14.12 112.4 14.12 112.4 13.08 112.88 13.08 112.88 11.4 112.4 11.4 112.4 10.36 112.88 10.36 112.88 8.68 112.4 8.68 112.4 7.64 112.88 7.64 112.88 5.96 112.4 5.96 112.4 4.92 112.88 4.92 112.88 3.24 112.4 3.24 112.4 2.2 112.88 2.2 112.88 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 ;
    LAYER li1 ;
      POLYGON 84.3 103.02 84.3 75.82 112.82 75.82 112.82 0.34 0.34 0.34 0.34 103.02 ;
    LAYER mcon ;
      RECT 84.325 103.275 84.495 103.445 ;
      RECT 83.865 103.275 84.035 103.445 ;
      RECT 83.405 103.275 83.575 103.445 ;
      RECT 82.945 103.275 83.115 103.445 ;
      RECT 82.485 103.275 82.655 103.445 ;
      RECT 82.025 103.275 82.195 103.445 ;
      RECT 81.565 103.275 81.735 103.445 ;
      RECT 81.105 103.275 81.275 103.445 ;
      RECT 80.645 103.275 80.815 103.445 ;
      RECT 80.185 103.275 80.355 103.445 ;
      RECT 79.725 103.275 79.895 103.445 ;
      RECT 79.265 103.275 79.435 103.445 ;
      RECT 78.805 103.275 78.975 103.445 ;
      RECT 78.345 103.275 78.515 103.445 ;
      RECT 77.885 103.275 78.055 103.445 ;
      RECT 77.425 103.275 77.595 103.445 ;
      RECT 76.965 103.275 77.135 103.445 ;
      RECT 76.505 103.275 76.675 103.445 ;
      RECT 76.045 103.275 76.215 103.445 ;
      RECT 75.585 103.275 75.755 103.445 ;
      RECT 75.125 103.275 75.295 103.445 ;
      RECT 74.665 103.275 74.835 103.445 ;
      RECT 74.205 103.275 74.375 103.445 ;
      RECT 73.745 103.275 73.915 103.445 ;
      RECT 73.285 103.275 73.455 103.445 ;
      RECT 72.825 103.275 72.995 103.445 ;
      RECT 72.365 103.275 72.535 103.445 ;
      RECT 71.905 103.275 72.075 103.445 ;
      RECT 71.445 103.275 71.615 103.445 ;
      RECT 70.985 103.275 71.155 103.445 ;
      RECT 70.525 103.275 70.695 103.445 ;
      RECT 70.065 103.275 70.235 103.445 ;
      RECT 69.605 103.275 69.775 103.445 ;
      RECT 69.145 103.275 69.315 103.445 ;
      RECT 68.685 103.275 68.855 103.445 ;
      RECT 68.225 103.275 68.395 103.445 ;
      RECT 67.765 103.275 67.935 103.445 ;
      RECT 67.305 103.275 67.475 103.445 ;
      RECT 66.845 103.275 67.015 103.445 ;
      RECT 66.385 103.275 66.555 103.445 ;
      RECT 65.925 103.275 66.095 103.445 ;
      RECT 65.465 103.275 65.635 103.445 ;
      RECT 65.005 103.275 65.175 103.445 ;
      RECT 64.545 103.275 64.715 103.445 ;
      RECT 64.085 103.275 64.255 103.445 ;
      RECT 63.625 103.275 63.795 103.445 ;
      RECT 63.165 103.275 63.335 103.445 ;
      RECT 62.705 103.275 62.875 103.445 ;
      RECT 62.245 103.275 62.415 103.445 ;
      RECT 61.785 103.275 61.955 103.445 ;
      RECT 61.325 103.275 61.495 103.445 ;
      RECT 60.865 103.275 61.035 103.445 ;
      RECT 60.405 103.275 60.575 103.445 ;
      RECT 59.945 103.275 60.115 103.445 ;
      RECT 59.485 103.275 59.655 103.445 ;
      RECT 59.025 103.275 59.195 103.445 ;
      RECT 58.565 103.275 58.735 103.445 ;
      RECT 58.105 103.275 58.275 103.445 ;
      RECT 57.645 103.275 57.815 103.445 ;
      RECT 57.185 103.275 57.355 103.445 ;
      RECT 56.725 103.275 56.895 103.445 ;
      RECT 56.265 103.275 56.435 103.445 ;
      RECT 55.805 103.275 55.975 103.445 ;
      RECT 55.345 103.275 55.515 103.445 ;
      RECT 54.885 103.275 55.055 103.445 ;
      RECT 54.425 103.275 54.595 103.445 ;
      RECT 53.965 103.275 54.135 103.445 ;
      RECT 53.505 103.275 53.675 103.445 ;
      RECT 53.045 103.275 53.215 103.445 ;
      RECT 52.585 103.275 52.755 103.445 ;
      RECT 52.125 103.275 52.295 103.445 ;
      RECT 51.665 103.275 51.835 103.445 ;
      RECT 51.205 103.275 51.375 103.445 ;
      RECT 50.745 103.275 50.915 103.445 ;
      RECT 50.285 103.275 50.455 103.445 ;
      RECT 49.825 103.275 49.995 103.445 ;
      RECT 49.365 103.275 49.535 103.445 ;
      RECT 48.905 103.275 49.075 103.445 ;
      RECT 48.445 103.275 48.615 103.445 ;
      RECT 47.985 103.275 48.155 103.445 ;
      RECT 47.525 103.275 47.695 103.445 ;
      RECT 47.065 103.275 47.235 103.445 ;
      RECT 46.605 103.275 46.775 103.445 ;
      RECT 46.145 103.275 46.315 103.445 ;
      RECT 45.685 103.275 45.855 103.445 ;
      RECT 45.225 103.275 45.395 103.445 ;
      RECT 44.765 103.275 44.935 103.445 ;
      RECT 44.305 103.275 44.475 103.445 ;
      RECT 43.845 103.275 44.015 103.445 ;
      RECT 43.385 103.275 43.555 103.445 ;
      RECT 42.925 103.275 43.095 103.445 ;
      RECT 42.465 103.275 42.635 103.445 ;
      RECT 42.005 103.275 42.175 103.445 ;
      RECT 41.545 103.275 41.715 103.445 ;
      RECT 41.085 103.275 41.255 103.445 ;
      RECT 40.625 103.275 40.795 103.445 ;
      RECT 40.165 103.275 40.335 103.445 ;
      RECT 39.705 103.275 39.875 103.445 ;
      RECT 39.245 103.275 39.415 103.445 ;
      RECT 38.785 103.275 38.955 103.445 ;
      RECT 38.325 103.275 38.495 103.445 ;
      RECT 37.865 103.275 38.035 103.445 ;
      RECT 37.405 103.275 37.575 103.445 ;
      RECT 36.945 103.275 37.115 103.445 ;
      RECT 36.485 103.275 36.655 103.445 ;
      RECT 36.025 103.275 36.195 103.445 ;
      RECT 35.565 103.275 35.735 103.445 ;
      RECT 35.105 103.275 35.275 103.445 ;
      RECT 34.645 103.275 34.815 103.445 ;
      RECT 34.185 103.275 34.355 103.445 ;
      RECT 33.725 103.275 33.895 103.445 ;
      RECT 33.265 103.275 33.435 103.445 ;
      RECT 32.805 103.275 32.975 103.445 ;
      RECT 32.345 103.275 32.515 103.445 ;
      RECT 31.885 103.275 32.055 103.445 ;
      RECT 31.425 103.275 31.595 103.445 ;
      RECT 30.965 103.275 31.135 103.445 ;
      RECT 30.505 103.275 30.675 103.445 ;
      RECT 30.045 103.275 30.215 103.445 ;
      RECT 29.585 103.275 29.755 103.445 ;
      RECT 29.125 103.275 29.295 103.445 ;
      RECT 28.665 103.275 28.835 103.445 ;
      RECT 28.205 103.275 28.375 103.445 ;
      RECT 27.745 103.275 27.915 103.445 ;
      RECT 27.285 103.275 27.455 103.445 ;
      RECT 26.825 103.275 26.995 103.445 ;
      RECT 26.365 103.275 26.535 103.445 ;
      RECT 25.905 103.275 26.075 103.445 ;
      RECT 25.445 103.275 25.615 103.445 ;
      RECT 24.985 103.275 25.155 103.445 ;
      RECT 24.525 103.275 24.695 103.445 ;
      RECT 24.065 103.275 24.235 103.445 ;
      RECT 23.605 103.275 23.775 103.445 ;
      RECT 23.145 103.275 23.315 103.445 ;
      RECT 22.685 103.275 22.855 103.445 ;
      RECT 22.225 103.275 22.395 103.445 ;
      RECT 21.765 103.275 21.935 103.445 ;
      RECT 21.305 103.275 21.475 103.445 ;
      RECT 20.845 103.275 21.015 103.445 ;
      RECT 20.385 103.275 20.555 103.445 ;
      RECT 19.925 103.275 20.095 103.445 ;
      RECT 19.465 103.275 19.635 103.445 ;
      RECT 19.005 103.275 19.175 103.445 ;
      RECT 18.545 103.275 18.715 103.445 ;
      RECT 18.085 103.275 18.255 103.445 ;
      RECT 17.625 103.275 17.795 103.445 ;
      RECT 17.165 103.275 17.335 103.445 ;
      RECT 16.705 103.275 16.875 103.445 ;
      RECT 16.245 103.275 16.415 103.445 ;
      RECT 15.785 103.275 15.955 103.445 ;
      RECT 15.325 103.275 15.495 103.445 ;
      RECT 14.865 103.275 15.035 103.445 ;
      RECT 14.405 103.275 14.575 103.445 ;
      RECT 13.945 103.275 14.115 103.445 ;
      RECT 13.485 103.275 13.655 103.445 ;
      RECT 13.025 103.275 13.195 103.445 ;
      RECT 12.565 103.275 12.735 103.445 ;
      RECT 12.105 103.275 12.275 103.445 ;
      RECT 11.645 103.275 11.815 103.445 ;
      RECT 11.185 103.275 11.355 103.445 ;
      RECT 10.725 103.275 10.895 103.445 ;
      RECT 10.265 103.275 10.435 103.445 ;
      RECT 9.805 103.275 9.975 103.445 ;
      RECT 9.345 103.275 9.515 103.445 ;
      RECT 8.885 103.275 9.055 103.445 ;
      RECT 8.425 103.275 8.595 103.445 ;
      RECT 7.965 103.275 8.135 103.445 ;
      RECT 7.505 103.275 7.675 103.445 ;
      RECT 7.045 103.275 7.215 103.445 ;
      RECT 6.585 103.275 6.755 103.445 ;
      RECT 6.125 103.275 6.295 103.445 ;
      RECT 5.665 103.275 5.835 103.445 ;
      RECT 5.205 103.275 5.375 103.445 ;
      RECT 4.745 103.275 4.915 103.445 ;
      RECT 4.285 103.275 4.455 103.445 ;
      RECT 3.825 103.275 3.995 103.445 ;
      RECT 3.365 103.275 3.535 103.445 ;
      RECT 2.905 103.275 3.075 103.445 ;
      RECT 2.445 103.275 2.615 103.445 ;
      RECT 1.985 103.275 2.155 103.445 ;
      RECT 1.525 103.275 1.695 103.445 ;
      RECT 1.065 103.275 1.235 103.445 ;
      RECT 0.605 103.275 0.775 103.445 ;
      RECT 0.145 103.275 0.315 103.445 ;
      RECT 84.325 100.555 84.495 100.725 ;
      RECT 83.865 100.555 84.035 100.725 ;
      RECT 0.605 100.555 0.775 100.725 ;
      RECT 0.145 100.555 0.315 100.725 ;
      RECT 84.325 97.835 84.495 98.005 ;
      RECT 83.865 97.835 84.035 98.005 ;
      RECT 0.605 97.835 0.775 98.005 ;
      RECT 0.145 97.835 0.315 98.005 ;
      RECT 84.325 95.115 84.495 95.285 ;
      RECT 83.865 95.115 84.035 95.285 ;
      RECT 0.605 95.115 0.775 95.285 ;
      RECT 0.145 95.115 0.315 95.285 ;
      RECT 84.325 92.395 84.495 92.565 ;
      RECT 83.865 92.395 84.035 92.565 ;
      RECT 0.605 92.395 0.775 92.565 ;
      RECT 0.145 92.395 0.315 92.565 ;
      RECT 84.325 89.675 84.495 89.845 ;
      RECT 83.865 89.675 84.035 89.845 ;
      RECT 0.605 89.675 0.775 89.845 ;
      RECT 0.145 89.675 0.315 89.845 ;
      RECT 84.325 86.955 84.495 87.125 ;
      RECT 83.865 86.955 84.035 87.125 ;
      RECT 0.605 86.955 0.775 87.125 ;
      RECT 0.145 86.955 0.315 87.125 ;
      RECT 84.325 84.235 84.495 84.405 ;
      RECT 83.865 84.235 84.035 84.405 ;
      RECT 0.605 84.235 0.775 84.405 ;
      RECT 0.145 84.235 0.315 84.405 ;
      RECT 84.325 81.515 84.495 81.685 ;
      RECT 83.865 81.515 84.035 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 84.325 78.795 84.495 78.965 ;
      RECT 83.865 78.795 84.035 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 112.845 76.075 113.015 76.245 ;
      RECT 112.385 76.075 112.555 76.245 ;
      RECT 111.925 76.075 112.095 76.245 ;
      RECT 111.465 76.075 111.635 76.245 ;
      RECT 111.005 76.075 111.175 76.245 ;
      RECT 110.545 76.075 110.715 76.245 ;
      RECT 110.085 76.075 110.255 76.245 ;
      RECT 109.625 76.075 109.795 76.245 ;
      RECT 109.165 76.075 109.335 76.245 ;
      RECT 108.705 76.075 108.875 76.245 ;
      RECT 108.245 76.075 108.415 76.245 ;
      RECT 107.785 76.075 107.955 76.245 ;
      RECT 107.325 76.075 107.495 76.245 ;
      RECT 106.865 76.075 107.035 76.245 ;
      RECT 106.405 76.075 106.575 76.245 ;
      RECT 105.945 76.075 106.115 76.245 ;
      RECT 105.485 76.075 105.655 76.245 ;
      RECT 105.025 76.075 105.195 76.245 ;
      RECT 104.565 76.075 104.735 76.245 ;
      RECT 104.105 76.075 104.275 76.245 ;
      RECT 103.645 76.075 103.815 76.245 ;
      RECT 103.185 76.075 103.355 76.245 ;
      RECT 102.725 76.075 102.895 76.245 ;
      RECT 102.265 76.075 102.435 76.245 ;
      RECT 101.805 76.075 101.975 76.245 ;
      RECT 101.345 76.075 101.515 76.245 ;
      RECT 100.885 76.075 101.055 76.245 ;
      RECT 100.425 76.075 100.595 76.245 ;
      RECT 99.965 76.075 100.135 76.245 ;
      RECT 99.505 76.075 99.675 76.245 ;
      RECT 99.045 76.075 99.215 76.245 ;
      RECT 98.585 76.075 98.755 76.245 ;
      RECT 98.125 76.075 98.295 76.245 ;
      RECT 97.665 76.075 97.835 76.245 ;
      RECT 97.205 76.075 97.375 76.245 ;
      RECT 96.745 76.075 96.915 76.245 ;
      RECT 96.285 76.075 96.455 76.245 ;
      RECT 95.825 76.075 95.995 76.245 ;
      RECT 95.365 76.075 95.535 76.245 ;
      RECT 94.905 76.075 95.075 76.245 ;
      RECT 94.445 76.075 94.615 76.245 ;
      RECT 93.985 76.075 94.155 76.245 ;
      RECT 93.525 76.075 93.695 76.245 ;
      RECT 93.065 76.075 93.235 76.245 ;
      RECT 92.605 76.075 92.775 76.245 ;
      RECT 92.145 76.075 92.315 76.245 ;
      RECT 91.685 76.075 91.855 76.245 ;
      RECT 91.225 76.075 91.395 76.245 ;
      RECT 90.765 76.075 90.935 76.245 ;
      RECT 90.305 76.075 90.475 76.245 ;
      RECT 89.845 76.075 90.015 76.245 ;
      RECT 89.385 76.075 89.555 76.245 ;
      RECT 88.925 76.075 89.095 76.245 ;
      RECT 88.465 76.075 88.635 76.245 ;
      RECT 88.005 76.075 88.175 76.245 ;
      RECT 87.545 76.075 87.715 76.245 ;
      RECT 87.085 76.075 87.255 76.245 ;
      RECT 86.625 76.075 86.795 76.245 ;
      RECT 86.165 76.075 86.335 76.245 ;
      RECT 85.705 76.075 85.875 76.245 ;
      RECT 85.245 76.075 85.415 76.245 ;
      RECT 84.785 76.075 84.955 76.245 ;
      RECT 84.325 76.075 84.495 76.245 ;
      RECT 83.865 76.075 84.035 76.245 ;
      RECT 83.405 76.075 83.575 76.245 ;
      RECT 82.945 76.075 83.115 76.245 ;
      RECT 82.485 76.075 82.655 76.245 ;
      RECT 82.025 76.075 82.195 76.245 ;
      RECT 81.565 76.075 81.735 76.245 ;
      RECT 81.105 76.075 81.275 76.245 ;
      RECT 80.645 76.075 80.815 76.245 ;
      RECT 80.185 76.075 80.355 76.245 ;
      RECT 79.725 76.075 79.895 76.245 ;
      RECT 79.265 76.075 79.435 76.245 ;
      RECT 78.805 76.075 78.975 76.245 ;
      RECT 78.345 76.075 78.515 76.245 ;
      RECT 77.885 76.075 78.055 76.245 ;
      RECT 77.425 76.075 77.595 76.245 ;
      RECT 76.965 76.075 77.135 76.245 ;
      RECT 76.505 76.075 76.675 76.245 ;
      RECT 76.045 76.075 76.215 76.245 ;
      RECT 75.585 76.075 75.755 76.245 ;
      RECT 75.125 76.075 75.295 76.245 ;
      RECT 74.665 76.075 74.835 76.245 ;
      RECT 74.205 76.075 74.375 76.245 ;
      RECT 73.745 76.075 73.915 76.245 ;
      RECT 73.285 76.075 73.455 76.245 ;
      RECT 72.825 76.075 72.995 76.245 ;
      RECT 72.365 76.075 72.535 76.245 ;
      RECT 71.905 76.075 72.075 76.245 ;
      RECT 71.445 76.075 71.615 76.245 ;
      RECT 70.985 76.075 71.155 76.245 ;
      RECT 70.525 76.075 70.695 76.245 ;
      RECT 70.065 76.075 70.235 76.245 ;
      RECT 69.605 76.075 69.775 76.245 ;
      RECT 69.145 76.075 69.315 76.245 ;
      RECT 68.685 76.075 68.855 76.245 ;
      RECT 68.225 76.075 68.395 76.245 ;
      RECT 67.765 76.075 67.935 76.245 ;
      RECT 67.305 76.075 67.475 76.245 ;
      RECT 66.845 76.075 67.015 76.245 ;
      RECT 66.385 76.075 66.555 76.245 ;
      RECT 65.925 76.075 66.095 76.245 ;
      RECT 65.465 76.075 65.635 76.245 ;
      RECT 65.005 76.075 65.175 76.245 ;
      RECT 64.545 76.075 64.715 76.245 ;
      RECT 64.085 76.075 64.255 76.245 ;
      RECT 63.625 76.075 63.795 76.245 ;
      RECT 63.165 76.075 63.335 76.245 ;
      RECT 62.705 76.075 62.875 76.245 ;
      RECT 62.245 76.075 62.415 76.245 ;
      RECT 61.785 76.075 61.955 76.245 ;
      RECT 61.325 76.075 61.495 76.245 ;
      RECT 60.865 76.075 61.035 76.245 ;
      RECT 60.405 76.075 60.575 76.245 ;
      RECT 59.945 76.075 60.115 76.245 ;
      RECT 59.485 76.075 59.655 76.245 ;
      RECT 59.025 76.075 59.195 76.245 ;
      RECT 58.565 76.075 58.735 76.245 ;
      RECT 58.105 76.075 58.275 76.245 ;
      RECT 57.645 76.075 57.815 76.245 ;
      RECT 57.185 76.075 57.355 76.245 ;
      RECT 56.725 76.075 56.895 76.245 ;
      RECT 56.265 76.075 56.435 76.245 ;
      RECT 55.805 76.075 55.975 76.245 ;
      RECT 55.345 76.075 55.515 76.245 ;
      RECT 54.885 76.075 55.055 76.245 ;
      RECT 54.425 76.075 54.595 76.245 ;
      RECT 53.965 76.075 54.135 76.245 ;
      RECT 53.505 76.075 53.675 76.245 ;
      RECT 53.045 76.075 53.215 76.245 ;
      RECT 52.585 76.075 52.755 76.245 ;
      RECT 52.125 76.075 52.295 76.245 ;
      RECT 51.665 76.075 51.835 76.245 ;
      RECT 51.205 76.075 51.375 76.245 ;
      RECT 50.745 76.075 50.915 76.245 ;
      RECT 50.285 76.075 50.455 76.245 ;
      RECT 49.825 76.075 49.995 76.245 ;
      RECT 49.365 76.075 49.535 76.245 ;
      RECT 48.905 76.075 49.075 76.245 ;
      RECT 48.445 76.075 48.615 76.245 ;
      RECT 47.985 76.075 48.155 76.245 ;
      RECT 47.525 76.075 47.695 76.245 ;
      RECT 47.065 76.075 47.235 76.245 ;
      RECT 46.605 76.075 46.775 76.245 ;
      RECT 46.145 76.075 46.315 76.245 ;
      RECT 45.685 76.075 45.855 76.245 ;
      RECT 45.225 76.075 45.395 76.245 ;
      RECT 44.765 76.075 44.935 76.245 ;
      RECT 44.305 76.075 44.475 76.245 ;
      RECT 43.845 76.075 44.015 76.245 ;
      RECT 43.385 76.075 43.555 76.245 ;
      RECT 42.925 76.075 43.095 76.245 ;
      RECT 42.465 76.075 42.635 76.245 ;
      RECT 42.005 76.075 42.175 76.245 ;
      RECT 41.545 76.075 41.715 76.245 ;
      RECT 41.085 76.075 41.255 76.245 ;
      RECT 40.625 76.075 40.795 76.245 ;
      RECT 40.165 76.075 40.335 76.245 ;
      RECT 39.705 76.075 39.875 76.245 ;
      RECT 39.245 76.075 39.415 76.245 ;
      RECT 38.785 76.075 38.955 76.245 ;
      RECT 38.325 76.075 38.495 76.245 ;
      RECT 37.865 76.075 38.035 76.245 ;
      RECT 37.405 76.075 37.575 76.245 ;
      RECT 36.945 76.075 37.115 76.245 ;
      RECT 36.485 76.075 36.655 76.245 ;
      RECT 36.025 76.075 36.195 76.245 ;
      RECT 35.565 76.075 35.735 76.245 ;
      RECT 35.105 76.075 35.275 76.245 ;
      RECT 34.645 76.075 34.815 76.245 ;
      RECT 34.185 76.075 34.355 76.245 ;
      RECT 33.725 76.075 33.895 76.245 ;
      RECT 33.265 76.075 33.435 76.245 ;
      RECT 32.805 76.075 32.975 76.245 ;
      RECT 32.345 76.075 32.515 76.245 ;
      RECT 31.885 76.075 32.055 76.245 ;
      RECT 31.425 76.075 31.595 76.245 ;
      RECT 30.965 76.075 31.135 76.245 ;
      RECT 30.505 76.075 30.675 76.245 ;
      RECT 30.045 76.075 30.215 76.245 ;
      RECT 29.585 76.075 29.755 76.245 ;
      RECT 29.125 76.075 29.295 76.245 ;
      RECT 28.665 76.075 28.835 76.245 ;
      RECT 28.205 76.075 28.375 76.245 ;
      RECT 27.745 76.075 27.915 76.245 ;
      RECT 27.285 76.075 27.455 76.245 ;
      RECT 26.825 76.075 26.995 76.245 ;
      RECT 26.365 76.075 26.535 76.245 ;
      RECT 25.905 76.075 26.075 76.245 ;
      RECT 25.445 76.075 25.615 76.245 ;
      RECT 24.985 76.075 25.155 76.245 ;
      RECT 24.525 76.075 24.695 76.245 ;
      RECT 24.065 76.075 24.235 76.245 ;
      RECT 23.605 76.075 23.775 76.245 ;
      RECT 23.145 76.075 23.315 76.245 ;
      RECT 22.685 76.075 22.855 76.245 ;
      RECT 22.225 76.075 22.395 76.245 ;
      RECT 21.765 76.075 21.935 76.245 ;
      RECT 21.305 76.075 21.475 76.245 ;
      RECT 20.845 76.075 21.015 76.245 ;
      RECT 20.385 76.075 20.555 76.245 ;
      RECT 19.925 76.075 20.095 76.245 ;
      RECT 19.465 76.075 19.635 76.245 ;
      RECT 19.005 76.075 19.175 76.245 ;
      RECT 18.545 76.075 18.715 76.245 ;
      RECT 18.085 76.075 18.255 76.245 ;
      RECT 17.625 76.075 17.795 76.245 ;
      RECT 17.165 76.075 17.335 76.245 ;
      RECT 16.705 76.075 16.875 76.245 ;
      RECT 16.245 76.075 16.415 76.245 ;
      RECT 15.785 76.075 15.955 76.245 ;
      RECT 15.325 76.075 15.495 76.245 ;
      RECT 14.865 76.075 15.035 76.245 ;
      RECT 14.405 76.075 14.575 76.245 ;
      RECT 13.945 76.075 14.115 76.245 ;
      RECT 13.485 76.075 13.655 76.245 ;
      RECT 13.025 76.075 13.195 76.245 ;
      RECT 12.565 76.075 12.735 76.245 ;
      RECT 12.105 76.075 12.275 76.245 ;
      RECT 11.645 76.075 11.815 76.245 ;
      RECT 11.185 76.075 11.355 76.245 ;
      RECT 10.725 76.075 10.895 76.245 ;
      RECT 10.265 76.075 10.435 76.245 ;
      RECT 9.805 76.075 9.975 76.245 ;
      RECT 9.345 76.075 9.515 76.245 ;
      RECT 8.885 76.075 9.055 76.245 ;
      RECT 8.425 76.075 8.595 76.245 ;
      RECT 7.965 76.075 8.135 76.245 ;
      RECT 7.505 76.075 7.675 76.245 ;
      RECT 7.045 76.075 7.215 76.245 ;
      RECT 6.585 76.075 6.755 76.245 ;
      RECT 6.125 76.075 6.295 76.245 ;
      RECT 5.665 76.075 5.835 76.245 ;
      RECT 5.205 76.075 5.375 76.245 ;
      RECT 4.745 76.075 4.915 76.245 ;
      RECT 4.285 76.075 4.455 76.245 ;
      RECT 3.825 76.075 3.995 76.245 ;
      RECT 3.365 76.075 3.535 76.245 ;
      RECT 2.905 76.075 3.075 76.245 ;
      RECT 2.445 76.075 2.615 76.245 ;
      RECT 1.985 76.075 2.155 76.245 ;
      RECT 1.525 76.075 1.695 76.245 ;
      RECT 1.065 76.075 1.235 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 112.845 73.355 113.015 73.525 ;
      RECT 112.385 73.355 112.555 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 112.845 70.635 113.015 70.805 ;
      RECT 112.385 70.635 112.555 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 112.845 67.915 113.015 68.085 ;
      RECT 112.385 67.915 112.555 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 112.845 65.195 113.015 65.365 ;
      RECT 112.385 65.195 112.555 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 112.845 62.475 113.015 62.645 ;
      RECT 112.385 62.475 112.555 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 112.845 59.755 113.015 59.925 ;
      RECT 112.385 59.755 112.555 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 112.845 57.035 113.015 57.205 ;
      RECT 112.385 57.035 112.555 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 112.845 54.315 113.015 54.485 ;
      RECT 112.385 54.315 112.555 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 112.845 51.595 113.015 51.765 ;
      RECT 112.385 51.595 112.555 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 112.845 48.875 113.015 49.045 ;
      RECT 112.385 48.875 112.555 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 112.845 46.155 113.015 46.325 ;
      RECT 112.385 46.155 112.555 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 112.845 43.435 113.015 43.605 ;
      RECT 112.385 43.435 112.555 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 112.845 40.715 113.015 40.885 ;
      RECT 112.385 40.715 112.555 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 112.845 37.995 113.015 38.165 ;
      RECT 112.385 37.995 112.555 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 112.845 35.275 113.015 35.445 ;
      RECT 112.385 35.275 112.555 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 112.845 32.555 113.015 32.725 ;
      RECT 112.385 32.555 112.555 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 112.845 29.835 113.015 30.005 ;
      RECT 112.385 29.835 112.555 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 112.845 27.115 113.015 27.285 ;
      RECT 112.385 27.115 112.555 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 112.845 24.395 113.015 24.565 ;
      RECT 112.385 24.395 112.555 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 112.845 21.675 113.015 21.845 ;
      RECT 112.385 21.675 112.555 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 112.845 18.955 113.015 19.125 ;
      RECT 112.385 18.955 112.555 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 112.845 16.235 113.015 16.405 ;
      RECT 112.385 16.235 112.555 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 112.845 13.515 113.015 13.685 ;
      RECT 112.385 13.515 112.555 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 112.845 10.795 113.015 10.965 ;
      RECT 112.385 10.795 112.555 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 112.845 8.075 113.015 8.245 ;
      RECT 112.385 8.075 112.555 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 112.845 5.355 113.015 5.525 ;
      RECT 112.385 5.355 112.555 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 112.845 2.635 113.015 2.805 ;
      RECT 112.385 2.635 112.555 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 112.845 -0.085 113.015 0.085 ;
      RECT 112.385 -0.085 112.555 0.085 ;
      RECT 111.925 -0.085 112.095 0.085 ;
      RECT 111.465 -0.085 111.635 0.085 ;
      RECT 111.005 -0.085 111.175 0.085 ;
      RECT 110.545 -0.085 110.715 0.085 ;
      RECT 110.085 -0.085 110.255 0.085 ;
      RECT 109.625 -0.085 109.795 0.085 ;
      RECT 109.165 -0.085 109.335 0.085 ;
      RECT 108.705 -0.085 108.875 0.085 ;
      RECT 108.245 -0.085 108.415 0.085 ;
      RECT 107.785 -0.085 107.955 0.085 ;
      RECT 107.325 -0.085 107.495 0.085 ;
      RECT 106.865 -0.085 107.035 0.085 ;
      RECT 106.405 -0.085 106.575 0.085 ;
      RECT 105.945 -0.085 106.115 0.085 ;
      RECT 105.485 -0.085 105.655 0.085 ;
      RECT 105.025 -0.085 105.195 0.085 ;
      RECT 104.565 -0.085 104.735 0.085 ;
      RECT 104.105 -0.085 104.275 0.085 ;
      RECT 103.645 -0.085 103.815 0.085 ;
      RECT 103.185 -0.085 103.355 0.085 ;
      RECT 102.725 -0.085 102.895 0.085 ;
      RECT 102.265 -0.085 102.435 0.085 ;
      RECT 101.805 -0.085 101.975 0.085 ;
      RECT 101.345 -0.085 101.515 0.085 ;
      RECT 100.885 -0.085 101.055 0.085 ;
      RECT 100.425 -0.085 100.595 0.085 ;
      RECT 99.965 -0.085 100.135 0.085 ;
      RECT 99.505 -0.085 99.675 0.085 ;
      RECT 99.045 -0.085 99.215 0.085 ;
      RECT 98.585 -0.085 98.755 0.085 ;
      RECT 98.125 -0.085 98.295 0.085 ;
      RECT 97.665 -0.085 97.835 0.085 ;
      RECT 97.205 -0.085 97.375 0.085 ;
      RECT 96.745 -0.085 96.915 0.085 ;
      RECT 96.285 -0.085 96.455 0.085 ;
      RECT 95.825 -0.085 95.995 0.085 ;
      RECT 95.365 -0.085 95.535 0.085 ;
      RECT 94.905 -0.085 95.075 0.085 ;
      RECT 94.445 -0.085 94.615 0.085 ;
      RECT 93.985 -0.085 94.155 0.085 ;
      RECT 93.525 -0.085 93.695 0.085 ;
      RECT 93.065 -0.085 93.235 0.085 ;
      RECT 92.605 -0.085 92.775 0.085 ;
      RECT 92.145 -0.085 92.315 0.085 ;
      RECT 91.685 -0.085 91.855 0.085 ;
      RECT 91.225 -0.085 91.395 0.085 ;
      RECT 90.765 -0.085 90.935 0.085 ;
      RECT 90.305 -0.085 90.475 0.085 ;
      RECT 89.845 -0.085 90.015 0.085 ;
      RECT 89.385 -0.085 89.555 0.085 ;
      RECT 88.925 -0.085 89.095 0.085 ;
      RECT 88.465 -0.085 88.635 0.085 ;
      RECT 88.005 -0.085 88.175 0.085 ;
      RECT 87.545 -0.085 87.715 0.085 ;
      RECT 87.085 -0.085 87.255 0.085 ;
      RECT 86.625 -0.085 86.795 0.085 ;
      RECT 86.165 -0.085 86.335 0.085 ;
      RECT 85.705 -0.085 85.875 0.085 ;
      RECT 85.245 -0.085 85.415 0.085 ;
      RECT 84.785 -0.085 84.955 0.085 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 56.965 103.285 57.115 103.435 ;
      RECT 27.525 103.285 27.675 103.435 ;
      RECT 62.025 101.585 62.175 101.735 ;
      RECT 48.225 101.585 48.375 101.735 ;
      RECT 56.965 76.085 57.115 76.235 ;
      RECT 27.525 76.085 27.675 76.235 ;
      RECT 108.025 74.385 108.175 74.535 ;
      RECT 109.865 1.625 110.015 1.775 ;
      RECT 56.965 -0.075 57.115 0.075 ;
      RECT 27.525 -0.075 27.675 0.075 ;
    LAYER via2 ;
      RECT 56.94 103.26 57.14 103.46 ;
      RECT 27.5 103.26 27.7 103.46 ;
      RECT 111.22 66.54 111.42 66.74 ;
      RECT 111.22 40.7 111.42 40.9 ;
      RECT 111.68 36.62 111.88 36.82 ;
      RECT 56.94 -0.1 57.14 0.1 ;
      RECT 27.5 -0.1 27.7 0.1 ;
    LAYER via3 ;
      RECT 56.94 103.26 57.14 103.46 ;
      RECT 27.5 103.26 27.7 103.46 ;
      RECT 82.7 91.7 82.9 91.9 ;
      RECT 56.94 -0.1 57.14 0.1 ;
      RECT 27.5 -0.1 27.7 0.1 ;
    LAYER via4 ;
      RECT 106.32 58.88 107.12 59.68 ;
      RECT 106.32 57.28 107.12 58.08 ;
      RECT 106.32 18.08 107.12 18.88 ;
      RECT 106.32 16.48 107.12 17.28 ;
    LAYER fieldpoly ;
      POLYGON 84.5 103.22 84.5 76.02 113.02 76.02 113.02 0.14 0.14 0.14 0.14 103.22 ;
    LAYER diff ;
      POLYGON 84.64 103.36 84.64 76.16 113.16 76.16 113.16 0 0 0 0 103.36 ;
    LAYER nwell ;
      POLYGON 84.83 102.055 84.83 99.225 83.53 99.225 83.53 100.45 80.77 100.45 80.77 102.055 ;
      RECT -0.19 99.225 3.87 102.055 ;
      POLYGON 84.83 96.615 84.83 93.785 80.77 93.785 80.77 95.39 83.53 95.39 83.53 96.615 ;
      RECT -0.19 93.785 3.87 96.615 ;
      RECT 83.99 88.345 84.83 91.175 ;
      RECT -0.19 88.345 3.87 91.175 ;
      RECT 83.99 82.905 84.83 85.735 ;
      RECT -0.19 82.905 3.87 85.735 ;
      POLYGON 84.83 80.295 84.83 77.465 80.77 77.465 80.77 79.07 83.53 79.07 83.53 80.295 ;
      RECT -0.19 77.465 3.87 80.295 ;
      POLYGON 113.35 74.855 113.35 72.025 112.51 72.025 112.51 73.25 111.13 73.25 111.13 74.855 ;
      RECT -0.19 72.025 3.87 74.855 ;
      RECT 112.05 66.585 113.35 69.415 ;
      POLYGON 2.03 69.415 2.03 68.19 3.87 68.19 3.87 66.585 -0.19 66.585 -0.19 69.415 ;
      POLYGON 113.35 63.975 113.35 61.145 112.51 61.145 112.51 62.37 112.05 62.37 112.05 63.975 ;
      RECT -0.19 61.145 3.87 63.975 ;
      RECT 112.05 55.705 113.35 58.535 ;
      RECT -0.19 55.705 3.87 58.535 ;
      RECT 112.05 50.265 113.35 53.095 ;
      RECT -0.19 50.265 3.87 53.095 ;
      POLYGON 113.35 47.655 113.35 44.825 112.05 44.825 112.05 46.05 111.13 46.05 111.13 47.655 ;
      RECT -0.19 44.825 3.87 47.655 ;
      RECT 112.05 39.385 113.35 42.215 ;
      RECT -0.19 39.385 3.87 42.215 ;
      POLYGON 113.35 36.775 113.35 33.945 111.13 33.945 111.13 35.55 112.05 35.55 112.05 36.775 ;
      RECT -0.19 33.945 3.87 36.775 ;
      RECT 112.05 28.505 113.35 31.335 ;
      RECT -0.19 28.505 3.87 31.335 ;
      RECT 112.05 23.065 113.35 25.895 ;
      RECT -0.19 23.065 3.87 25.895 ;
      RECT 112.05 17.625 113.35 20.455 ;
      RECT -0.19 17.625 3.87 20.455 ;
      RECT 112.05 12.185 113.35 15.015 ;
      RECT -0.19 12.185 3.87 15.015 ;
      RECT 112.05 6.745 113.35 9.575 ;
      RECT -0.19 6.745 3.87 9.575 ;
      RECT 112.05 1.305 113.35 4.135 ;
      RECT -0.19 1.305 3.87 4.135 ;
      POLYGON 84.64 103.36 84.64 76.16 113.16 76.16 113.16 0 0 0 0 103.36 ;
    LAYER pwell ;
      RECT 81.09 103.31 81.31 103.48 ;
      RECT 77.41 103.31 77.63 103.48 ;
      RECT 73.73 103.31 73.95 103.48 ;
      RECT 70.05 103.31 70.27 103.48 ;
      RECT 66.37 103.31 66.59 103.48 ;
      RECT 62.69 103.31 62.91 103.48 ;
      RECT 59.01 103.31 59.23 103.48 ;
      RECT 55.33 103.31 55.55 103.48 ;
      RECT 51.65 103.31 51.87 103.48 ;
      RECT 47.97 103.31 48.19 103.48 ;
      RECT 44.29 103.31 44.51 103.48 ;
      RECT 40.61 103.31 40.83 103.48 ;
      RECT 36.93 103.31 37.15 103.48 ;
      RECT 33.25 103.31 33.47 103.48 ;
      RECT 29.57 103.31 29.79 103.48 ;
      RECT 25.89 103.31 26.11 103.48 ;
      RECT 22.21 103.31 22.43 103.48 ;
      RECT 18.53 103.31 18.75 103.48 ;
      RECT 14.85 103.31 15.07 103.48 ;
      RECT 11.17 103.31 11.39 103.48 ;
      RECT 7.49 103.31 7.71 103.48 ;
      RECT 3.81 103.31 4.03 103.48 ;
      RECT 0.13 103.31 0.35 103.48 ;
      RECT 107.77 76.11 107.99 76.28 ;
      RECT 104.09 76.11 104.31 76.28 ;
      RECT 100.41 76.11 100.63 76.28 ;
      RECT 96.73 76.11 96.95 76.28 ;
      RECT 93.05 76.11 93.27 76.28 ;
      RECT 89.37 76.11 89.59 76.28 ;
      RECT 85.69 76.11 85.91 76.28 ;
      RECT 111.495 76.1 111.605 76.22 ;
      RECT 112.395 -0.05 112.555 0.06 ;
      RECT 110.575 -0.06 110.685 0.06 ;
      RECT 106.85 -0.12 107.07 0.05 ;
      RECT 103.17 -0.12 103.39 0.05 ;
      RECT 99.49 -0.12 99.71 0.05 ;
      RECT 95.81 -0.12 96.03 0.05 ;
      RECT 92.13 -0.12 92.35 0.05 ;
      RECT 88.45 -0.12 88.67 0.05 ;
      RECT 84.77 -0.12 84.99 0.05 ;
      RECT 81.09 -0.12 81.31 0.05 ;
      RECT 77.41 -0.12 77.63 0.05 ;
      RECT 73.73 -0.12 73.95 0.05 ;
      RECT 70.05 -0.12 70.27 0.05 ;
      RECT 66.37 -0.12 66.59 0.05 ;
      RECT 62.69 -0.12 62.91 0.05 ;
      RECT 59.01 -0.12 59.23 0.05 ;
      RECT 55.33 -0.12 55.55 0.05 ;
      RECT 51.65 -0.12 51.87 0.05 ;
      RECT 47.97 -0.12 48.19 0.05 ;
      RECT 44.29 -0.12 44.51 0.05 ;
      RECT 40.61 -0.12 40.83 0.05 ;
      RECT 36.93 -0.12 37.15 0.05 ;
      RECT 33.25 -0.12 33.47 0.05 ;
      RECT 29.57 -0.12 29.79 0.05 ;
      RECT 25.89 -0.12 26.11 0.05 ;
      RECT 22.21 -0.12 22.43 0.05 ;
      RECT 18.53 -0.12 18.75 0.05 ;
      RECT 14.85 -0.12 15.07 0.05 ;
      RECT 11.17 -0.12 11.39 0.05 ;
      RECT 7.49 -0.12 7.71 0.05 ;
      RECT 3.81 -0.12 4.03 0.05 ;
      RECT 0.13 -0.12 0.35 0.05 ;
      POLYGON 84.64 103.36 84.64 76.16 113.16 76.16 113.16 0 0 0 0 103.36 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 103.36 84.64 103.36 84.64 76.16 113.16 76.16 113.16 0 ;
  END
END sb_0__0_

END LIBRARY
