VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_0__2_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 92 BY 97.92 ;
  SYMMETRY X Y ;
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 90.63 92 90.93 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 74.99 92 75.29 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 65.47 92 65.77 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 76.35 92 76.65 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 32.15 92 32.45 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 60.03 92 60.33 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 51.19 92 51.49 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 45.07 92 45.37 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 64.11 92 64.41 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 29.43 92 29.73 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 69.55 92 69.85 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 73.63 92 73.93 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 35.55 92 35.85 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 19.23 92 19.53 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 36.91 92 37.21 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 40.99 92 41.29 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 57.31 92 57.61 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 70.91 92 71.21 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 49.83 92 50.13 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 68.19 92 68.49 ;
    END
  END chanx_right_in[19]
  PIN right_top_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 43.71 92 44.01 ;
    END
  END right_top_grid_pin_1_[0]
  PIN right_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.28 10.88 79.42 11.365 ;
    END
  END right_bottom_grid_pin_34_[0]
  PIN right_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.72 10.88 85.86 11.365 ;
    END
  END right_bottom_grid_pin_35_[0]
  PIN right_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.04 10.88 82.18 11.365 ;
    END
  END right_bottom_grid_pin_36_[0]
  PIN right_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.1 10.88 87.24 11.365 ;
    END
  END right_bottom_grid_pin_37_[0]
  PIN right_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.12 10.88 81.26 11.365 ;
    END
  END right_bottom_grid_pin_38_[0]
  PIN right_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.36 10.88 78.5 11.365 ;
    END
  END right_bottom_grid_pin_39_[0]
  PIN right_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.2 10.88 80.34 11.365 ;
    END
  END right_bottom_grid_pin_40_[0]
  PIN right_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.96 10.88 83.1 11.365 ;
    END
  END right_bottom_grid_pin_41_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.84 0 49.98 0.485 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.96 0 60.1 0.485 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.88 0 61.02 0.485 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.64 0 63.78 0.485 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.6 0 52.74 0.485 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 0 39.4 0.485 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 0 35.72 0.485 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.72 0 62.86 0.485 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.36 0 9.5 0.485 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.44 0 8.58 0.485 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.38 0 26.52 0.485 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.68 0 51.82 0.485 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.52 0 53.66 0.485 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 0 56.42 0.485 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.12 0 58.26 0.485 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 0 38.48 0.485 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.8 0 61.94 0.485 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.82 0 32.96 0.485 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.32 0 21.46 0.485 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.18 0 40.32 0.485 ;
    END
  END chany_bottom_in[19]
  PIN bottom_left_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.4 0 20.54 0.485 ;
    END
  END bottom_left_grid_pin_1_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 61.39 92 61.69 ;
    END
  END ccff_head[0]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 17.87 92 18.17 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 46.43 92 46.73 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 39.63 92 39.93 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 25.35 92 25.65 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 47.79 92 48.09 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 28.07 92 28.37 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 58.67 92 58.97 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 23.99 92 24.29 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 42.35 92 42.65 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 30.79 92 31.09 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 53.23 92 53.53 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 26.71 92 27.01 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 72.27 92 72.57 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 20.59 92 20.89 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 55.95 92 56.25 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 33.51 92 33.81 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 66.83 92 67.13 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 38.27 92 38.57 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 54.59 92 54.89 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 22.63 92 22.93 ;
    END
  END chanx_right_out[19]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.76 0 50.9 0.485 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.2 0 57.34 0.485 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 0 41.24 0.485 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.2 0 11.34 0.485 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.74 0 33.88 0.485 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.48 0 19.62 0.485 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.12 0 12.26 0.485 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.5 0 36.64 0.485 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.56 0 18.7 0.485 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.04 0 13.18 0.485 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.04 0 59.18 0.485 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.64 0 17.78 0.485 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.28 0 10.42 0.485 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.96 0 14.1 0.485 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.42 0 37.56 0.485 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.72 0 16.86 0.485 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.44 0 54.58 0.485 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.88 0 15.02 0.485 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.46 0 2.6 0.485 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.8 0 15.94 0.485 ;
    END
  END chany_bottom_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.66 0 34.8 0.485 ;
    END
  END ccff_tail[0]
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.7 10.88 68.84 11.365 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 14.47 92 14.77 ;
    END
  END SC_OUT_BOT
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met3 ;
        RECT 91.2 62.75 92 63.05 ;
    END
  END prog_clk_0_E_in
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 22.2 3.2 25.4 ;
        RECT 88.8 22.2 92 25.4 ;
        RECT 0 63 3.2 66.2 ;
        RECT 88.8 63 92 66.2 ;
      LAYER met4 ;
        RECT 10.74 0 11.34 0.6 ;
        RECT 40.18 0 40.78 0.6 ;
        RECT 80.66 10.88 81.26 11.48 ;
        RECT 10.74 97.32 11.34 97.92 ;
        RECT 40.18 97.32 40.78 97.92 ;
        RECT 80.66 97.32 81.26 97.92 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 65.76 2.48 66.24 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 65.76 7.92 66.24 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 91.52 13.36 92 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 91.52 18.8 92 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 91.52 24.24 92 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 91.52 29.68 92 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 91.52 35.12 92 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 91.52 40.56 92 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 91.52 46 92 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 91.52 51.44 92 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 91.52 56.88 92 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 91.52 62.32 92 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 91.52 67.76 92 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 91.52 73.2 92 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 91.52 78.64 92 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 91.52 84.08 92 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 91.52 89.52 92 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 91.52 94.96 92 95.44 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 25.46 0 26.06 0.6 ;
        RECT 54.9 0 55.5 0.6 ;
        RECT 25.46 97.32 26.06 97.92 ;
        RECT 54.9 97.32 55.5 97.92 ;
      LAYER met5 ;
        RECT 0 42.6 3.2 45.8 ;
        RECT 88.8 42.6 92 45.8 ;
        RECT 0 83.4 3.2 86.6 ;
        RECT 88.8 83.4 92 86.6 ;
      LAYER met1 ;
        RECT 0 0 45.4 0.24 ;
        RECT 46.6 0 66.24 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 65.76 5.2 66.24 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 46.6 10.64 92 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 91.52 16.08 92 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 91.52 21.52 92 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 91.52 26.96 92 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 91.52 32.4 92 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 91.52 37.84 92 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 91.52 43.28 92 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 91.52 48.72 92 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 91.52 54.16 92 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 91.52 59.6 92 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 91.52 65.04 92 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 91.52 70.48 92 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 91.52 75.92 92 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 91.52 81.36 92 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 91.52 86.8 92 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 91.52 92.24 92 92.72 ;
        RECT 0 97.68 45.4 97.92 ;
        RECT 46.6 97.68 92 97.92 ;
    END
  END VSS
  OBS
    LAYER met3 ;
      POLYGON 55.365 98.085 55.365 98.08 55.58 98.08 55.58 97.76 55.365 97.76 55.365 97.755 55.035 97.755 55.035 97.76 54.82 97.76 54.82 98.08 55.035 98.08 55.035 98.085 ;
      POLYGON 25.925 98.085 25.925 98.08 26.14 98.08 26.14 97.76 25.925 97.76 25.925 97.755 25.595 97.755 25.595 97.76 25.38 97.76 25.38 98.08 25.595 98.08 25.595 98.085 ;
      POLYGON 74.915 11.385 74.915 11.055 74.585 11.055 74.585 11.07 58.04 11.07 58.04 11.37 74.585 11.37 74.585 11.385 ;
      POLYGON 55.365 0.165 55.365 0.16 55.58 0.16 55.58 -0.16 55.365 -0.16 55.365 -0.165 55.035 -0.165 55.035 -0.16 54.82 -0.16 54.82 0.16 55.035 0.16 55.035 0.165 ;
      POLYGON 25.925 0.165 25.925 0.16 26.14 0.16 26.14 -0.16 25.925 -0.16 25.925 -0.165 25.595 -0.165 25.595 -0.16 25.38 -0.16 25.38 0.16 25.595 0.16 25.595 0.165 ;
      POLYGON 91.6 97.52 91.6 91.33 90.8 91.33 90.8 90.23 91.6 90.23 91.6 77.05 90.8 77.05 90.8 75.95 91.6 75.95 91.6 75.69 90.8 75.69 90.8 74.59 91.6 74.59 91.6 74.33 90.8 74.33 90.8 73.23 91.6 73.23 91.6 72.97 90.8 72.97 90.8 71.87 91.6 71.87 91.6 71.61 90.8 71.61 90.8 70.51 91.6 70.51 91.6 70.25 90.8 70.25 90.8 69.15 91.6 69.15 91.6 68.89 90.8 68.89 90.8 67.79 91.6 67.79 91.6 67.53 90.8 67.53 90.8 66.43 91.6 66.43 91.6 66.17 90.8 66.17 90.8 65.07 91.6 65.07 91.6 64.81 90.8 64.81 90.8 63.71 91.6 63.71 91.6 63.45 90.8 63.45 90.8 62.35 91.6 62.35 91.6 62.09 90.8 62.09 90.8 60.99 91.6 60.99 91.6 60.73 90.8 60.73 90.8 59.63 91.6 59.63 91.6 59.37 90.8 59.37 90.8 58.27 91.6 58.27 91.6 58.01 90.8 58.01 90.8 56.91 91.6 56.91 91.6 56.65 90.8 56.65 90.8 55.55 91.6 55.55 91.6 55.29 90.8 55.29 90.8 54.19 91.6 54.19 91.6 53.93 90.8 53.93 90.8 52.83 91.6 52.83 91.6 51.89 90.8 51.89 90.8 50.79 91.6 50.79 91.6 50.53 90.8 50.53 90.8 49.43 91.6 49.43 91.6 48.49 90.8 48.49 90.8 47.39 91.6 47.39 91.6 47.13 90.8 47.13 90.8 46.03 91.6 46.03 91.6 45.77 90.8 45.77 90.8 44.67 91.6 44.67 91.6 44.41 90.8 44.41 90.8 43.31 91.6 43.31 91.6 43.05 90.8 43.05 90.8 41.95 91.6 41.95 91.6 41.69 90.8 41.69 90.8 40.59 91.6 40.59 91.6 40.33 90.8 40.33 90.8 39.23 91.6 39.23 91.6 38.97 90.8 38.97 90.8 37.87 91.6 37.87 91.6 37.61 90.8 37.61 90.8 36.51 91.6 36.51 91.6 36.25 90.8 36.25 90.8 35.15 91.6 35.15 91.6 34.21 90.8 34.21 90.8 33.11 91.6 33.11 91.6 32.85 90.8 32.85 90.8 31.75 91.6 31.75 91.6 31.49 90.8 31.49 90.8 30.39 91.6 30.39 91.6 30.13 90.8 30.13 90.8 29.03 91.6 29.03 91.6 28.77 90.8 28.77 90.8 27.67 91.6 27.67 91.6 27.41 90.8 27.41 90.8 26.31 91.6 26.31 91.6 26.05 90.8 26.05 90.8 24.95 91.6 24.95 91.6 24.69 90.8 24.69 90.8 23.59 91.6 23.59 91.6 23.33 90.8 23.33 90.8 22.23 91.6 22.23 91.6 21.29 90.8 21.29 90.8 20.19 91.6 20.19 91.6 19.93 90.8 19.93 90.8 18.83 91.6 18.83 91.6 18.57 90.8 18.57 90.8 17.47 91.6 17.47 91.6 15.17 90.8 15.17 90.8 14.07 91.6 14.07 91.6 11.28 65.84 11.28 65.84 0.4 0.4 0.4 0.4 97.52 ;
    LAYER met2 ;
      RECT 55.06 97.735 55.34 98.105 ;
      RECT 25.62 97.735 25.9 98.105 ;
      POLYGON 39.86 21.32 39.86 0.24 39.9 0.24 39.9 0.1 39.72 0.1 39.72 21.32 ;
      POLYGON 74.82 12.14 74.82 11.405 74.89 11.405 74.89 11.035 74.61 11.035 74.61 11.405 74.68 11.405 74.68 12.14 ;
      POLYGON 63.32 6.02 63.32 0.24 63.36 0.24 63.36 0.1 63.18 0.1 63.18 6.02 ;
      POLYGON 14.56 5.17 14.56 0.1 14.38 0.1 14.38 0.24 14.42 0.24 14.42 5.17 ;
      RECT 64.04 0.35 64.3 0.67 ;
      RECT 55.06 -0.185 55.34 0.185 ;
      RECT 25.62 -0.185 25.9 0.185 ;
      POLYGON 91.72 97.64 91.72 11.16 87.52 11.16 87.52 11.645 86.82 11.645 86.82 11.16 86.14 11.16 86.14 11.645 85.44 11.645 85.44 11.16 83.38 11.16 83.38 11.645 82.68 11.645 82.68 11.16 82.46 11.16 82.46 11.645 81.76 11.645 81.76 11.16 81.54 11.16 81.54 11.645 80.84 11.645 80.84 11.16 80.62 11.16 80.62 11.645 79.92 11.645 79.92 11.16 79.7 11.16 79.7 11.645 79 11.645 79 11.16 78.78 11.16 78.78 11.645 78.08 11.645 78.08 11.16 69.12 11.16 69.12 11.645 68.42 11.645 68.42 11.16 65.96 11.16 65.96 0.28 64.06 0.28 64.06 0.765 63.36 0.765 63.36 0.28 63.14 0.28 63.14 0.765 62.44 0.765 62.44 0.28 62.22 0.28 62.22 0.765 61.52 0.765 61.52 0.28 61.3 0.28 61.3 0.765 60.6 0.765 60.6 0.28 60.38 0.28 60.38 0.765 59.68 0.765 59.68 0.28 59.46 0.28 59.46 0.765 58.76 0.765 58.76 0.28 58.54 0.28 58.54 0.765 57.84 0.765 57.84 0.28 57.62 0.28 57.62 0.765 56.92 0.765 56.92 0.28 56.7 0.28 56.7 0.765 56 0.765 56 0.28 54.86 0.28 54.86 0.765 54.16 0.765 54.16 0.28 53.94 0.28 53.94 0.765 53.24 0.765 53.24 0.28 53.02 0.28 53.02 0.765 52.32 0.765 52.32 0.28 52.1 0.28 52.1 0.765 51.4 0.765 51.4 0.28 51.18 0.28 51.18 0.765 50.48 0.765 50.48 0.28 50.26 0.28 50.26 0.765 49.56 0.765 49.56 0.28 41.52 0.28 41.52 0.765 40.82 0.765 40.82 0.28 40.6 0.28 40.6 0.765 39.9 0.765 39.9 0.28 39.68 0.28 39.68 0.765 38.98 0.765 38.98 0.28 38.76 0.28 38.76 0.765 38.06 0.765 38.06 0.28 37.84 0.28 37.84 0.765 37.14 0.765 37.14 0.28 36.92 0.28 36.92 0.765 36.22 0.765 36.22 0.28 36 0.28 36 0.765 35.3 0.765 35.3 0.28 35.08 0.28 35.08 0.765 34.38 0.765 34.38 0.28 34.16 0.28 34.16 0.765 33.46 0.765 33.46 0.28 33.24 0.28 33.24 0.765 32.54 0.765 32.54 0.28 26.8 0.28 26.8 0.765 26.1 0.765 26.1 0.28 21.74 0.28 21.74 0.765 21.04 0.765 21.04 0.28 20.82 0.28 20.82 0.765 20.12 0.765 20.12 0.28 19.9 0.28 19.9 0.765 19.2 0.765 19.2 0.28 18.98 0.28 18.98 0.765 18.28 0.765 18.28 0.28 18.06 0.28 18.06 0.765 17.36 0.765 17.36 0.28 17.14 0.28 17.14 0.765 16.44 0.765 16.44 0.28 16.22 0.28 16.22 0.765 15.52 0.765 15.52 0.28 15.3 0.28 15.3 0.765 14.6 0.765 14.6 0.28 14.38 0.28 14.38 0.765 13.68 0.765 13.68 0.28 13.46 0.28 13.46 0.765 12.76 0.765 12.76 0.28 12.54 0.28 12.54 0.765 11.84 0.765 11.84 0.28 11.62 0.28 11.62 0.765 10.92 0.765 10.92 0.28 10.7 0.28 10.7 0.765 10 0.765 10 0.28 9.78 0.28 9.78 0.765 9.08 0.765 9.08 0.28 8.86 0.28 8.86 0.765 8.16 0.765 8.16 0.28 2.88 0.28 2.88 0.765 2.18 0.765 2.18 0.28 0.28 0.28 0.28 97.64 ;
    LAYER met1 ;
      RECT 45.68 97.68 46.32 98.16 ;
      POLYGON 82.27 11.52 82.27 11.26 81.95 11.26 81.95 11.32 80.015 11.32 80.015 11.275 79.725 11.275 79.725 11.32 76.29 11.32 76.29 11.26 75.97 11.26 75.97 11.52 76.29 11.52 76.29 11.46 79.725 11.46 79.725 11.505 80.015 11.505 80.015 11.46 81.95 11.46 81.95 11.52 ;
      POLYGON 65.71 11.52 65.71 11.26 65.39 11.26 65.39 11.32 62.935 11.32 62.935 11.275 62.645 11.275 62.645 11.505 62.935 11.505 62.935 11.46 65.39 11.46 65.39 11.52 ;
      POLYGON 56.97 11.52 56.97 11.505 57.015 11.505 57.015 11.275 56.97 11.275 56.97 11.26 56.65 11.26 56.65 11.52 ;
      POLYGON 56.05 11.52 56.05 11.26 55.73 11.26 55.73 11.32 55.115 11.32 55.115 11.275 54.825 11.275 54.825 11.505 55.115 11.505 55.115 11.46 55.73 11.46 55.73 11.52 ;
      POLYGON 52.37 11.52 52.37 11.26 52.05 11.26 52.05 11.32 51.435 11.32 51.435 11.275 51.145 11.275 51.145 11.505 51.435 11.505 51.435 11.46 52.05 11.46 52.05 11.52 ;
      RECT 55.73 10.24 56.05 10.5 ;
      POLYGON 52.37 10.5 52.37 10.24 52.05 10.24 52.05 10.3 51.895 10.3 51.895 10.255 51.605 10.255 51.605 10.485 51.895 10.485 51.895 10.44 52.05 10.44 52.05 10.5 ;
      POLYGON 50.99 10.5 50.99 10.24 50.67 10.24 50.67 10.3 49.595 10.3 49.595 10.255 49.305 10.255 49.305 10.485 49.595 10.485 49.595 10.44 50.67 10.44 50.67 10.5 ;
      POLYGON 64.33 0.64 64.33 0.38 64.01 0.38 64.01 0.44 59.255 0.44 59.255 0.395 58.965 0.395 58.965 0.625 59.255 0.625 59.255 0.58 64.01 0.58 64.01 0.64 ;
      POLYGON 58.35 0.64 58.35 0.38 58.03 0.38 58.03 0.44 56.955 0.44 56.955 0.395 56.665 0.395 56.665 0.625 56.955 0.625 56.955 0.58 58.03 0.58 58.03 0.64 ;
      POLYGON 50.99 0.64 50.99 0.38 50.67 0.38 50.67 0.44 49.225 0.44 49.225 0.395 48.935 0.395 48.935 0.625 49.225 0.625 49.225 0.58 50.67 0.58 50.67 0.64 ;
      RECT 45.61 0.38 45.93 0.64 ;
      POLYGON 38.57 0.64 38.57 0.58 43.325 0.58 43.325 0.625 43.615 0.625 43.615 0.395 43.325 0.395 43.325 0.44 38.57 0.44 38.57 0.38 38.25 0.38 38.25 0.64 ;
      RECT 45.68 -0.24 46.32 0.24 ;
      POLYGON 46.32 97.64 46.32 97.4 91.72 97.4 91.72 95.72 91.24 95.72 91.24 94.68 91.72 94.68 91.72 93 91.24 93 91.24 91.96 91.72 91.96 91.72 90.28 91.24 90.28 91.24 89.24 91.72 89.24 91.72 87.56 91.24 87.56 91.24 86.52 91.72 86.52 91.72 84.84 91.24 84.84 91.24 83.8 91.72 83.8 91.72 82.12 91.24 82.12 91.24 81.08 91.72 81.08 91.72 79.4 91.24 79.4 91.24 78.36 91.72 78.36 91.72 76.68 91.24 76.68 91.24 75.64 91.72 75.64 91.72 73.96 91.24 73.96 91.24 72.92 91.72 72.92 91.72 71.24 91.24 71.24 91.24 70.2 91.72 70.2 91.72 68.52 91.24 68.52 91.24 67.48 91.72 67.48 91.72 65.8 91.24 65.8 91.24 64.76 91.72 64.76 91.72 63.08 91.24 63.08 91.24 62.04 91.72 62.04 91.72 60.36 91.24 60.36 91.24 59.32 91.72 59.32 91.72 57.64 91.24 57.64 91.24 56.6 91.72 56.6 91.72 54.92 91.24 54.92 91.24 53.88 91.72 53.88 91.72 52.2 91.24 52.2 91.24 51.16 91.72 51.16 91.72 49.48 91.24 49.48 91.24 48.44 91.72 48.44 91.72 46.76 91.24 46.76 91.24 45.72 91.72 45.72 91.72 44.04 91.24 44.04 91.24 43 91.72 43 91.72 41.32 91.24 41.32 91.24 40.28 91.72 40.28 91.72 38.6 91.24 38.6 91.24 37.56 91.72 37.56 91.72 35.88 91.24 35.88 91.24 34.84 91.72 34.84 91.72 33.16 91.24 33.16 91.24 32.12 91.72 32.12 91.72 30.44 91.24 30.44 91.24 29.4 91.72 29.4 91.72 27.72 91.24 27.72 91.24 26.68 91.72 26.68 91.72 25 91.24 25 91.24 23.96 91.72 23.96 91.72 22.28 91.24 22.28 91.24 21.24 91.72 21.24 91.72 19.56 91.24 19.56 91.24 18.52 91.72 18.52 91.72 16.84 91.24 16.84 91.24 15.8 91.72 15.8 91.72 14.12 91.24 14.12 91.24 13.08 91.72 13.08 91.72 11.4 46.32 11.4 46.32 10.36 65.96 10.36 65.96 8.68 65.48 8.68 65.48 7.64 65.96 7.64 65.96 5.96 65.48 5.96 65.48 4.92 65.96 4.92 65.96 3.24 65.48 3.24 65.48 2.2 65.96 2.2 65.96 0.52 46.32 0.52 46.32 0.28 45.68 0.28 45.68 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 45.68 97.4 45.68 97.64 ;
    LAYER met4 ;
      POLYGON 91.6 97.52 91.6 11.28 81.66 11.28 81.66 11.88 80.26 11.88 80.26 11.28 65.84 11.28 65.84 0.4 55.9 0.4 55.9 1 54.5 1 54.5 0.4 41.18 0.4 41.18 1 39.78 1 39.78 0.4 26.46 0.4 26.46 1 25.06 1 25.06 0.4 11.74 0.4 11.74 1 10.34 1 10.34 0.4 0.4 0.4 0.4 97.52 10.34 97.52 10.34 96.92 11.74 96.92 11.74 97.52 25.06 97.52 25.06 96.92 26.46 96.92 26.46 97.52 39.78 97.52 39.78 96.92 41.18 96.92 41.18 97.52 54.5 97.52 54.5 96.92 55.9 96.92 55.9 97.52 80.26 97.52 80.26 96.92 81.66 96.92 81.66 97.52 ;
    LAYER met5 ;
      POLYGON 90.4 96.32 90.4 88.2 87.2 88.2 87.2 81.8 90.4 81.8 90.4 67.8 87.2 67.8 87.2 61.4 90.4 61.4 90.4 47.4 87.2 47.4 87.2 41 90.4 41 90.4 27 87.2 27 87.2 20.6 90.4 20.6 90.4 12.48 64.64 12.48 64.64 1.6 1.6 1.6 1.6 20.6 4.8 20.6 4.8 27 1.6 27 1.6 41 4.8 41 4.8 47.4 1.6 47.4 1.6 61.4 4.8 61.4 4.8 67.8 1.6 67.8 1.6 81.8 4.8 81.8 4.8 88.2 1.6 88.2 1.6 96.32 ;
    LAYER li1 ;
      POLYGON 92 98.005 92 97.835 89.615 97.835 89.615 97.11 89.325 97.11 89.325 97.835 82.255 97.835 82.255 97.11 81.965 97.11 81.965 97.835 67.535 97.835 67.535 97.11 67.245 97.11 67.245 97.835 52.355 97.835 52.355 97.11 52.065 97.11 52.065 97.835 37.635 97.835 37.635 97.11 37.345 97.11 37.345 97.835 22.455 97.835 22.455 97.11 22.165 97.11 22.165 97.835 7.735 97.835 7.735 97.11 7.445 97.11 7.445 97.835 0 97.835 0 98.005 ;
      RECT 91.54 95.115 92 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 91.54 92.395 92 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 91.54 89.675 92 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 91.54 86.955 92 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 91.54 84.235 92 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 91.54 81.515 92 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 91.54 78.795 92 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 91.08 76.075 92 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 91.08 73.355 92 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 88.32 70.635 92 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 88.32 67.915 92 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 91.54 65.195 92 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 91.54 62.475 92 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 90.16 59.755 92 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 90.16 57.035 92 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 91.54 54.315 92 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 91.54 51.595 92 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 91.08 48.875 92 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 91.08 46.155 92 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 91.54 43.435 92 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 91.54 40.715 92 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 91.08 37.995 92 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 91.08 35.275 92 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 91.08 32.555 92 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 91.08 29.835 92 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 91.08 27.115 92 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 91.08 24.395 92 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 91.08 21.675 92 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 91.08 18.955 92 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 91.08 16.235 92 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 91.08 13.515 92 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      POLYGON 75.07 11.785 75.07 10.965 78.255 10.965 78.255 11.365 78.585 11.365 78.585 10.965 80.545 10.965 80.545 11.5 81.055 11.5 81.055 10.965 81.965 10.965 81.965 11.69 82.255 11.69 82.255 10.965 84.615 10.965 84.615 11.445 84.785 11.445 84.785 10.965 85.455 10.965 85.455 11.445 85.625 11.445 85.625 10.965 86.215 10.965 86.215 11.445 86.545 11.445 86.545 10.965 87.055 10.965 87.055 11.445 87.385 11.445 87.385 10.965 87.895 10.965 87.895 11.765 88.225 11.765 88.225 10.965 89.325 10.965 89.325 11.69 89.615 11.69 89.615 10.965 92 10.965 92 10.795 63.02 10.795 63.02 10.965 67.245 10.965 67.245 11.69 67.535 11.69 67.535 10.965 69.095 10.965 69.095 11.765 69.425 11.765 69.425 10.965 69.935 10.965 69.935 11.445 70.265 11.445 70.265 10.965 70.775 10.965 70.775 11.445 71.105 11.445 71.105 10.965 71.695 10.965 71.695 11.445 71.865 11.445 71.865 10.965 72.535 10.965 72.535 11.445 72.705 11.445 72.705 10.965 74.84 10.965 74.84 11.785 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 65.32 8.075 66.24 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 65.32 5.355 66.24 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 65.32 2.635 66.24 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      POLYGON 50.505 0.885 50.505 0.085 52.065 0.085 52.065 0.81 52.355 0.81 52.355 0.085 56.025 0.085 56.025 0.62 56.535 0.62 56.535 0.085 58.495 0.085 58.495 0.485 58.825 0.485 58.825 0.085 59.425 0.085 59.425 0.81 59.715 0.81 59.715 0.085 66.24 0.085 66.24 -0.085 0 -0.085 0 0.085 3.315 0.085 3.315 0.885 3.645 0.885 3.645 0.085 4.155 0.085 4.155 0.565 4.485 0.565 4.485 0.085 4.995 0.085 4.995 0.565 5.325 0.565 5.325 0.085 5.915 0.085 5.915 0.565 6.085 0.565 6.085 0.085 6.755 0.085 6.755 0.565 6.925 0.565 6.925 0.085 7.445 0.085 7.445 0.81 7.735 0.81 7.735 0.085 13.855 0.085 13.855 0.465 14.185 0.465 14.185 0.085 14.795 0.085 14.795 0.545 15.045 0.545 15.045 0.085 16.74 0.085 16.74 0.585 17.11 0.585 17.11 0.085 18.965 0.085 18.965 0.615 19.135 0.615 19.135 0.085 19.965 0.085 19.965 0.565 20.135 0.565 20.135 0.085 20.835 0.085 20.835 0.56 21.005 0.56 21.005 0.085 21.685 0.085 21.685 0.56 21.855 0.56 21.855 0.085 22.165 0.085 22.165 0.81 22.455 0.81 22.455 0.085 22.975 0.085 22.975 0.565 23.145 0.565 23.145 0.085 23.815 0.085 23.815 0.565 23.985 0.565 23.985 0.085 24.575 0.085 24.575 0.565 24.905 0.565 24.905 0.085 25.415 0.085 25.415 0.565 25.745 0.565 25.745 0.085 26.255 0.085 26.255 0.885 26.585 0.885 26.585 0.085 29.875 0.085 29.875 0.565 30.045 0.565 30.045 0.085 30.715 0.085 30.715 0.565 30.885 0.565 30.885 0.085 31.475 0.085 31.475 0.565 31.805 0.565 31.805 0.085 32.315 0.085 32.315 0.565 32.645 0.565 32.645 0.085 33.155 0.085 33.155 0.885 33.485 0.885 33.485 0.085 37.345 0.085 37.345 0.81 37.635 0.81 37.635 0.085 38.155 0.085 38.155 0.565 38.325 0.565 38.325 0.085 38.995 0.085 38.995 0.565 39.165 0.565 39.165 0.085 39.755 0.085 39.755 0.565 40.085 0.565 40.085 0.085 40.595 0.085 40.595 0.565 40.925 0.565 40.925 0.085 41.435 0.085 41.435 0.885 41.765 0.885 41.765 0.085 42.685 0.085 42.685 0.62 43.195 0.62 43.195 0.085 45.155 0.085 45.155 0.485 45.485 0.485 45.485 0.085 46.895 0.085 46.895 0.565 47.065 0.565 47.065 0.085 47.735 0.085 47.735 0.565 47.905 0.565 47.905 0.085 48.495 0.085 48.495 0.565 48.825 0.565 48.825 0.085 49.335 0.085 49.335 0.565 49.665 0.565 49.665 0.085 50.175 0.085 50.175 0.885 ;
      POLYGON 91.83 97.75 91.83 11.05 66.07 11.05 66.07 0.17 0.17 0.17 0.17 97.75 ;
    LAYER mcon ;
      RECT 79.785 11.305 79.955 11.475 ;
      RECT 62.705 11.305 62.875 11.475 ;
      RECT 56.785 11.305 56.955 11.475 ;
      RECT 54.885 11.305 55.055 11.475 ;
      RECT 51.205 11.305 51.375 11.475 ;
      RECT 55.805 10.285 55.975 10.455 ;
      RECT 51.665 10.285 51.835 10.455 ;
      RECT 49.365 10.285 49.535 10.455 ;
      RECT 59.025 0.425 59.195 0.595 ;
      RECT 56.725 0.425 56.895 0.595 ;
      RECT 48.995 0.425 49.165 0.595 ;
      RECT 43.385 0.425 43.555 0.595 ;
    LAYER via ;
      RECT 55.125 97.845 55.275 97.995 ;
      RECT 25.685 97.845 25.835 97.995 ;
      RECT 82.035 11.315 82.185 11.465 ;
      RECT 76.055 11.315 76.205 11.465 ;
      RECT 65.475 11.315 65.625 11.465 ;
      RECT 56.735 11.315 56.885 11.465 ;
      RECT 55.815 11.315 55.965 11.465 ;
      RECT 52.135 11.315 52.285 11.465 ;
      RECT 55.125 10.805 55.275 10.955 ;
      RECT 55.815 10.295 55.965 10.445 ;
      RECT 52.135 10.295 52.285 10.445 ;
      RECT 50.755 10.295 50.905 10.445 ;
      RECT 64.095 0.435 64.245 0.585 ;
      RECT 58.115 0.435 58.265 0.585 ;
      RECT 50.755 0.435 50.905 0.585 ;
      RECT 38.335 0.435 38.485 0.585 ;
      RECT 55.125 -0.075 55.275 0.075 ;
      RECT 25.685 -0.075 25.835 0.075 ;
    LAYER via2 ;
      RECT 55.1 97.82 55.3 98.02 ;
      RECT 25.66 97.82 25.86 98.02 ;
      RECT 90.75 64.16 90.95 64.36 ;
      RECT 74.65 11.12 74.85 11.32 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER via3 ;
      RECT 55.1 97.82 55.3 98.02 ;
      RECT 25.66 97.82 25.86 98.02 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 97.92 92 97.92 92 10.88 66.24 10.88 66.24 0 ;
  END
END sb_0__2_

END LIBRARY
