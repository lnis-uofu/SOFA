VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_0__0_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 95.68 BY 97.92 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met3 ;
        RECT 94.3 6.65 95.68 6.95 ;
    END
  END prog_clk[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.33 96.56 41.47 97.92 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.11 96.56 61.25 97.92 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.37 96.56 52.51 97.92 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.19 96.56 60.33 97.92 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.55 96.56 44.69 97.92 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.03 96.56 62.17 97.92 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.33 96.56 18.47 97.92 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.41 96.56 40.55 97.92 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.49 96.56 39.63 97.92 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 17.33 96.56 17.63 97.92 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 54.13 96.56 54.43 97.92 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 96.56 57.57 97.92 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.21 96.56 54.35 97.92 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.95 96.56 63.09 97.92 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.73 96.56 13.87 97.92 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.41 96.56 17.55 97.92 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.97 96.56 34.11 97.92 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.33 96.56 63.63 97.92 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.89 96.56 34.19 97.92 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.89 96.56 35.03 97.92 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.45 96.56 51.59 97.92 ;
    END
  END top_left_grid_pin_1_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 76.69 95.68 76.99 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 25.69 95.68 25.99 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 13.45 95.68 13.75 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 39.29 95.68 39.59 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 37.93 95.68 38.23 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 40.65 95.68 40.95 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 27.05 95.68 27.35 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 52.89 95.68 53.19 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 75.33 95.68 75.63 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 46.09 95.68 46.39 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 44.73 95.68 45.03 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 21.61 95.68 21.91 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 10.73 95.68 11.03 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 70.57 95.68 70.87 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 61.73 95.68 62.03 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 71.93 95.68 72.23 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 22.97 95.68 23.27 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 9.37 95.68 9.67 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 31.13 95.68 31.43 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 28.41 95.68 28.71 ;
    END
  END chanx_right_in[19]
  PIN right_bottom_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 60.37 95.68 60.67 ;
    END
  END right_bottom_grid_pin_1_[0]
  PIN right_bottom_grid_pin_3_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 56.97 95.68 57.27 ;
    END
  END right_bottom_grid_pin_3_[0]
  PIN right_bottom_grid_pin_5_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 66.49 95.68 66.79 ;
    END
  END right_bottom_grid_pin_5_[0]
  PIN right_bottom_grid_pin_7_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 43.37 95.68 43.67 ;
    END
  END right_bottom_grid_pin_7_[0]
  PIN right_bottom_grid_pin_9_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 69.21 95.68 69.51 ;
    END
  END right_bottom_grid_pin_9_[0]
  PIN right_bottom_grid_pin_11_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 55.61 95.68 55.91 ;
    END
  END right_bottom_grid_pin_11_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 12.09 95.68 12.39 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.29 96.56 53.43 97.92 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.65 96.56 14.79 97.92 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.71 96.56 65.85 97.92 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.49 96.56 16.63 97.92 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.33 96.56 64.47 97.92 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.81 96.56 35.95 97.92 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.57 96.56 38.71 97.92 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.73 96.56 36.87 97.92 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.57 96.56 15.71 97.92 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.65 96.56 37.79 97.92 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.13 96.56 55.27 97.92 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.49 96.56 61.79 97.92 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.35 96.56 58.49 97.92 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.41 96.56 39.71 97.92 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.49 96.56 15.79 97.92 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.73 96.56 36.03 97.92 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.27 96.56 59.41 97.92 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.65 96.56 59.95 97.92 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 57.81 96.56 58.11 97.92 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.57 96.56 37.87 97.92 ;
    END
  END chany_top_out[19]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 81.45 95.68 81.75 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 65.13 95.68 65.43 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 80.09 95.68 80.39 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 58.33 95.68 58.63 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 24.33 95.68 24.63 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 63.77 95.68 64.07 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 78.73 95.68 79.03 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 42.01 95.68 42.31 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 54.25 95.68 54.55 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 73.97 95.68 74.27 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 47.45 95.68 47.75 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 82.81 95.68 83.11 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 32.49 95.68 32.79 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 35.21 95.68 35.51 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 33.85 95.68 34.15 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 51.53 95.68 51.83 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 48.81 95.68 49.11 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 50.17 95.68 50.47 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 67.85 95.68 68.15 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 29.77 95.68 30.07 ;
    END
  END chanx_right_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.69 0 25.83 1.36 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 95.2 2.48 95.68 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 95.2 7.92 95.68 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 95.2 13.36 95.68 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 95.2 18.8 95.68 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 95.2 24.24 95.68 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 95.2 29.68 95.68 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 95.2 35.12 95.68 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 95.2 40.56 95.68 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 95.2 46 95.68 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 95.2 51.44 95.68 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 95.2 56.88 95.68 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 95.2 62.32 95.68 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 95.2 67.76 95.68 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 95.2 73.2 95.68 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 95.2 78.64 95.68 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 95.2 84.08 95.68 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 67.6 89.52 68.08 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 67.6 94.96 68.08 95.44 ;
      LAYER met4 ;
        RECT 11.66 0 12.26 0.6 ;
        RECT 41.1 0 41.7 0.6 ;
        RECT 85.26 0 85.86 0.6 ;
        RECT 85.26 86.44 85.86 87.04 ;
        RECT 11.66 97.32 12.26 97.92 ;
        RECT 41.1 97.32 41.7 97.92 ;
      LAYER met5 ;
        RECT 0 11.32 3.2 14.52 ;
        RECT 92.48 11.32 95.68 14.52 ;
        RECT 0 52.12 3.2 55.32 ;
        RECT 92.48 52.12 95.68 55.32 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 0 95.68 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 95.2 5.2 95.68 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 95.2 10.64 95.68 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 95.2 16.08 95.68 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 95.2 21.52 95.68 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 95.2 26.96 95.68 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 95.2 32.4 95.68 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 95.2 37.84 95.68 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 95.2 43.28 95.68 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 95.2 48.72 95.68 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 95.2 54.16 95.68 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 95.2 59.6 95.68 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 95.2 65.04 95.68 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 95.2 70.48 95.68 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 95.2 75.92 95.68 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 95.2 81.36 95.68 81.84 ;
        RECT 0 86.8 95.68 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 67.6 92.24 68.08 92.72 ;
        RECT 0 97.68 68.08 97.92 ;
      LAYER met4 ;
        RECT 26.38 0 26.98 0.6 ;
        RECT 55.82 0 56.42 0.6 ;
        RECT 26.38 97.32 26.98 97.92 ;
        RECT 55.82 97.32 56.42 97.92 ;
      LAYER met5 ;
        RECT 0 31.72 3.2 34.92 ;
        RECT 92.48 31.72 95.68 34.92 ;
        RECT 0 72.52 3.2 75.72 ;
        RECT 92.48 72.52 95.68 75.72 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 0 97.835 68.08 98.005 ;
      RECT 67.16 95.115 68.08 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 67.16 92.395 68.08 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 67.16 89.675 68.08 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 65.32 86.955 95.68 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 95.22 84.235 95.68 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 95.22 81.515 95.68 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 94.76 78.795 95.68 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 94.76 76.075 95.68 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 94.76 73.355 95.68 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 94.76 70.635 95.68 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 94.76 67.915 95.68 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 94.76 65.195 95.68 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 94.76 62.475 95.68 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 94.76 59.755 95.68 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 94.76 57.035 95.68 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 94.76 54.315 95.68 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 94.76 51.595 95.68 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 94.76 48.875 95.68 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 94.76 46.155 95.68 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 94.76 43.435 95.68 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 94.76 40.715 95.68 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 94.76 37.995 95.68 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 93.84 35.275 95.68 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 93.84 32.555 95.68 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 94.76 29.835 95.68 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 94.76 27.115 95.68 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 95.22 24.395 95.68 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 95.22 21.675 95.68 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 95.22 18.955 95.68 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 94.76 16.235 95.68 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 92 13.515 95.68 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 92 10.795 95.68 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 95.22 8.075 95.68 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 95.22 5.355 95.68 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 95.22 2.635 95.68 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 95.68 0.085 ;
    LAYER met3 ;
      POLYGON 56.285 98.085 56.285 98.08 56.5 98.08 56.5 97.76 56.285 97.76 56.285 97.755 55.955 97.755 55.955 97.76 55.74 97.76 55.74 98.08 55.955 98.08 55.955 98.085 ;
      POLYGON 26.845 98.085 26.845 98.08 27.06 98.08 27.06 97.76 26.845 97.76 26.845 97.755 26.515 97.755 26.515 97.76 26.3 97.76 26.3 98.08 26.515 98.08 26.515 98.085 ;
      POLYGON 94.45 67.47 94.45 67.19 93.9 67.19 93.9 67.17 79.89 67.17 79.89 67.47 ;
      POLYGON 56.285 0.165 56.285 0.16 56.5 0.16 56.5 -0.16 56.285 -0.16 56.285 -0.165 55.955 -0.165 55.955 -0.16 55.74 -0.16 55.74 0.16 55.955 0.16 55.955 0.165 ;
      POLYGON 26.845 0.165 26.845 0.16 27.06 0.16 27.06 -0.16 26.845 -0.16 26.845 -0.165 26.515 -0.165 26.515 -0.16 26.3 -0.16 26.3 0.16 26.515 0.16 26.515 0.165 ;
      POLYGON 67.68 97.52 67.68 86.64 95.28 86.64 95.28 83.51 93.9 83.51 93.9 82.41 95.28 82.41 95.28 82.15 93.9 82.15 93.9 81.05 95.28 81.05 95.28 80.79 93.9 80.79 93.9 79.69 95.28 79.69 95.28 79.43 93.9 79.43 93.9 78.33 95.28 78.33 95.28 77.39 93.9 77.39 93.9 76.29 95.28 76.29 95.28 76.03 93.9 76.03 93.9 74.93 95.28 74.93 95.28 74.67 93.9 74.67 93.9 73.57 95.28 73.57 95.28 72.63 93.9 72.63 93.9 71.53 95.28 71.53 95.28 71.27 93.9 71.27 93.9 70.17 95.28 70.17 95.28 69.91 93.9 69.91 93.9 68.81 95.28 68.81 95.28 68.55 93.9 68.55 93.9 67.45 95.28 67.45 95.28 67.19 93.9 67.19 93.9 66.09 95.28 66.09 95.28 65.83 93.9 65.83 93.9 64.73 95.28 64.73 95.28 64.47 93.9 64.47 93.9 63.37 95.28 63.37 95.28 62.43 93.9 62.43 93.9 61.33 95.28 61.33 95.28 61.07 93.9 61.07 93.9 59.97 95.28 59.97 95.28 59.03 93.9 59.03 93.9 57.93 95.28 57.93 95.28 57.67 93.9 57.67 93.9 56.57 95.28 56.57 95.28 56.31 93.9 56.31 93.9 55.21 95.28 55.21 95.28 54.95 93.9 54.95 93.9 53.85 95.28 53.85 95.28 53.59 93.9 53.59 93.9 52.49 95.28 52.49 95.28 52.23 93.9 52.23 93.9 51.13 95.28 51.13 95.28 50.87 93.9 50.87 93.9 49.77 95.28 49.77 95.28 49.51 93.9 49.51 93.9 48.41 95.28 48.41 95.28 48.15 93.9 48.15 93.9 47.05 95.28 47.05 95.28 46.79 93.9 46.79 93.9 45.69 95.28 45.69 95.28 45.43 93.9 45.43 93.9 44.33 95.28 44.33 95.28 44.07 93.9 44.07 93.9 42.97 95.28 42.97 95.28 42.71 93.9 42.71 93.9 41.61 95.28 41.61 95.28 41.35 93.9 41.35 93.9 40.25 95.28 40.25 95.28 39.99 93.9 39.99 93.9 38.89 95.28 38.89 95.28 38.63 93.9 38.63 93.9 37.53 95.28 37.53 95.28 35.91 93.9 35.91 93.9 34.81 95.28 34.81 95.28 34.55 93.9 34.55 93.9 33.45 95.28 33.45 95.28 33.19 93.9 33.19 93.9 32.09 95.28 32.09 95.28 31.83 93.9 31.83 93.9 30.73 95.28 30.73 95.28 30.47 93.9 30.47 93.9 29.37 95.28 29.37 95.28 29.11 93.9 29.11 93.9 28.01 95.28 28.01 95.28 27.75 93.9 27.75 93.9 26.65 95.28 26.65 95.28 26.39 93.9 26.39 93.9 25.29 95.28 25.29 95.28 25.03 93.9 25.03 93.9 23.93 95.28 23.93 95.28 23.67 93.9 23.67 93.9 22.57 95.28 22.57 95.28 22.31 93.9 22.31 93.9 21.21 95.28 21.21 95.28 14.15 93.9 14.15 93.9 13.05 95.28 13.05 95.28 12.79 93.9 12.79 93.9 11.69 95.28 11.69 95.28 11.43 93.9 11.43 93.9 10.33 95.28 10.33 95.28 10.07 93.9 10.07 93.9 8.97 95.28 8.97 95.28 7.35 93.9 7.35 93.9 6.25 95.28 6.25 95.28 0.4 0.4 0.4 0.4 97.52 ;
    LAYER met2 ;
      RECT 55.98 97.735 56.26 98.105 ;
      RECT 26.54 97.735 26.82 98.105 ;
      RECT 66.11 96.06 66.37 96.38 ;
      RECT 56.91 96.06 57.17 96.38 ;
      RECT 52.77 96.06 53.03 96.38 ;
      RECT 39.89 96.06 40.15 96.38 ;
      RECT 18.73 96.06 18.99 96.38 ;
      RECT 55.98 -0.185 56.26 0.185 ;
      RECT 26.54 -0.185 26.82 0.185 ;
      POLYGON 67.8 97.64 67.8 86.76 95.4 86.76 95.4 0.28 26.11 0.28 26.11 1.64 25.41 1.64 25.41 0.28 0.28 0.28 0.28 97.64 13.45 97.64 13.45 96.28 14.15 96.28 14.15 97.64 14.37 97.64 14.37 96.28 15.07 96.28 15.07 97.64 15.29 97.64 15.29 96.28 15.99 96.28 15.99 97.64 16.21 97.64 16.21 96.28 16.91 96.28 16.91 97.64 17.13 97.64 17.13 96.28 17.83 96.28 17.83 97.64 18.05 97.64 18.05 96.28 18.75 96.28 18.75 97.64 33.69 97.64 33.69 96.28 34.39 96.28 34.39 97.64 34.61 97.64 34.61 96.28 35.31 96.28 35.31 97.64 35.53 97.64 35.53 96.28 36.23 96.28 36.23 97.64 36.45 97.64 36.45 96.28 37.15 96.28 37.15 97.64 37.37 97.64 37.37 96.28 38.07 96.28 38.07 97.64 38.29 97.64 38.29 96.28 38.99 96.28 38.99 97.64 39.21 97.64 39.21 96.28 39.91 96.28 39.91 97.64 40.13 97.64 40.13 96.28 40.83 96.28 40.83 97.64 41.05 97.64 41.05 96.28 41.75 96.28 41.75 97.64 44.27 97.64 44.27 96.28 44.97 96.28 44.97 97.64 51.17 97.64 51.17 96.28 51.87 96.28 51.87 97.64 52.09 97.64 52.09 96.28 52.79 96.28 52.79 97.64 53.01 97.64 53.01 96.28 53.71 96.28 53.71 97.64 53.93 97.64 53.93 96.28 54.63 96.28 54.63 97.64 54.85 97.64 54.85 96.28 55.55 96.28 55.55 97.64 57.15 97.64 57.15 96.28 57.85 96.28 57.85 97.64 58.07 97.64 58.07 96.28 58.77 96.28 58.77 97.64 58.99 97.64 58.99 96.28 59.69 96.28 59.69 97.64 59.91 97.64 59.91 96.28 60.61 96.28 60.61 97.64 60.83 97.64 60.83 96.28 61.53 96.28 61.53 97.64 61.75 97.64 61.75 96.28 62.45 96.28 62.45 97.64 62.67 97.64 62.67 96.28 63.37 96.28 63.37 97.64 64.05 97.64 64.05 96.28 64.75 96.28 64.75 97.64 65.43 97.64 65.43 96.28 66.13 96.28 66.13 97.64 ;
    LAYER met4 ;
      POLYGON 67.68 97.52 67.68 86.64 84.86 86.64 84.86 86.04 86.26 86.04 86.26 86.64 95.28 86.64 95.28 0.4 86.26 0.4 86.26 1 84.86 1 84.86 0.4 56.82 0.4 56.82 1 55.42 1 55.42 0.4 42.1 0.4 42.1 1 40.7 1 40.7 0.4 27.38 0.4 27.38 1 25.98 1 25.98 0.4 12.66 0.4 12.66 1 11.26 1 11.26 0.4 0.4 0.4 0.4 97.52 11.26 97.52 11.26 96.92 12.66 96.92 12.66 97.52 15.09 97.52 15.09 96.16 16.19 96.16 16.19 97.52 16.93 97.52 16.93 96.16 18.03 96.16 18.03 97.52 25.98 97.52 25.98 96.92 27.38 96.92 27.38 97.52 33.49 97.52 33.49 96.16 34.59 96.16 34.59 97.52 35.33 97.52 35.33 96.16 36.43 96.16 36.43 97.52 37.17 97.52 37.17 96.16 38.27 96.16 38.27 97.52 39.01 97.52 39.01 96.16 40.11 96.16 40.11 97.52 40.7 97.52 40.7 96.92 42.1 96.92 42.1 97.52 53.73 97.52 53.73 96.16 54.83 96.16 54.83 97.52 55.42 97.52 55.42 96.92 56.82 96.92 56.82 97.52 57.41 97.52 57.41 96.16 58.51 96.16 58.51 97.52 59.25 97.52 59.25 96.16 60.35 96.16 60.35 97.52 61.09 97.52 61.09 96.16 62.19 96.16 62.19 97.52 62.93 97.52 62.93 96.16 64.03 96.16 64.03 97.52 ;
    LAYER met5 ;
      POLYGON 66.48 96.32 66.48 85.44 94.08 85.44 94.08 77.32 90.88 77.32 90.88 70.92 94.08 70.92 94.08 56.92 90.88 56.92 90.88 50.52 94.08 50.52 94.08 36.52 90.88 36.52 90.88 30.12 94.08 30.12 94.08 16.12 90.88 16.12 90.88 9.72 94.08 9.72 94.08 1.6 1.6 1.6 1.6 9.72 4.8 9.72 4.8 16.12 1.6 16.12 1.6 30.12 4.8 30.12 4.8 36.52 1.6 36.52 1.6 50.52 4.8 50.52 4.8 56.92 1.6 56.92 1.6 70.92 4.8 70.92 4.8 77.32 1.6 77.32 1.6 96.32 ;
    LAYER met1 ;
      POLYGON 67.8 97.4 67.8 95.72 67.32 95.72 67.32 94.68 67.8 94.68 67.8 93 67.32 93 67.32 91.96 67.8 91.96 67.8 90.28 67.32 90.28 67.32 89.24 67.8 89.24 67.8 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 ;
      POLYGON 95.4 86.52 95.4 84.84 94.92 84.84 94.92 83.8 95.4 83.8 95.4 82.12 94.92 82.12 94.92 81.08 95.4 81.08 95.4 79.4 94.92 79.4 94.92 78.36 95.4 78.36 95.4 76.68 94.92 76.68 94.92 75.64 95.4 75.64 95.4 73.96 94.92 73.96 94.92 72.92 95.4 72.92 95.4 71.24 94.92 71.24 94.92 70.2 95.4 70.2 95.4 68.52 94.92 68.52 94.92 67.48 95.4 67.48 95.4 65.8 94.92 65.8 94.92 64.76 95.4 64.76 95.4 63.08 94.92 63.08 94.92 62.04 95.4 62.04 95.4 60.36 94.92 60.36 94.92 59.32 95.4 59.32 95.4 57.64 94.92 57.64 94.92 56.6 95.4 56.6 95.4 54.92 94.92 54.92 94.92 53.88 95.4 53.88 95.4 52.2 94.92 52.2 94.92 51.16 95.4 51.16 95.4 49.48 94.92 49.48 94.92 48.44 95.4 48.44 95.4 46.76 94.92 46.76 94.92 45.72 95.4 45.72 95.4 44.04 94.92 44.04 94.92 43 95.4 43 95.4 41.32 94.92 41.32 94.92 40.28 95.4 40.28 95.4 38.6 94.92 38.6 94.92 37.56 95.4 37.56 95.4 35.88 94.92 35.88 94.92 34.84 95.4 34.84 95.4 33.16 94.92 33.16 94.92 32.12 95.4 32.12 95.4 30.44 94.92 30.44 94.92 29.4 95.4 29.4 95.4 27.72 94.92 27.72 94.92 26.68 95.4 26.68 95.4 25 94.92 25 94.92 23.96 95.4 23.96 95.4 22.28 94.92 22.28 94.92 21.24 95.4 21.24 95.4 19.56 94.92 19.56 94.92 18.52 95.4 18.52 95.4 16.84 94.92 16.84 94.92 15.8 95.4 15.8 95.4 14.12 94.92 14.12 94.92 13.08 95.4 13.08 95.4 11.4 94.92 11.4 94.92 10.36 95.4 10.36 95.4 8.68 94.92 8.68 94.92 7.64 95.4 7.64 95.4 5.96 94.92 5.96 94.92 4.92 95.4 4.92 95.4 3.24 94.92 3.24 94.92 2.2 95.4 2.2 95.4 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 ;
    LAYER li1 ;
      POLYGON 67.91 97.75 67.91 86.87 95.51 86.87 95.51 0.17 0.17 0.17 0.17 97.75 ;
    LAYER mcon ;
      RECT 67.765 97.835 67.935 98.005 ;
      RECT 67.305 97.835 67.475 98.005 ;
      RECT 66.845 97.835 67.015 98.005 ;
      RECT 66.385 97.835 66.555 98.005 ;
      RECT 65.925 97.835 66.095 98.005 ;
      RECT 65.465 97.835 65.635 98.005 ;
      RECT 65.005 97.835 65.175 98.005 ;
      RECT 64.545 97.835 64.715 98.005 ;
      RECT 64.085 97.835 64.255 98.005 ;
      RECT 63.625 97.835 63.795 98.005 ;
      RECT 63.165 97.835 63.335 98.005 ;
      RECT 62.705 97.835 62.875 98.005 ;
      RECT 62.245 97.835 62.415 98.005 ;
      RECT 61.785 97.835 61.955 98.005 ;
      RECT 61.325 97.835 61.495 98.005 ;
      RECT 60.865 97.835 61.035 98.005 ;
      RECT 60.405 97.835 60.575 98.005 ;
      RECT 59.945 97.835 60.115 98.005 ;
      RECT 59.485 97.835 59.655 98.005 ;
      RECT 59.025 97.835 59.195 98.005 ;
      RECT 58.565 97.835 58.735 98.005 ;
      RECT 58.105 97.835 58.275 98.005 ;
      RECT 57.645 97.835 57.815 98.005 ;
      RECT 57.185 97.835 57.355 98.005 ;
      RECT 56.725 97.835 56.895 98.005 ;
      RECT 56.265 97.835 56.435 98.005 ;
      RECT 55.805 97.835 55.975 98.005 ;
      RECT 55.345 97.835 55.515 98.005 ;
      RECT 54.885 97.835 55.055 98.005 ;
      RECT 54.425 97.835 54.595 98.005 ;
      RECT 53.965 97.835 54.135 98.005 ;
      RECT 53.505 97.835 53.675 98.005 ;
      RECT 53.045 97.835 53.215 98.005 ;
      RECT 52.585 97.835 52.755 98.005 ;
      RECT 52.125 97.835 52.295 98.005 ;
      RECT 51.665 97.835 51.835 98.005 ;
      RECT 51.205 97.835 51.375 98.005 ;
      RECT 50.745 97.835 50.915 98.005 ;
      RECT 50.285 97.835 50.455 98.005 ;
      RECT 49.825 97.835 49.995 98.005 ;
      RECT 49.365 97.835 49.535 98.005 ;
      RECT 48.905 97.835 49.075 98.005 ;
      RECT 48.445 97.835 48.615 98.005 ;
      RECT 47.985 97.835 48.155 98.005 ;
      RECT 47.525 97.835 47.695 98.005 ;
      RECT 47.065 97.835 47.235 98.005 ;
      RECT 46.605 97.835 46.775 98.005 ;
      RECT 46.145 97.835 46.315 98.005 ;
      RECT 45.685 97.835 45.855 98.005 ;
      RECT 45.225 97.835 45.395 98.005 ;
      RECT 44.765 97.835 44.935 98.005 ;
      RECT 44.305 97.835 44.475 98.005 ;
      RECT 43.845 97.835 44.015 98.005 ;
      RECT 43.385 97.835 43.555 98.005 ;
      RECT 42.925 97.835 43.095 98.005 ;
      RECT 42.465 97.835 42.635 98.005 ;
      RECT 42.005 97.835 42.175 98.005 ;
      RECT 41.545 97.835 41.715 98.005 ;
      RECT 41.085 97.835 41.255 98.005 ;
      RECT 40.625 97.835 40.795 98.005 ;
      RECT 40.165 97.835 40.335 98.005 ;
      RECT 39.705 97.835 39.875 98.005 ;
      RECT 39.245 97.835 39.415 98.005 ;
      RECT 38.785 97.835 38.955 98.005 ;
      RECT 38.325 97.835 38.495 98.005 ;
      RECT 37.865 97.835 38.035 98.005 ;
      RECT 37.405 97.835 37.575 98.005 ;
      RECT 36.945 97.835 37.115 98.005 ;
      RECT 36.485 97.835 36.655 98.005 ;
      RECT 36.025 97.835 36.195 98.005 ;
      RECT 35.565 97.835 35.735 98.005 ;
      RECT 35.105 97.835 35.275 98.005 ;
      RECT 34.645 97.835 34.815 98.005 ;
      RECT 34.185 97.835 34.355 98.005 ;
      RECT 33.725 97.835 33.895 98.005 ;
      RECT 33.265 97.835 33.435 98.005 ;
      RECT 32.805 97.835 32.975 98.005 ;
      RECT 32.345 97.835 32.515 98.005 ;
      RECT 31.885 97.835 32.055 98.005 ;
      RECT 31.425 97.835 31.595 98.005 ;
      RECT 30.965 97.835 31.135 98.005 ;
      RECT 30.505 97.835 30.675 98.005 ;
      RECT 30.045 97.835 30.215 98.005 ;
      RECT 29.585 97.835 29.755 98.005 ;
      RECT 29.125 97.835 29.295 98.005 ;
      RECT 28.665 97.835 28.835 98.005 ;
      RECT 28.205 97.835 28.375 98.005 ;
      RECT 27.745 97.835 27.915 98.005 ;
      RECT 27.285 97.835 27.455 98.005 ;
      RECT 26.825 97.835 26.995 98.005 ;
      RECT 26.365 97.835 26.535 98.005 ;
      RECT 25.905 97.835 26.075 98.005 ;
      RECT 25.445 97.835 25.615 98.005 ;
      RECT 24.985 97.835 25.155 98.005 ;
      RECT 24.525 97.835 24.695 98.005 ;
      RECT 24.065 97.835 24.235 98.005 ;
      RECT 23.605 97.835 23.775 98.005 ;
      RECT 23.145 97.835 23.315 98.005 ;
      RECT 22.685 97.835 22.855 98.005 ;
      RECT 22.225 97.835 22.395 98.005 ;
      RECT 21.765 97.835 21.935 98.005 ;
      RECT 21.305 97.835 21.475 98.005 ;
      RECT 20.845 97.835 21.015 98.005 ;
      RECT 20.385 97.835 20.555 98.005 ;
      RECT 19.925 97.835 20.095 98.005 ;
      RECT 19.465 97.835 19.635 98.005 ;
      RECT 19.005 97.835 19.175 98.005 ;
      RECT 18.545 97.835 18.715 98.005 ;
      RECT 18.085 97.835 18.255 98.005 ;
      RECT 17.625 97.835 17.795 98.005 ;
      RECT 17.165 97.835 17.335 98.005 ;
      RECT 16.705 97.835 16.875 98.005 ;
      RECT 16.245 97.835 16.415 98.005 ;
      RECT 15.785 97.835 15.955 98.005 ;
      RECT 15.325 97.835 15.495 98.005 ;
      RECT 14.865 97.835 15.035 98.005 ;
      RECT 14.405 97.835 14.575 98.005 ;
      RECT 13.945 97.835 14.115 98.005 ;
      RECT 13.485 97.835 13.655 98.005 ;
      RECT 13.025 97.835 13.195 98.005 ;
      RECT 12.565 97.835 12.735 98.005 ;
      RECT 12.105 97.835 12.275 98.005 ;
      RECT 11.645 97.835 11.815 98.005 ;
      RECT 11.185 97.835 11.355 98.005 ;
      RECT 10.725 97.835 10.895 98.005 ;
      RECT 10.265 97.835 10.435 98.005 ;
      RECT 9.805 97.835 9.975 98.005 ;
      RECT 9.345 97.835 9.515 98.005 ;
      RECT 8.885 97.835 9.055 98.005 ;
      RECT 8.425 97.835 8.595 98.005 ;
      RECT 7.965 97.835 8.135 98.005 ;
      RECT 7.505 97.835 7.675 98.005 ;
      RECT 7.045 97.835 7.215 98.005 ;
      RECT 6.585 97.835 6.755 98.005 ;
      RECT 6.125 97.835 6.295 98.005 ;
      RECT 5.665 97.835 5.835 98.005 ;
      RECT 5.205 97.835 5.375 98.005 ;
      RECT 4.745 97.835 4.915 98.005 ;
      RECT 4.285 97.835 4.455 98.005 ;
      RECT 3.825 97.835 3.995 98.005 ;
      RECT 3.365 97.835 3.535 98.005 ;
      RECT 2.905 97.835 3.075 98.005 ;
      RECT 2.445 97.835 2.615 98.005 ;
      RECT 1.985 97.835 2.155 98.005 ;
      RECT 1.525 97.835 1.695 98.005 ;
      RECT 1.065 97.835 1.235 98.005 ;
      RECT 0.605 97.835 0.775 98.005 ;
      RECT 0.145 97.835 0.315 98.005 ;
      RECT 67.765 95.115 67.935 95.285 ;
      RECT 67.305 95.115 67.475 95.285 ;
      RECT 0.605 95.115 0.775 95.285 ;
      RECT 0.145 95.115 0.315 95.285 ;
      RECT 67.765 92.395 67.935 92.565 ;
      RECT 67.305 92.395 67.475 92.565 ;
      RECT 0.605 92.395 0.775 92.565 ;
      RECT 0.145 92.395 0.315 92.565 ;
      RECT 67.765 89.675 67.935 89.845 ;
      RECT 67.305 89.675 67.475 89.845 ;
      RECT 0.605 89.675 0.775 89.845 ;
      RECT 0.145 89.675 0.315 89.845 ;
      RECT 95.365 86.955 95.535 87.125 ;
      RECT 94.905 86.955 95.075 87.125 ;
      RECT 94.445 86.955 94.615 87.125 ;
      RECT 93.985 86.955 94.155 87.125 ;
      RECT 93.525 86.955 93.695 87.125 ;
      RECT 93.065 86.955 93.235 87.125 ;
      RECT 92.605 86.955 92.775 87.125 ;
      RECT 92.145 86.955 92.315 87.125 ;
      RECT 91.685 86.955 91.855 87.125 ;
      RECT 91.225 86.955 91.395 87.125 ;
      RECT 90.765 86.955 90.935 87.125 ;
      RECT 90.305 86.955 90.475 87.125 ;
      RECT 89.845 86.955 90.015 87.125 ;
      RECT 89.385 86.955 89.555 87.125 ;
      RECT 88.925 86.955 89.095 87.125 ;
      RECT 88.465 86.955 88.635 87.125 ;
      RECT 88.005 86.955 88.175 87.125 ;
      RECT 87.545 86.955 87.715 87.125 ;
      RECT 87.085 86.955 87.255 87.125 ;
      RECT 86.625 86.955 86.795 87.125 ;
      RECT 86.165 86.955 86.335 87.125 ;
      RECT 85.705 86.955 85.875 87.125 ;
      RECT 85.245 86.955 85.415 87.125 ;
      RECT 84.785 86.955 84.955 87.125 ;
      RECT 84.325 86.955 84.495 87.125 ;
      RECT 83.865 86.955 84.035 87.125 ;
      RECT 83.405 86.955 83.575 87.125 ;
      RECT 82.945 86.955 83.115 87.125 ;
      RECT 82.485 86.955 82.655 87.125 ;
      RECT 82.025 86.955 82.195 87.125 ;
      RECT 81.565 86.955 81.735 87.125 ;
      RECT 81.105 86.955 81.275 87.125 ;
      RECT 80.645 86.955 80.815 87.125 ;
      RECT 80.185 86.955 80.355 87.125 ;
      RECT 79.725 86.955 79.895 87.125 ;
      RECT 79.265 86.955 79.435 87.125 ;
      RECT 78.805 86.955 78.975 87.125 ;
      RECT 78.345 86.955 78.515 87.125 ;
      RECT 77.885 86.955 78.055 87.125 ;
      RECT 77.425 86.955 77.595 87.125 ;
      RECT 76.965 86.955 77.135 87.125 ;
      RECT 76.505 86.955 76.675 87.125 ;
      RECT 76.045 86.955 76.215 87.125 ;
      RECT 75.585 86.955 75.755 87.125 ;
      RECT 75.125 86.955 75.295 87.125 ;
      RECT 74.665 86.955 74.835 87.125 ;
      RECT 74.205 86.955 74.375 87.125 ;
      RECT 73.745 86.955 73.915 87.125 ;
      RECT 73.285 86.955 73.455 87.125 ;
      RECT 72.825 86.955 72.995 87.125 ;
      RECT 72.365 86.955 72.535 87.125 ;
      RECT 71.905 86.955 72.075 87.125 ;
      RECT 71.445 86.955 71.615 87.125 ;
      RECT 70.985 86.955 71.155 87.125 ;
      RECT 70.525 86.955 70.695 87.125 ;
      RECT 70.065 86.955 70.235 87.125 ;
      RECT 69.605 86.955 69.775 87.125 ;
      RECT 69.145 86.955 69.315 87.125 ;
      RECT 68.685 86.955 68.855 87.125 ;
      RECT 68.225 86.955 68.395 87.125 ;
      RECT 67.765 86.955 67.935 87.125 ;
      RECT 67.305 86.955 67.475 87.125 ;
      RECT 66.845 86.955 67.015 87.125 ;
      RECT 66.385 86.955 66.555 87.125 ;
      RECT 65.925 86.955 66.095 87.125 ;
      RECT 65.465 86.955 65.635 87.125 ;
      RECT 65.005 86.955 65.175 87.125 ;
      RECT 64.545 86.955 64.715 87.125 ;
      RECT 64.085 86.955 64.255 87.125 ;
      RECT 63.625 86.955 63.795 87.125 ;
      RECT 63.165 86.955 63.335 87.125 ;
      RECT 62.705 86.955 62.875 87.125 ;
      RECT 62.245 86.955 62.415 87.125 ;
      RECT 61.785 86.955 61.955 87.125 ;
      RECT 61.325 86.955 61.495 87.125 ;
      RECT 60.865 86.955 61.035 87.125 ;
      RECT 60.405 86.955 60.575 87.125 ;
      RECT 59.945 86.955 60.115 87.125 ;
      RECT 59.485 86.955 59.655 87.125 ;
      RECT 59.025 86.955 59.195 87.125 ;
      RECT 58.565 86.955 58.735 87.125 ;
      RECT 58.105 86.955 58.275 87.125 ;
      RECT 57.645 86.955 57.815 87.125 ;
      RECT 57.185 86.955 57.355 87.125 ;
      RECT 56.725 86.955 56.895 87.125 ;
      RECT 56.265 86.955 56.435 87.125 ;
      RECT 55.805 86.955 55.975 87.125 ;
      RECT 55.345 86.955 55.515 87.125 ;
      RECT 54.885 86.955 55.055 87.125 ;
      RECT 54.425 86.955 54.595 87.125 ;
      RECT 53.965 86.955 54.135 87.125 ;
      RECT 53.505 86.955 53.675 87.125 ;
      RECT 53.045 86.955 53.215 87.125 ;
      RECT 52.585 86.955 52.755 87.125 ;
      RECT 52.125 86.955 52.295 87.125 ;
      RECT 51.665 86.955 51.835 87.125 ;
      RECT 51.205 86.955 51.375 87.125 ;
      RECT 50.745 86.955 50.915 87.125 ;
      RECT 50.285 86.955 50.455 87.125 ;
      RECT 49.825 86.955 49.995 87.125 ;
      RECT 49.365 86.955 49.535 87.125 ;
      RECT 48.905 86.955 49.075 87.125 ;
      RECT 48.445 86.955 48.615 87.125 ;
      RECT 47.985 86.955 48.155 87.125 ;
      RECT 47.525 86.955 47.695 87.125 ;
      RECT 47.065 86.955 47.235 87.125 ;
      RECT 46.605 86.955 46.775 87.125 ;
      RECT 46.145 86.955 46.315 87.125 ;
      RECT 45.685 86.955 45.855 87.125 ;
      RECT 45.225 86.955 45.395 87.125 ;
      RECT 44.765 86.955 44.935 87.125 ;
      RECT 44.305 86.955 44.475 87.125 ;
      RECT 43.845 86.955 44.015 87.125 ;
      RECT 43.385 86.955 43.555 87.125 ;
      RECT 42.925 86.955 43.095 87.125 ;
      RECT 42.465 86.955 42.635 87.125 ;
      RECT 42.005 86.955 42.175 87.125 ;
      RECT 41.545 86.955 41.715 87.125 ;
      RECT 41.085 86.955 41.255 87.125 ;
      RECT 40.625 86.955 40.795 87.125 ;
      RECT 40.165 86.955 40.335 87.125 ;
      RECT 39.705 86.955 39.875 87.125 ;
      RECT 39.245 86.955 39.415 87.125 ;
      RECT 38.785 86.955 38.955 87.125 ;
      RECT 38.325 86.955 38.495 87.125 ;
      RECT 37.865 86.955 38.035 87.125 ;
      RECT 37.405 86.955 37.575 87.125 ;
      RECT 36.945 86.955 37.115 87.125 ;
      RECT 36.485 86.955 36.655 87.125 ;
      RECT 36.025 86.955 36.195 87.125 ;
      RECT 35.565 86.955 35.735 87.125 ;
      RECT 35.105 86.955 35.275 87.125 ;
      RECT 34.645 86.955 34.815 87.125 ;
      RECT 34.185 86.955 34.355 87.125 ;
      RECT 33.725 86.955 33.895 87.125 ;
      RECT 33.265 86.955 33.435 87.125 ;
      RECT 32.805 86.955 32.975 87.125 ;
      RECT 32.345 86.955 32.515 87.125 ;
      RECT 31.885 86.955 32.055 87.125 ;
      RECT 31.425 86.955 31.595 87.125 ;
      RECT 30.965 86.955 31.135 87.125 ;
      RECT 30.505 86.955 30.675 87.125 ;
      RECT 30.045 86.955 30.215 87.125 ;
      RECT 29.585 86.955 29.755 87.125 ;
      RECT 29.125 86.955 29.295 87.125 ;
      RECT 28.665 86.955 28.835 87.125 ;
      RECT 28.205 86.955 28.375 87.125 ;
      RECT 27.745 86.955 27.915 87.125 ;
      RECT 27.285 86.955 27.455 87.125 ;
      RECT 26.825 86.955 26.995 87.125 ;
      RECT 26.365 86.955 26.535 87.125 ;
      RECT 25.905 86.955 26.075 87.125 ;
      RECT 25.445 86.955 25.615 87.125 ;
      RECT 24.985 86.955 25.155 87.125 ;
      RECT 24.525 86.955 24.695 87.125 ;
      RECT 24.065 86.955 24.235 87.125 ;
      RECT 23.605 86.955 23.775 87.125 ;
      RECT 23.145 86.955 23.315 87.125 ;
      RECT 22.685 86.955 22.855 87.125 ;
      RECT 22.225 86.955 22.395 87.125 ;
      RECT 21.765 86.955 21.935 87.125 ;
      RECT 21.305 86.955 21.475 87.125 ;
      RECT 20.845 86.955 21.015 87.125 ;
      RECT 20.385 86.955 20.555 87.125 ;
      RECT 19.925 86.955 20.095 87.125 ;
      RECT 19.465 86.955 19.635 87.125 ;
      RECT 19.005 86.955 19.175 87.125 ;
      RECT 18.545 86.955 18.715 87.125 ;
      RECT 18.085 86.955 18.255 87.125 ;
      RECT 17.625 86.955 17.795 87.125 ;
      RECT 17.165 86.955 17.335 87.125 ;
      RECT 16.705 86.955 16.875 87.125 ;
      RECT 16.245 86.955 16.415 87.125 ;
      RECT 15.785 86.955 15.955 87.125 ;
      RECT 15.325 86.955 15.495 87.125 ;
      RECT 14.865 86.955 15.035 87.125 ;
      RECT 14.405 86.955 14.575 87.125 ;
      RECT 13.945 86.955 14.115 87.125 ;
      RECT 13.485 86.955 13.655 87.125 ;
      RECT 13.025 86.955 13.195 87.125 ;
      RECT 12.565 86.955 12.735 87.125 ;
      RECT 12.105 86.955 12.275 87.125 ;
      RECT 11.645 86.955 11.815 87.125 ;
      RECT 11.185 86.955 11.355 87.125 ;
      RECT 10.725 86.955 10.895 87.125 ;
      RECT 10.265 86.955 10.435 87.125 ;
      RECT 9.805 86.955 9.975 87.125 ;
      RECT 9.345 86.955 9.515 87.125 ;
      RECT 8.885 86.955 9.055 87.125 ;
      RECT 8.425 86.955 8.595 87.125 ;
      RECT 7.965 86.955 8.135 87.125 ;
      RECT 7.505 86.955 7.675 87.125 ;
      RECT 7.045 86.955 7.215 87.125 ;
      RECT 6.585 86.955 6.755 87.125 ;
      RECT 6.125 86.955 6.295 87.125 ;
      RECT 5.665 86.955 5.835 87.125 ;
      RECT 5.205 86.955 5.375 87.125 ;
      RECT 4.745 86.955 4.915 87.125 ;
      RECT 4.285 86.955 4.455 87.125 ;
      RECT 3.825 86.955 3.995 87.125 ;
      RECT 3.365 86.955 3.535 87.125 ;
      RECT 2.905 86.955 3.075 87.125 ;
      RECT 2.445 86.955 2.615 87.125 ;
      RECT 1.985 86.955 2.155 87.125 ;
      RECT 1.525 86.955 1.695 87.125 ;
      RECT 1.065 86.955 1.235 87.125 ;
      RECT 0.605 86.955 0.775 87.125 ;
      RECT 0.145 86.955 0.315 87.125 ;
      RECT 95.365 84.235 95.535 84.405 ;
      RECT 94.905 84.235 95.075 84.405 ;
      RECT 0.605 84.235 0.775 84.405 ;
      RECT 0.145 84.235 0.315 84.405 ;
      RECT 95.365 81.515 95.535 81.685 ;
      RECT 94.905 81.515 95.075 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 95.365 78.795 95.535 78.965 ;
      RECT 94.905 78.795 95.075 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 95.365 76.075 95.535 76.245 ;
      RECT 94.905 76.075 95.075 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 95.365 73.355 95.535 73.525 ;
      RECT 94.905 73.355 95.075 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 95.365 70.635 95.535 70.805 ;
      RECT 94.905 70.635 95.075 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 95.365 67.915 95.535 68.085 ;
      RECT 94.905 67.915 95.075 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 95.365 65.195 95.535 65.365 ;
      RECT 94.905 65.195 95.075 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 95.365 62.475 95.535 62.645 ;
      RECT 94.905 62.475 95.075 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 95.365 59.755 95.535 59.925 ;
      RECT 94.905 59.755 95.075 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 95.365 57.035 95.535 57.205 ;
      RECT 94.905 57.035 95.075 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 95.365 54.315 95.535 54.485 ;
      RECT 94.905 54.315 95.075 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 95.365 51.595 95.535 51.765 ;
      RECT 94.905 51.595 95.075 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 95.365 48.875 95.535 49.045 ;
      RECT 94.905 48.875 95.075 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 95.365 46.155 95.535 46.325 ;
      RECT 94.905 46.155 95.075 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 95.365 43.435 95.535 43.605 ;
      RECT 94.905 43.435 95.075 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 95.365 40.715 95.535 40.885 ;
      RECT 94.905 40.715 95.075 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 95.365 37.995 95.535 38.165 ;
      RECT 94.905 37.995 95.075 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 95.365 35.275 95.535 35.445 ;
      RECT 94.905 35.275 95.075 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 95.365 32.555 95.535 32.725 ;
      RECT 94.905 32.555 95.075 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 95.365 29.835 95.535 30.005 ;
      RECT 94.905 29.835 95.075 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 95.365 27.115 95.535 27.285 ;
      RECT 94.905 27.115 95.075 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 95.365 24.395 95.535 24.565 ;
      RECT 94.905 24.395 95.075 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 95.365 21.675 95.535 21.845 ;
      RECT 94.905 21.675 95.075 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 95.365 18.955 95.535 19.125 ;
      RECT 94.905 18.955 95.075 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 95.365 16.235 95.535 16.405 ;
      RECT 94.905 16.235 95.075 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 95.365 13.515 95.535 13.685 ;
      RECT 94.905 13.515 95.075 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 95.365 10.795 95.535 10.965 ;
      RECT 94.905 10.795 95.075 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 95.365 8.075 95.535 8.245 ;
      RECT 94.905 8.075 95.075 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 95.365 5.355 95.535 5.525 ;
      RECT 94.905 5.355 95.075 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 95.365 2.635 95.535 2.805 ;
      RECT 94.905 2.635 95.075 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 95.365 -0.085 95.535 0.085 ;
      RECT 94.905 -0.085 95.075 0.085 ;
      RECT 94.445 -0.085 94.615 0.085 ;
      RECT 93.985 -0.085 94.155 0.085 ;
      RECT 93.525 -0.085 93.695 0.085 ;
      RECT 93.065 -0.085 93.235 0.085 ;
      RECT 92.605 -0.085 92.775 0.085 ;
      RECT 92.145 -0.085 92.315 0.085 ;
      RECT 91.685 -0.085 91.855 0.085 ;
      RECT 91.225 -0.085 91.395 0.085 ;
      RECT 90.765 -0.085 90.935 0.085 ;
      RECT 90.305 -0.085 90.475 0.085 ;
      RECT 89.845 -0.085 90.015 0.085 ;
      RECT 89.385 -0.085 89.555 0.085 ;
      RECT 88.925 -0.085 89.095 0.085 ;
      RECT 88.465 -0.085 88.635 0.085 ;
      RECT 88.005 -0.085 88.175 0.085 ;
      RECT 87.545 -0.085 87.715 0.085 ;
      RECT 87.085 -0.085 87.255 0.085 ;
      RECT 86.625 -0.085 86.795 0.085 ;
      RECT 86.165 -0.085 86.335 0.085 ;
      RECT 85.705 -0.085 85.875 0.085 ;
      RECT 85.245 -0.085 85.415 0.085 ;
      RECT 84.785 -0.085 84.955 0.085 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 56.045 97.845 56.195 97.995 ;
      RECT 26.605 97.845 26.755 97.995 ;
      RECT 55.125 96.145 55.275 96.295 ;
      RECT 44.545 96.145 44.695 96.295 ;
      RECT 36.725 96.145 36.875 96.295 ;
      RECT 56.045 86.965 56.195 87.115 ;
      RECT 26.605 86.965 26.755 87.115 ;
      RECT 56.045 -0.075 56.195 0.075 ;
      RECT 26.605 -0.075 26.755 0.075 ;
    LAYER via2 ;
      RECT 56.02 97.82 56.22 98.02 ;
      RECT 26.58 97.82 26.78 98.02 ;
      RECT 93.74 61.78 93.94 61.98 ;
      RECT 93.74 47.5 93.94 47.7 ;
      RECT 94.2 25.74 94.4 25.94 ;
      RECT 94.2 12.14 94.4 12.34 ;
      RECT 56.02 -0.1 56.22 0.1 ;
      RECT 26.58 -0.1 26.78 0.1 ;
    LAYER via3 ;
      RECT 56.02 97.82 56.22 98.02 ;
      RECT 26.58 97.82 26.78 98.02 ;
      RECT 56.02 -0.1 56.22 0.1 ;
      RECT 26.58 -0.1 26.78 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 97.92 68.08 97.92 68.08 87.04 95.68 87.04 95.68 0 ;
  END
END sb_0__0_

END LIBRARY
