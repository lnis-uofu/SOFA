VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_0__0_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 92 BY 97.92 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 73.53 85.68 73.67 87.04 ;
    END
  END prog_clk[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.55 96.56 44.69 97.92 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.75 96.56 53.89 97.92 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.89 96.56 58.03 97.92 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 96.56 46.53 97.92 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.95 96.56 40.09 97.92 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.53 96.56 27.67 97.92 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.21 96.56 8.35 97.92 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.45 96.56 28.59 97.92 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.37 96.56 29.51 97.92 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.65 96.56 36.95 97.92 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.93 96.56 45.23 97.92 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 96.56 50.21 97.92 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.15 96.56 49.29 97.92 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.97 96.56 57.11 97.92 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.13 96.56 9.27 97.92 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.29 96.56 30.43 97.92 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.51 96.56 33.65 97.92 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.89 96.56 57.19 97.92 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.93 96.56 22.23 97.92 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 96.56 52.97 97.92 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.19 96.56 60.33 97.92 ;
    END
  END top_left_grid_pin_1_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 73.29 92 73.59 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 71.93 92 72.23 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 9.37 92 9.67 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 21.61 92 21.91 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 76.01 92 76.31 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 22.97 92 23.27 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 42.01 92 42.31 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 36.57 92 36.87 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 24.33 92 24.63 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 44.73 92 45.03 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 54.93 92 55.23 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 31.13 92 31.43 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 12.09 92 12.39 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 83.49 92 83.79 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 77.37 92 77.67 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 26.37 92 26.67 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 32.49 92 32.79 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 10.73 92 11.03 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 35.21 92 35.51 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 28.41 92 28.71 ;
    END
  END chanx_right_in[19]
  PIN right_bottom_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 74.65 92 74.95 ;
    END
  END right_bottom_grid_pin_1_[0]
  PIN right_bottom_grid_pin_3_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 59.69 92 59.99 ;
    END
  END right_bottom_grid_pin_3_[0]
  PIN right_bottom_grid_pin_5_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 66.49 92 66.79 ;
    END
  END right_bottom_grid_pin_5_[0]
  PIN right_bottom_grid_pin_7_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 50.17 92 50.47 ;
    END
  END right_bottom_grid_pin_7_[0]
  PIN right_bottom_grid_pin_9_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 61.73 92 62.03 ;
    END
  END right_bottom_grid_pin_9_[0]
  PIN right_bottom_grid_pin_11_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 48.81 92 49.11 ;
    END
  END right_bottom_grid_pin_11_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 13.45 92 13.75 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 96.56 45.61 97.92 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 12.73 96.56 13.03 97.92 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 96.56 47.45 97.92 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 5.37 96.56 5.67 97.92 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.05 96.56 56.19 97.92 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.77 96.56 47.07 97.92 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 34.81 96.56 35.11 97.92 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.77 96.56 24.07 97.92 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.21 96.56 7.51 97.92 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 32.97 96.56 33.27 97.92 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 96.56 48.37 97.92 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.61 96.56 48.91 97.92 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 96.56 51.13 97.92 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 31.13 96.56 31.43 97.92 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 9.05 96.56 9.35 97.92 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 27.45 96.56 27.75 97.92 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 96.56 52.05 97.92 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.29 96.56 52.59 97.92 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 50.45 96.56 50.75 97.92 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.29 96.56 29.59 97.92 ;
    END
  END chany_top_out[19]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 56.97 92 57.27 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 67.85 92 68.15 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 43.37 92 43.67 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 80.09 92 80.39 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 33.85 92 34.15 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 82.13 92 82.43 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 39.29 92 39.59 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 53.57 92 53.87 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 47.45 92 47.75 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 78.73 92 79.03 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 46.09 92 46.39 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 69.21 92 69.51 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 40.65 92 40.95 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 37.93 92 38.23 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 29.77 92 30.07 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 52.21 92 52.51 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 58.33 92 58.63 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 63.09 92 63.39 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 70.57 92 70.87 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.62 65.13 92 65.43 ;
    END
  END chanx_right_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.85 0 23.99 1.36 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 91.52 2.48 92 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 91.52 7.92 92 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 91.52 13.36 92 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 91.52 18.8 92 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 91.52 24.24 92 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 91.52 29.68 92 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 91.52 35.12 92 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 91.52 40.56 92 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 91.52 46 92 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 91.52 51.44 92 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 91.52 56.88 92 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 91.52 62.32 92 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 91.52 67.76 92 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 91.52 73.2 92 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 91.52 78.64 92 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 91.52 84.08 92 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 65.76 89.52 66.24 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 65.76 94.96 66.24 95.44 ;
      LAYER met4 ;
        RECT 10.74 0 11.34 0.6 ;
        RECT 40.18 0 40.78 0.6 ;
        RECT 80.66 0 81.26 0.6 ;
        RECT 80.66 86.44 81.26 87.04 ;
        RECT 10.74 97.32 11.34 97.92 ;
        RECT 40.18 97.32 40.78 97.92 ;
      LAYER met5 ;
        RECT 0 11.32 3.2 14.52 ;
        RECT 88.8 11.32 92 14.52 ;
        RECT 0 52.12 3.2 55.32 ;
        RECT 88.8 52.12 92 55.32 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 0 92 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 91.52 5.2 92 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 91.52 10.64 92 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 91.52 16.08 92 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 91.52 21.52 92 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 91.52 26.96 92 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 91.52 32.4 92 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 91.52 37.84 92 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 91.52 43.28 92 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 91.52 48.72 92 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 91.52 54.16 92 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 91.52 59.6 92 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 91.52 65.04 92 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 91.52 70.48 92 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 91.52 75.92 92 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 91.52 81.36 92 81.84 ;
        RECT 0 86.8 92 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 65.76 92.24 66.24 92.72 ;
        RECT 0 97.68 66.24 97.92 ;
      LAYER met4 ;
        RECT 25.46 0 26.06 0.6 ;
        RECT 54.9 0 55.5 0.6 ;
        RECT 25.46 97.32 26.06 97.92 ;
        RECT 54.9 97.32 55.5 97.92 ;
      LAYER met5 ;
        RECT 0 31.72 3.2 34.92 ;
        RECT 88.8 31.72 92 34.92 ;
        RECT 0 72.52 3.2 75.72 ;
        RECT 88.8 72.52 92 75.72 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 0 97.835 66.24 98.005 ;
      RECT 65.32 95.115 66.24 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 65.32 92.395 66.24 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 65.32 89.675 66.24 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 62.56 86.955 92 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 91.54 84.235 92 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 91.08 81.515 92 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 91.08 78.795 92 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 91.54 76.075 92 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 91.54 73.355 92 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 91.08 70.635 92 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 91.08 67.915 92 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 91.08 65.195 92 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 91.08 62.475 92 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 91.08 59.755 92 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 91.08 57.035 92 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 91.08 54.315 92 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 91.08 51.595 92 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 91.08 48.875 92 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 91.08 46.155 92 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 91.08 43.435 92 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 91.08 40.715 92 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 91.08 37.995 92 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 91.08 35.275 92 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 91.54 32.555 92 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 91.54 29.835 92 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 91.54 27.115 92 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 91.54 24.395 92 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 91.54 21.675 92 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 91.54 18.955 92 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 91.54 16.235 92 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 91.54 13.515 92 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 91.54 10.795 92 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 91.54 8.075 92 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 91.54 5.355 92 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 91.54 2.635 92 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 92 0.085 ;
    LAYER met2 ;
      RECT 55.06 97.735 55.34 98.105 ;
      RECT 25.62 97.735 25.9 98.105 ;
      RECT 55.06 -0.185 55.34 0.185 ;
      RECT 25.62 -0.185 25.9 0.185 ;
      POLYGON 65.96 97.64 65.96 86.76 73.25 86.76 73.25 85.4 73.95 85.4 73.95 86.76 91.72 86.76 91.72 0.28 24.27 0.28 24.27 1.64 23.57 1.64 23.57 0.28 0.28 0.28 0.28 97.64 7.93 97.64 7.93 96.28 8.63 96.28 8.63 97.64 8.85 97.64 8.85 96.28 9.55 96.28 9.55 97.64 27.25 97.64 27.25 96.28 27.95 96.28 27.95 97.64 28.17 97.64 28.17 96.28 28.87 96.28 28.87 97.64 29.09 97.64 29.09 96.28 29.79 96.28 29.79 97.64 30.01 97.64 30.01 96.28 30.71 96.28 30.71 97.64 33.23 97.64 33.23 96.28 33.93 96.28 33.93 97.64 39.67 97.64 39.67 96.28 40.37 96.28 40.37 97.64 44.27 97.64 44.27 96.28 44.97 96.28 44.97 97.64 45.19 97.64 45.19 96.28 45.89 96.28 45.89 97.64 46.11 97.64 46.11 96.28 46.81 96.28 46.81 97.64 47.03 97.64 47.03 96.28 47.73 96.28 47.73 97.64 47.95 97.64 47.95 96.28 48.65 96.28 48.65 97.64 48.87 97.64 48.87 96.28 49.57 96.28 49.57 97.64 49.79 97.64 49.79 96.28 50.49 96.28 50.49 97.64 50.71 97.64 50.71 96.28 51.41 96.28 51.41 97.64 51.63 97.64 51.63 96.28 52.33 96.28 52.33 97.64 52.55 97.64 52.55 96.28 53.25 96.28 53.25 97.64 53.47 97.64 53.47 96.28 54.17 96.28 54.17 97.64 55.77 97.64 55.77 96.28 56.47 96.28 56.47 97.64 56.69 97.64 56.69 96.28 57.39 96.28 57.39 97.64 57.61 97.64 57.61 96.28 58.31 96.28 58.31 97.64 59.91 97.64 59.91 96.28 60.61 96.28 60.61 97.64 ;
    LAYER met4 ;
      POLYGON 65.84 97.52 65.84 86.64 80.26 86.64 80.26 86.04 81.66 86.04 81.66 86.64 91.6 86.64 91.6 0.4 81.66 0.4 81.66 1 80.26 1 80.26 0.4 55.9 0.4 55.9 1 54.5 1 54.5 0.4 41.18 0.4 41.18 1 39.78 1 39.78 0.4 26.46 0.4 26.46 1 25.06 1 25.06 0.4 11.74 0.4 11.74 1 10.34 1 10.34 0.4 0.4 0.4 0.4 97.52 4.97 97.52 4.97 96.16 6.07 96.16 6.07 97.52 6.81 97.52 6.81 96.16 7.91 96.16 7.91 97.52 8.65 97.52 8.65 96.16 9.75 96.16 9.75 97.52 10.34 97.52 10.34 96.92 11.74 96.92 11.74 97.52 12.33 97.52 12.33 96.16 13.43 96.16 13.43 97.52 21.53 97.52 21.53 96.16 22.63 96.16 22.63 97.52 23.37 97.52 23.37 96.16 24.47 96.16 24.47 97.52 25.06 97.52 25.06 96.92 26.46 96.92 26.46 97.52 27.05 97.52 27.05 96.16 28.15 96.16 28.15 97.52 28.89 97.52 28.89 96.16 29.99 96.16 29.99 97.52 30.73 97.52 30.73 96.16 31.83 96.16 31.83 97.52 32.57 97.52 32.57 96.16 33.67 96.16 33.67 97.52 34.41 97.52 34.41 96.16 35.51 96.16 35.51 97.52 36.25 97.52 36.25 96.16 37.35 96.16 37.35 97.52 39.78 97.52 39.78 96.92 41.18 96.92 41.18 97.52 44.53 97.52 44.53 96.16 45.63 96.16 45.63 97.52 46.37 97.52 46.37 96.16 47.47 96.16 47.47 97.52 48.21 97.52 48.21 96.16 49.31 96.16 49.31 97.52 50.05 97.52 50.05 96.16 51.15 96.16 51.15 97.52 51.89 97.52 51.89 96.16 52.99 96.16 52.99 97.52 54.5 97.52 54.5 96.92 55.9 96.92 55.9 97.52 56.49 97.52 56.49 96.16 57.59 96.16 57.59 97.52 ;
    LAYER met3 ;
      POLYGON 55.365 98.085 55.365 98.08 55.58 98.08 55.58 97.76 55.365 97.76 55.365 97.755 55.035 97.755 55.035 97.76 54.82 97.76 54.82 98.08 55.035 98.08 55.035 98.085 ;
      POLYGON 25.925 98.085 25.925 98.08 26.14 98.08 26.14 97.76 25.925 97.76 25.925 97.755 25.595 97.755 25.595 97.76 25.38 97.76 25.38 98.08 25.595 98.08 25.595 98.085 ;
      POLYGON 90.785 56.605 90.785 56.275 90.455 56.275 90.455 56.29 76.67 56.29 76.67 56.59 90.455 56.59 90.455 56.605 ;
      POLYGON 90.77 30.75 90.77 30.47 90.22 30.47 90.22 30.45 72.53 30.45 72.53 30.75 ;
      POLYGON 55.365 0.165 55.365 0.16 55.58 0.16 55.58 -0.16 55.365 -0.16 55.365 -0.165 55.035 -0.165 55.035 -0.16 54.82 -0.16 54.82 0.16 55.035 0.16 55.035 0.165 ;
      POLYGON 25.925 0.165 25.925 0.16 26.14 0.16 26.14 -0.16 25.925 -0.16 25.925 -0.165 25.595 -0.165 25.595 -0.16 25.38 -0.16 25.38 0.16 25.595 0.16 25.595 0.165 ;
      POLYGON 65.84 97.52 65.84 86.64 91.6 86.64 91.6 84.19 90.22 84.19 90.22 83.09 91.6 83.09 91.6 82.83 90.22 82.83 90.22 81.73 91.6 81.73 91.6 80.79 90.22 80.79 90.22 79.69 91.6 79.69 91.6 79.43 90.22 79.43 90.22 78.33 91.6 78.33 91.6 78.07 90.22 78.07 90.22 76.97 91.6 76.97 91.6 76.71 90.22 76.71 90.22 75.61 91.6 75.61 91.6 75.35 90.22 75.35 90.22 74.25 91.6 74.25 91.6 73.99 90.22 73.99 90.22 72.89 91.6 72.89 91.6 72.63 90.22 72.63 90.22 71.53 91.6 71.53 91.6 71.27 90.22 71.27 90.22 70.17 91.6 70.17 91.6 69.91 90.22 69.91 90.22 68.81 91.6 68.81 91.6 68.55 90.22 68.55 90.22 67.45 91.6 67.45 91.6 67.19 90.22 67.19 90.22 66.09 91.6 66.09 91.6 65.83 90.22 65.83 90.22 64.73 91.6 64.73 91.6 63.79 90.22 63.79 90.22 62.69 91.6 62.69 91.6 62.43 90.22 62.43 90.22 61.33 91.6 61.33 91.6 60.39 90.22 60.39 90.22 59.29 91.6 59.29 91.6 59.03 90.22 59.03 90.22 57.93 91.6 57.93 91.6 57.67 90.22 57.67 90.22 56.57 91.6 56.57 91.6 55.63 90.22 55.63 90.22 54.53 91.6 54.53 91.6 54.27 90.22 54.27 90.22 53.17 91.6 53.17 91.6 52.91 90.22 52.91 90.22 51.81 91.6 51.81 91.6 50.87 90.22 50.87 90.22 49.77 91.6 49.77 91.6 49.51 90.22 49.51 90.22 48.41 91.6 48.41 91.6 48.15 90.22 48.15 90.22 47.05 91.6 47.05 91.6 46.79 90.22 46.79 90.22 45.69 91.6 45.69 91.6 45.43 90.22 45.43 90.22 44.33 91.6 44.33 91.6 44.07 90.22 44.07 90.22 42.97 91.6 42.97 91.6 42.71 90.22 42.71 90.22 41.61 91.6 41.61 91.6 41.35 90.22 41.35 90.22 40.25 91.6 40.25 91.6 39.99 90.22 39.99 90.22 38.89 91.6 38.89 91.6 38.63 90.22 38.63 90.22 37.53 91.6 37.53 91.6 37.27 90.22 37.27 90.22 36.17 91.6 36.17 91.6 35.91 90.22 35.91 90.22 34.81 91.6 34.81 91.6 34.55 90.22 34.55 90.22 33.45 91.6 33.45 91.6 33.19 90.22 33.19 90.22 32.09 91.6 32.09 91.6 31.83 90.22 31.83 90.22 30.73 91.6 30.73 91.6 30.47 90.22 30.47 90.22 29.37 91.6 29.37 91.6 29.11 90.22 29.11 90.22 28.01 91.6 28.01 91.6 27.07 90.22 27.07 90.22 25.97 91.6 25.97 91.6 25.03 90.22 25.03 90.22 23.93 91.6 23.93 91.6 23.67 90.22 23.67 90.22 22.57 91.6 22.57 91.6 22.31 90.22 22.31 90.22 21.21 91.6 21.21 91.6 14.15 90.22 14.15 90.22 13.05 91.6 13.05 91.6 12.79 90.22 12.79 90.22 11.69 91.6 11.69 91.6 11.43 90.22 11.43 90.22 10.33 91.6 10.33 91.6 10.07 90.22 10.07 90.22 8.97 91.6 8.97 91.6 0.4 0.4 0.4 0.4 97.52 ;
    LAYER met5 ;
      POLYGON 64.64 96.32 64.64 85.44 90.4 85.44 90.4 77.32 87.2 77.32 87.2 70.92 90.4 70.92 90.4 56.92 87.2 56.92 87.2 50.52 90.4 50.52 90.4 36.52 87.2 36.52 87.2 30.12 90.4 30.12 90.4 16.12 87.2 16.12 87.2 9.72 90.4 9.72 90.4 1.6 1.6 1.6 1.6 9.72 4.8 9.72 4.8 16.12 1.6 16.12 1.6 30.12 4.8 30.12 4.8 36.52 1.6 36.52 1.6 50.52 4.8 50.52 4.8 56.92 1.6 56.92 1.6 70.92 4.8 70.92 4.8 77.32 1.6 77.32 1.6 96.32 ;
    LAYER met1 ;
      POLYGON 65.96 97.4 65.96 95.72 65.48 95.72 65.48 94.68 65.96 94.68 65.96 93 65.48 93 65.48 91.96 65.96 91.96 65.96 90.28 65.48 90.28 65.48 89.24 65.96 89.24 65.96 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 ;
      POLYGON 91.72 86.52 91.72 84.84 91.24 84.84 91.24 83.8 91.72 83.8 91.72 82.12 91.24 82.12 91.24 81.08 91.72 81.08 91.72 79.4 91.24 79.4 91.24 78.36 91.72 78.36 91.72 76.68 91.24 76.68 91.24 75.64 91.72 75.64 91.72 73.96 91.24 73.96 91.24 72.92 91.72 72.92 91.72 71.24 91.24 71.24 91.24 70.2 91.72 70.2 91.72 68.52 91.24 68.52 91.24 67.48 91.72 67.48 91.72 65.8 91.24 65.8 91.24 64.76 91.72 64.76 91.72 63.08 91.24 63.08 91.24 62.04 91.72 62.04 91.72 60.36 91.24 60.36 91.24 59.32 91.72 59.32 91.72 57.64 91.24 57.64 91.24 56.6 91.72 56.6 91.72 54.92 91.24 54.92 91.24 53.88 91.72 53.88 91.72 52.2 91.24 52.2 91.24 51.16 91.72 51.16 91.72 49.48 91.24 49.48 91.24 48.44 91.72 48.44 91.72 46.76 91.24 46.76 91.24 45.72 91.72 45.72 91.72 44.04 91.24 44.04 91.24 43 91.72 43 91.72 41.32 91.24 41.32 91.24 40.28 91.72 40.28 91.72 38.6 91.24 38.6 91.24 37.56 91.72 37.56 91.72 35.88 91.24 35.88 91.24 34.84 91.72 34.84 91.72 33.16 91.24 33.16 91.24 32.12 91.72 32.12 91.72 30.44 91.24 30.44 91.24 29.4 91.72 29.4 91.72 27.72 91.24 27.72 91.24 26.68 91.72 26.68 91.72 25 91.24 25 91.24 23.96 91.72 23.96 91.72 22.28 91.24 22.28 91.24 21.24 91.72 21.24 91.72 19.56 91.24 19.56 91.24 18.52 91.72 18.52 91.72 16.84 91.24 16.84 91.24 15.8 91.72 15.8 91.72 14.12 91.24 14.12 91.24 13.08 91.72 13.08 91.72 11.4 91.24 11.4 91.24 10.36 91.72 10.36 91.72 8.68 91.24 8.68 91.24 7.64 91.72 7.64 91.72 5.96 91.24 5.96 91.24 4.92 91.72 4.92 91.72 3.24 91.24 3.24 91.24 2.2 91.72 2.2 91.72 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 ;
    LAYER li1 ;
      POLYGON 66.07 97.75 66.07 86.87 91.83 86.87 91.83 0.17 0.17 0.17 0.17 97.75 ;
    LAYER mcon ;
      RECT 65.925 97.835 66.095 98.005 ;
      RECT 65.465 97.835 65.635 98.005 ;
      RECT 65.005 97.835 65.175 98.005 ;
      RECT 64.545 97.835 64.715 98.005 ;
      RECT 64.085 97.835 64.255 98.005 ;
      RECT 63.625 97.835 63.795 98.005 ;
      RECT 63.165 97.835 63.335 98.005 ;
      RECT 62.705 97.835 62.875 98.005 ;
      RECT 62.245 97.835 62.415 98.005 ;
      RECT 61.785 97.835 61.955 98.005 ;
      RECT 61.325 97.835 61.495 98.005 ;
      RECT 60.865 97.835 61.035 98.005 ;
      RECT 60.405 97.835 60.575 98.005 ;
      RECT 59.945 97.835 60.115 98.005 ;
      RECT 59.485 97.835 59.655 98.005 ;
      RECT 59.025 97.835 59.195 98.005 ;
      RECT 58.565 97.835 58.735 98.005 ;
      RECT 58.105 97.835 58.275 98.005 ;
      RECT 57.645 97.835 57.815 98.005 ;
      RECT 57.185 97.835 57.355 98.005 ;
      RECT 56.725 97.835 56.895 98.005 ;
      RECT 56.265 97.835 56.435 98.005 ;
      RECT 55.805 97.835 55.975 98.005 ;
      RECT 55.345 97.835 55.515 98.005 ;
      RECT 54.885 97.835 55.055 98.005 ;
      RECT 54.425 97.835 54.595 98.005 ;
      RECT 53.965 97.835 54.135 98.005 ;
      RECT 53.505 97.835 53.675 98.005 ;
      RECT 53.045 97.835 53.215 98.005 ;
      RECT 52.585 97.835 52.755 98.005 ;
      RECT 52.125 97.835 52.295 98.005 ;
      RECT 51.665 97.835 51.835 98.005 ;
      RECT 51.205 97.835 51.375 98.005 ;
      RECT 50.745 97.835 50.915 98.005 ;
      RECT 50.285 97.835 50.455 98.005 ;
      RECT 49.825 97.835 49.995 98.005 ;
      RECT 49.365 97.835 49.535 98.005 ;
      RECT 48.905 97.835 49.075 98.005 ;
      RECT 48.445 97.835 48.615 98.005 ;
      RECT 47.985 97.835 48.155 98.005 ;
      RECT 47.525 97.835 47.695 98.005 ;
      RECT 47.065 97.835 47.235 98.005 ;
      RECT 46.605 97.835 46.775 98.005 ;
      RECT 46.145 97.835 46.315 98.005 ;
      RECT 45.685 97.835 45.855 98.005 ;
      RECT 45.225 97.835 45.395 98.005 ;
      RECT 44.765 97.835 44.935 98.005 ;
      RECT 44.305 97.835 44.475 98.005 ;
      RECT 43.845 97.835 44.015 98.005 ;
      RECT 43.385 97.835 43.555 98.005 ;
      RECT 42.925 97.835 43.095 98.005 ;
      RECT 42.465 97.835 42.635 98.005 ;
      RECT 42.005 97.835 42.175 98.005 ;
      RECT 41.545 97.835 41.715 98.005 ;
      RECT 41.085 97.835 41.255 98.005 ;
      RECT 40.625 97.835 40.795 98.005 ;
      RECT 40.165 97.835 40.335 98.005 ;
      RECT 39.705 97.835 39.875 98.005 ;
      RECT 39.245 97.835 39.415 98.005 ;
      RECT 38.785 97.835 38.955 98.005 ;
      RECT 38.325 97.835 38.495 98.005 ;
      RECT 37.865 97.835 38.035 98.005 ;
      RECT 37.405 97.835 37.575 98.005 ;
      RECT 36.945 97.835 37.115 98.005 ;
      RECT 36.485 97.835 36.655 98.005 ;
      RECT 36.025 97.835 36.195 98.005 ;
      RECT 35.565 97.835 35.735 98.005 ;
      RECT 35.105 97.835 35.275 98.005 ;
      RECT 34.645 97.835 34.815 98.005 ;
      RECT 34.185 97.835 34.355 98.005 ;
      RECT 33.725 97.835 33.895 98.005 ;
      RECT 33.265 97.835 33.435 98.005 ;
      RECT 32.805 97.835 32.975 98.005 ;
      RECT 32.345 97.835 32.515 98.005 ;
      RECT 31.885 97.835 32.055 98.005 ;
      RECT 31.425 97.835 31.595 98.005 ;
      RECT 30.965 97.835 31.135 98.005 ;
      RECT 30.505 97.835 30.675 98.005 ;
      RECT 30.045 97.835 30.215 98.005 ;
      RECT 29.585 97.835 29.755 98.005 ;
      RECT 29.125 97.835 29.295 98.005 ;
      RECT 28.665 97.835 28.835 98.005 ;
      RECT 28.205 97.835 28.375 98.005 ;
      RECT 27.745 97.835 27.915 98.005 ;
      RECT 27.285 97.835 27.455 98.005 ;
      RECT 26.825 97.835 26.995 98.005 ;
      RECT 26.365 97.835 26.535 98.005 ;
      RECT 25.905 97.835 26.075 98.005 ;
      RECT 25.445 97.835 25.615 98.005 ;
      RECT 24.985 97.835 25.155 98.005 ;
      RECT 24.525 97.835 24.695 98.005 ;
      RECT 24.065 97.835 24.235 98.005 ;
      RECT 23.605 97.835 23.775 98.005 ;
      RECT 23.145 97.835 23.315 98.005 ;
      RECT 22.685 97.835 22.855 98.005 ;
      RECT 22.225 97.835 22.395 98.005 ;
      RECT 21.765 97.835 21.935 98.005 ;
      RECT 21.305 97.835 21.475 98.005 ;
      RECT 20.845 97.835 21.015 98.005 ;
      RECT 20.385 97.835 20.555 98.005 ;
      RECT 19.925 97.835 20.095 98.005 ;
      RECT 19.465 97.835 19.635 98.005 ;
      RECT 19.005 97.835 19.175 98.005 ;
      RECT 18.545 97.835 18.715 98.005 ;
      RECT 18.085 97.835 18.255 98.005 ;
      RECT 17.625 97.835 17.795 98.005 ;
      RECT 17.165 97.835 17.335 98.005 ;
      RECT 16.705 97.835 16.875 98.005 ;
      RECT 16.245 97.835 16.415 98.005 ;
      RECT 15.785 97.835 15.955 98.005 ;
      RECT 15.325 97.835 15.495 98.005 ;
      RECT 14.865 97.835 15.035 98.005 ;
      RECT 14.405 97.835 14.575 98.005 ;
      RECT 13.945 97.835 14.115 98.005 ;
      RECT 13.485 97.835 13.655 98.005 ;
      RECT 13.025 97.835 13.195 98.005 ;
      RECT 12.565 97.835 12.735 98.005 ;
      RECT 12.105 97.835 12.275 98.005 ;
      RECT 11.645 97.835 11.815 98.005 ;
      RECT 11.185 97.835 11.355 98.005 ;
      RECT 10.725 97.835 10.895 98.005 ;
      RECT 10.265 97.835 10.435 98.005 ;
      RECT 9.805 97.835 9.975 98.005 ;
      RECT 9.345 97.835 9.515 98.005 ;
      RECT 8.885 97.835 9.055 98.005 ;
      RECT 8.425 97.835 8.595 98.005 ;
      RECT 7.965 97.835 8.135 98.005 ;
      RECT 7.505 97.835 7.675 98.005 ;
      RECT 7.045 97.835 7.215 98.005 ;
      RECT 6.585 97.835 6.755 98.005 ;
      RECT 6.125 97.835 6.295 98.005 ;
      RECT 5.665 97.835 5.835 98.005 ;
      RECT 5.205 97.835 5.375 98.005 ;
      RECT 4.745 97.835 4.915 98.005 ;
      RECT 4.285 97.835 4.455 98.005 ;
      RECT 3.825 97.835 3.995 98.005 ;
      RECT 3.365 97.835 3.535 98.005 ;
      RECT 2.905 97.835 3.075 98.005 ;
      RECT 2.445 97.835 2.615 98.005 ;
      RECT 1.985 97.835 2.155 98.005 ;
      RECT 1.525 97.835 1.695 98.005 ;
      RECT 1.065 97.835 1.235 98.005 ;
      RECT 0.605 97.835 0.775 98.005 ;
      RECT 0.145 97.835 0.315 98.005 ;
      RECT 65.925 95.115 66.095 95.285 ;
      RECT 65.465 95.115 65.635 95.285 ;
      RECT 0.605 95.115 0.775 95.285 ;
      RECT 0.145 95.115 0.315 95.285 ;
      RECT 65.925 92.395 66.095 92.565 ;
      RECT 65.465 92.395 65.635 92.565 ;
      RECT 0.605 92.395 0.775 92.565 ;
      RECT 0.145 92.395 0.315 92.565 ;
      RECT 65.925 89.675 66.095 89.845 ;
      RECT 65.465 89.675 65.635 89.845 ;
      RECT 0.605 89.675 0.775 89.845 ;
      RECT 0.145 89.675 0.315 89.845 ;
      RECT 91.685 86.955 91.855 87.125 ;
      RECT 91.225 86.955 91.395 87.125 ;
      RECT 90.765 86.955 90.935 87.125 ;
      RECT 90.305 86.955 90.475 87.125 ;
      RECT 89.845 86.955 90.015 87.125 ;
      RECT 89.385 86.955 89.555 87.125 ;
      RECT 88.925 86.955 89.095 87.125 ;
      RECT 88.465 86.955 88.635 87.125 ;
      RECT 88.005 86.955 88.175 87.125 ;
      RECT 87.545 86.955 87.715 87.125 ;
      RECT 87.085 86.955 87.255 87.125 ;
      RECT 86.625 86.955 86.795 87.125 ;
      RECT 86.165 86.955 86.335 87.125 ;
      RECT 85.705 86.955 85.875 87.125 ;
      RECT 85.245 86.955 85.415 87.125 ;
      RECT 84.785 86.955 84.955 87.125 ;
      RECT 84.325 86.955 84.495 87.125 ;
      RECT 83.865 86.955 84.035 87.125 ;
      RECT 83.405 86.955 83.575 87.125 ;
      RECT 82.945 86.955 83.115 87.125 ;
      RECT 82.485 86.955 82.655 87.125 ;
      RECT 82.025 86.955 82.195 87.125 ;
      RECT 81.565 86.955 81.735 87.125 ;
      RECT 81.105 86.955 81.275 87.125 ;
      RECT 80.645 86.955 80.815 87.125 ;
      RECT 80.185 86.955 80.355 87.125 ;
      RECT 79.725 86.955 79.895 87.125 ;
      RECT 79.265 86.955 79.435 87.125 ;
      RECT 78.805 86.955 78.975 87.125 ;
      RECT 78.345 86.955 78.515 87.125 ;
      RECT 77.885 86.955 78.055 87.125 ;
      RECT 77.425 86.955 77.595 87.125 ;
      RECT 76.965 86.955 77.135 87.125 ;
      RECT 76.505 86.955 76.675 87.125 ;
      RECT 76.045 86.955 76.215 87.125 ;
      RECT 75.585 86.955 75.755 87.125 ;
      RECT 75.125 86.955 75.295 87.125 ;
      RECT 74.665 86.955 74.835 87.125 ;
      RECT 74.205 86.955 74.375 87.125 ;
      RECT 73.745 86.955 73.915 87.125 ;
      RECT 73.285 86.955 73.455 87.125 ;
      RECT 72.825 86.955 72.995 87.125 ;
      RECT 72.365 86.955 72.535 87.125 ;
      RECT 71.905 86.955 72.075 87.125 ;
      RECT 71.445 86.955 71.615 87.125 ;
      RECT 70.985 86.955 71.155 87.125 ;
      RECT 70.525 86.955 70.695 87.125 ;
      RECT 70.065 86.955 70.235 87.125 ;
      RECT 69.605 86.955 69.775 87.125 ;
      RECT 69.145 86.955 69.315 87.125 ;
      RECT 68.685 86.955 68.855 87.125 ;
      RECT 68.225 86.955 68.395 87.125 ;
      RECT 67.765 86.955 67.935 87.125 ;
      RECT 67.305 86.955 67.475 87.125 ;
      RECT 66.845 86.955 67.015 87.125 ;
      RECT 66.385 86.955 66.555 87.125 ;
      RECT 65.925 86.955 66.095 87.125 ;
      RECT 65.465 86.955 65.635 87.125 ;
      RECT 65.005 86.955 65.175 87.125 ;
      RECT 64.545 86.955 64.715 87.125 ;
      RECT 64.085 86.955 64.255 87.125 ;
      RECT 63.625 86.955 63.795 87.125 ;
      RECT 63.165 86.955 63.335 87.125 ;
      RECT 62.705 86.955 62.875 87.125 ;
      RECT 62.245 86.955 62.415 87.125 ;
      RECT 61.785 86.955 61.955 87.125 ;
      RECT 61.325 86.955 61.495 87.125 ;
      RECT 60.865 86.955 61.035 87.125 ;
      RECT 60.405 86.955 60.575 87.125 ;
      RECT 59.945 86.955 60.115 87.125 ;
      RECT 59.485 86.955 59.655 87.125 ;
      RECT 59.025 86.955 59.195 87.125 ;
      RECT 58.565 86.955 58.735 87.125 ;
      RECT 58.105 86.955 58.275 87.125 ;
      RECT 57.645 86.955 57.815 87.125 ;
      RECT 57.185 86.955 57.355 87.125 ;
      RECT 56.725 86.955 56.895 87.125 ;
      RECT 56.265 86.955 56.435 87.125 ;
      RECT 55.805 86.955 55.975 87.125 ;
      RECT 55.345 86.955 55.515 87.125 ;
      RECT 54.885 86.955 55.055 87.125 ;
      RECT 54.425 86.955 54.595 87.125 ;
      RECT 53.965 86.955 54.135 87.125 ;
      RECT 53.505 86.955 53.675 87.125 ;
      RECT 53.045 86.955 53.215 87.125 ;
      RECT 52.585 86.955 52.755 87.125 ;
      RECT 52.125 86.955 52.295 87.125 ;
      RECT 51.665 86.955 51.835 87.125 ;
      RECT 51.205 86.955 51.375 87.125 ;
      RECT 50.745 86.955 50.915 87.125 ;
      RECT 50.285 86.955 50.455 87.125 ;
      RECT 49.825 86.955 49.995 87.125 ;
      RECT 49.365 86.955 49.535 87.125 ;
      RECT 48.905 86.955 49.075 87.125 ;
      RECT 48.445 86.955 48.615 87.125 ;
      RECT 47.985 86.955 48.155 87.125 ;
      RECT 47.525 86.955 47.695 87.125 ;
      RECT 47.065 86.955 47.235 87.125 ;
      RECT 46.605 86.955 46.775 87.125 ;
      RECT 46.145 86.955 46.315 87.125 ;
      RECT 45.685 86.955 45.855 87.125 ;
      RECT 45.225 86.955 45.395 87.125 ;
      RECT 44.765 86.955 44.935 87.125 ;
      RECT 44.305 86.955 44.475 87.125 ;
      RECT 43.845 86.955 44.015 87.125 ;
      RECT 43.385 86.955 43.555 87.125 ;
      RECT 42.925 86.955 43.095 87.125 ;
      RECT 42.465 86.955 42.635 87.125 ;
      RECT 42.005 86.955 42.175 87.125 ;
      RECT 41.545 86.955 41.715 87.125 ;
      RECT 41.085 86.955 41.255 87.125 ;
      RECT 40.625 86.955 40.795 87.125 ;
      RECT 40.165 86.955 40.335 87.125 ;
      RECT 39.705 86.955 39.875 87.125 ;
      RECT 39.245 86.955 39.415 87.125 ;
      RECT 38.785 86.955 38.955 87.125 ;
      RECT 38.325 86.955 38.495 87.125 ;
      RECT 37.865 86.955 38.035 87.125 ;
      RECT 37.405 86.955 37.575 87.125 ;
      RECT 36.945 86.955 37.115 87.125 ;
      RECT 36.485 86.955 36.655 87.125 ;
      RECT 36.025 86.955 36.195 87.125 ;
      RECT 35.565 86.955 35.735 87.125 ;
      RECT 35.105 86.955 35.275 87.125 ;
      RECT 34.645 86.955 34.815 87.125 ;
      RECT 34.185 86.955 34.355 87.125 ;
      RECT 33.725 86.955 33.895 87.125 ;
      RECT 33.265 86.955 33.435 87.125 ;
      RECT 32.805 86.955 32.975 87.125 ;
      RECT 32.345 86.955 32.515 87.125 ;
      RECT 31.885 86.955 32.055 87.125 ;
      RECT 31.425 86.955 31.595 87.125 ;
      RECT 30.965 86.955 31.135 87.125 ;
      RECT 30.505 86.955 30.675 87.125 ;
      RECT 30.045 86.955 30.215 87.125 ;
      RECT 29.585 86.955 29.755 87.125 ;
      RECT 29.125 86.955 29.295 87.125 ;
      RECT 28.665 86.955 28.835 87.125 ;
      RECT 28.205 86.955 28.375 87.125 ;
      RECT 27.745 86.955 27.915 87.125 ;
      RECT 27.285 86.955 27.455 87.125 ;
      RECT 26.825 86.955 26.995 87.125 ;
      RECT 26.365 86.955 26.535 87.125 ;
      RECT 25.905 86.955 26.075 87.125 ;
      RECT 25.445 86.955 25.615 87.125 ;
      RECT 24.985 86.955 25.155 87.125 ;
      RECT 24.525 86.955 24.695 87.125 ;
      RECT 24.065 86.955 24.235 87.125 ;
      RECT 23.605 86.955 23.775 87.125 ;
      RECT 23.145 86.955 23.315 87.125 ;
      RECT 22.685 86.955 22.855 87.125 ;
      RECT 22.225 86.955 22.395 87.125 ;
      RECT 21.765 86.955 21.935 87.125 ;
      RECT 21.305 86.955 21.475 87.125 ;
      RECT 20.845 86.955 21.015 87.125 ;
      RECT 20.385 86.955 20.555 87.125 ;
      RECT 19.925 86.955 20.095 87.125 ;
      RECT 19.465 86.955 19.635 87.125 ;
      RECT 19.005 86.955 19.175 87.125 ;
      RECT 18.545 86.955 18.715 87.125 ;
      RECT 18.085 86.955 18.255 87.125 ;
      RECT 17.625 86.955 17.795 87.125 ;
      RECT 17.165 86.955 17.335 87.125 ;
      RECT 16.705 86.955 16.875 87.125 ;
      RECT 16.245 86.955 16.415 87.125 ;
      RECT 15.785 86.955 15.955 87.125 ;
      RECT 15.325 86.955 15.495 87.125 ;
      RECT 14.865 86.955 15.035 87.125 ;
      RECT 14.405 86.955 14.575 87.125 ;
      RECT 13.945 86.955 14.115 87.125 ;
      RECT 13.485 86.955 13.655 87.125 ;
      RECT 13.025 86.955 13.195 87.125 ;
      RECT 12.565 86.955 12.735 87.125 ;
      RECT 12.105 86.955 12.275 87.125 ;
      RECT 11.645 86.955 11.815 87.125 ;
      RECT 11.185 86.955 11.355 87.125 ;
      RECT 10.725 86.955 10.895 87.125 ;
      RECT 10.265 86.955 10.435 87.125 ;
      RECT 9.805 86.955 9.975 87.125 ;
      RECT 9.345 86.955 9.515 87.125 ;
      RECT 8.885 86.955 9.055 87.125 ;
      RECT 8.425 86.955 8.595 87.125 ;
      RECT 7.965 86.955 8.135 87.125 ;
      RECT 7.505 86.955 7.675 87.125 ;
      RECT 7.045 86.955 7.215 87.125 ;
      RECT 6.585 86.955 6.755 87.125 ;
      RECT 6.125 86.955 6.295 87.125 ;
      RECT 5.665 86.955 5.835 87.125 ;
      RECT 5.205 86.955 5.375 87.125 ;
      RECT 4.745 86.955 4.915 87.125 ;
      RECT 4.285 86.955 4.455 87.125 ;
      RECT 3.825 86.955 3.995 87.125 ;
      RECT 3.365 86.955 3.535 87.125 ;
      RECT 2.905 86.955 3.075 87.125 ;
      RECT 2.445 86.955 2.615 87.125 ;
      RECT 1.985 86.955 2.155 87.125 ;
      RECT 1.525 86.955 1.695 87.125 ;
      RECT 1.065 86.955 1.235 87.125 ;
      RECT 0.605 86.955 0.775 87.125 ;
      RECT 0.145 86.955 0.315 87.125 ;
      RECT 91.685 84.235 91.855 84.405 ;
      RECT 91.225 84.235 91.395 84.405 ;
      RECT 0.605 84.235 0.775 84.405 ;
      RECT 0.145 84.235 0.315 84.405 ;
      RECT 91.685 81.515 91.855 81.685 ;
      RECT 91.225 81.515 91.395 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 91.685 78.795 91.855 78.965 ;
      RECT 91.225 78.795 91.395 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 91.685 76.075 91.855 76.245 ;
      RECT 91.225 76.075 91.395 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 91.685 73.355 91.855 73.525 ;
      RECT 91.225 73.355 91.395 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 91.685 70.635 91.855 70.805 ;
      RECT 91.225 70.635 91.395 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 91.685 67.915 91.855 68.085 ;
      RECT 91.225 67.915 91.395 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 91.685 65.195 91.855 65.365 ;
      RECT 91.225 65.195 91.395 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 91.685 62.475 91.855 62.645 ;
      RECT 91.225 62.475 91.395 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 91.685 59.755 91.855 59.925 ;
      RECT 91.225 59.755 91.395 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 91.685 57.035 91.855 57.205 ;
      RECT 91.225 57.035 91.395 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 91.685 54.315 91.855 54.485 ;
      RECT 91.225 54.315 91.395 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 91.685 51.595 91.855 51.765 ;
      RECT 91.225 51.595 91.395 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 91.685 48.875 91.855 49.045 ;
      RECT 91.225 48.875 91.395 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 91.685 46.155 91.855 46.325 ;
      RECT 91.225 46.155 91.395 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 91.685 43.435 91.855 43.605 ;
      RECT 91.225 43.435 91.395 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 91.685 40.715 91.855 40.885 ;
      RECT 91.225 40.715 91.395 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 91.685 37.995 91.855 38.165 ;
      RECT 91.225 37.995 91.395 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 91.685 35.275 91.855 35.445 ;
      RECT 91.225 35.275 91.395 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 91.685 32.555 91.855 32.725 ;
      RECT 91.225 32.555 91.395 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 91.685 29.835 91.855 30.005 ;
      RECT 91.225 29.835 91.395 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 91.685 27.115 91.855 27.285 ;
      RECT 91.225 27.115 91.395 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 91.685 24.395 91.855 24.565 ;
      RECT 91.225 24.395 91.395 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 91.685 21.675 91.855 21.845 ;
      RECT 91.225 21.675 91.395 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 91.685 18.955 91.855 19.125 ;
      RECT 91.225 18.955 91.395 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 91.685 16.235 91.855 16.405 ;
      RECT 91.225 16.235 91.395 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 91.685 13.515 91.855 13.685 ;
      RECT 91.225 13.515 91.395 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 91.685 10.795 91.855 10.965 ;
      RECT 91.225 10.795 91.395 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 91.685 8.075 91.855 8.245 ;
      RECT 91.225 8.075 91.395 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 91.685 5.355 91.855 5.525 ;
      RECT 91.225 5.355 91.395 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 91.685 2.635 91.855 2.805 ;
      RECT 91.225 2.635 91.395 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 91.685 -0.085 91.855 0.085 ;
      RECT 91.225 -0.085 91.395 0.085 ;
      RECT 90.765 -0.085 90.935 0.085 ;
      RECT 90.305 -0.085 90.475 0.085 ;
      RECT 89.845 -0.085 90.015 0.085 ;
      RECT 89.385 -0.085 89.555 0.085 ;
      RECT 88.925 -0.085 89.095 0.085 ;
      RECT 88.465 -0.085 88.635 0.085 ;
      RECT 88.005 -0.085 88.175 0.085 ;
      RECT 87.545 -0.085 87.715 0.085 ;
      RECT 87.085 -0.085 87.255 0.085 ;
      RECT 86.625 -0.085 86.795 0.085 ;
      RECT 86.165 -0.085 86.335 0.085 ;
      RECT 85.705 -0.085 85.875 0.085 ;
      RECT 85.245 -0.085 85.415 0.085 ;
      RECT 84.785 -0.085 84.955 0.085 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 55.125 97.845 55.275 97.995 ;
      RECT 25.685 97.845 25.835 97.995 ;
      RECT 46.385 96.145 46.535 96.295 ;
      RECT 29.365 96.145 29.515 96.295 ;
      RECT 55.125 86.965 55.275 87.115 ;
      RECT 25.685 86.965 25.835 87.115 ;
      RECT 55.125 -0.075 55.275 0.075 ;
      RECT 25.685 -0.075 25.835 0.075 ;
    LAYER via2 ;
      RECT 55.1 97.82 55.3 98.02 ;
      RECT 25.66 97.82 25.86 98.02 ;
      RECT 90.52 78.78 90.72 78.98 ;
      RECT 90.52 70.62 90.72 70.82 ;
      RECT 90.52 61.78 90.72 61.98 ;
      RECT 90.52 52.26 90.72 52.46 ;
      RECT 90.52 46.14 90.72 46.34 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER via3 ;
      RECT 55.1 97.82 55.3 98.02 ;
      RECT 25.66 97.82 25.86 98.02 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 97.92 66.24 97.92 66.24 87.04 92 87.04 92 0 ;
  END
END sb_0__0_

END LIBRARY
