VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_2__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 92 BY 108.8 ;
  SYMMETRY X Y ;
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.74 108.315 56.88 108.8 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.04 108.315 59.18 108.8 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 108.315 65.16 108.8 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.08 108.315 70.22 108.8 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.18 108.315 63.32 108.8 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.78 108.315 67.92 108.8 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.14 108.315 52.28 108.8 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.06 108.315 53.2 108.8 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.7 108.315 45.84 108.8 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.94 108.315 66.08 108.8 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 108.315 64.24 108.8 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.68 108.315 74.82 108.8 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 108.315 62.4 108.8 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.84 108.315 72.98 108.8 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.98 108.315 54.12 108.8 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.12 108.315 58.26 108.8 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.46 108.315 48.6 108.8 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.76 108.315 73.9 108.8 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.78 108.315 44.92 108.8 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.16 108.315 69.3 108.8 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.5 97.435 13.64 97.92 ;
    END
  END top_left_grid_pin_42_[0]
  PIN top_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.66 97.435 11.8 97.92 ;
    END
  END top_left_grid_pin_43_[0]
  PIN top_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.44 97.435 8.58 97.92 ;
    END
  END top_left_grid_pin_44_[0]
  PIN top_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.58 97.435 12.72 97.92 ;
    END
  END top_left_grid_pin_45_[0]
  PIN top_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.28 97.435 10.42 97.92 ;
    END
  END top_left_grid_pin_46_[0]
  PIN top_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.3 97.435 4.44 97.92 ;
    END
  END top_left_grid_pin_47_[0]
  PIN top_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.36 97.435 9.5 97.92 ;
    END
  END top_left_grid_pin_48_[0]
  PIN top_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.06 97.435 7.2 97.92 ;
    END
  END top_left_grid_pin_49_[0]
  PIN top_right_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.44 108.315 31.58 108.8 ;
    END
  END top_right_grid_pin_1_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.08 0 70.22 0.485 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.58 0 81.72 0.485 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.2 0 57.34 0.485 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.2 0 80.34 0.485 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.56 0 64.7 0.485 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.52 0 76.66 0.485 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.36 0 55.5 0.485 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.76 0 73.9 0.485 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.64 0 63.78 0.485 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.16 0 69.3 0.485 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.14 0 52.28 0.485 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71 0 71.14 0.485 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.6 0 75.74 0.485 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.36 0 78.5 0.485 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.44 0 54.58 0.485 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.4 0 66.54 0.485 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.08 0 47.22 0.485 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.44 0 77.58 0.485 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.06 0 53.2 0.485 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.28 0 79.42 0.485 ;
    END
  END chany_bottom_in[19]
  PIN bottom_right_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.36 0 32.5 0.485 ;
    END
  END bottom_right_grid_pin_1_[0]
  PIN bottom_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.42 10.88 14.56 11.365 ;
    END
  END bottom_left_grid_pin_42_[0]
  PIN bottom_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.34 10.88 15.48 11.365 ;
    END
  END bottom_left_grid_pin_43_[0]
  PIN bottom_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.92 10.88 3.06 11.365 ;
    END
  END bottom_left_grid_pin_44_[0]
  PIN bottom_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.28 10.88 10.42 11.365 ;
    END
  END bottom_left_grid_pin_45_[0]
  PIN bottom_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.22 10.88 5.36 11.365 ;
    END
  END bottom_left_grid_pin_46_[0]
  PIN bottom_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.3 10.88 4.44 11.365 ;
    END
  END bottom_left_grid_pin_47_[0]
  PIN bottom_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.5 10.88 13.64 11.365 ;
    END
  END bottom_left_grid_pin_48_[0]
  PIN bottom_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.06 10.88 7.2 11.365 ;
    END
  END bottom_left_grid_pin_49_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.35 0.8 59.65 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 53.91 0.8 54.21 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 62.07 0.8 62.37 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.63 0.8 56.93 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.63 0.8 22.93 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 47.11 0.8 47.41 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.03 0.8 43.33 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.47 0.8 48.77 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 66.83 0.8 67.13 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 72.27 0.8 72.57 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 41.67 0.8 41.97 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 57.99 0.8 58.29 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 60.71 0.8 61.01 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 87.91 0.8 88.21 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 45.75 0.8 46.05 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.55 0.8 69.85 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 63.43 0.8 63.73 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 70.91 0.8 71.21 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 85.19 0.8 85.49 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 68.19 0.8 68.49 ;
    END
  END chanx_left_in[19]
  PIN left_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 6.75 10.88 7.05 11.68 ;
    END
  END left_bottom_grid_pin_34_[0]
  PIN left_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 8.59 10.88 8.89 11.68 ;
    END
  END left_bottom_grid_pin_35_[0]
  PIN left_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.9 10.88 9.04 11.365 ;
    END
  END left_bottom_grid_pin_36_[0]
  PIN left_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.98 10.88 8.12 11.365 ;
    END
  END left_bottom_grid_pin_37_[0]
  PIN left_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.66 10.88 11.8 11.365 ;
    END
  END left_bottom_grid_pin_38_[0]
  PIN left_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.58 10.88 12.72 11.365 ;
    END
  END left_bottom_grid_pin_39_[0]
  PIN left_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.56 10.88 18.7 11.365 ;
    END
  END left_bottom_grid_pin_40_[0]
  PIN left_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.14 10.88 6.28 11.365 ;
    END
  END left_bottom_grid_pin_41_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.52 108.315 30.66 108.8 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.52 108.315 76.66 108.8 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.86 108.315 44 108.8 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.6 108.315 75.74 108.8 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.44 108.315 77.58 108.8 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.96 108.315 60.1 108.8 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.62 108.315 46.76 108.8 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.9 108.315 55.04 108.8 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.36 108.315 78.5 108.8 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.86 108.315 67 108.8 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.82 108.315 55.96 108.8 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.54 108.315 47.68 108.8 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 108.315 61.48 108.8 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 108.315 38.48 108.8 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.28 108.315 79.42 108.8 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.76 108.315 50.9 108.8 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.84 108.315 49.98 108.8 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.36 108.315 32.5 108.8 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.92 108.315 72.06 108.8 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.28 108.315 33.42 108.8 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71 108.315 71.14 108.8 ;
    END
  END chany_top_out[19]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 0 38.48 0.485 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.68 0 74.82 0.485 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.44 0 31.58 0.485 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 0 62.4 0.485 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.48 0 65.62 0.485 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.38 0 49.52 0.485 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.32 0 67.46 0.485 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.24 0 68.38 0.485 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.04 0 59.18 0.485 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.3 0 50.44 0.485 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.12 0 35.26 0.485 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 0 61.48 0.485 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.96 0 60.1 0.485 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.5 0 82.64 0.485 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 0 56.42 0.485 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.12 0 58.26 0.485 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48 0 48.14 0.485 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.84 0 72.98 0.485 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.74 0 33.88 0.485 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.92 0 72.06 0.485 ;
    END
  END chany_bottom_out[19]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 23.99 0.8 24.29 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 64.79 0.8 65.09 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 34.87 0.8 35.17 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 55.27 0.8 55.57 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 15.83 0.8 16.13 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.39 0.8 44.69 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.51 0.8 33.81 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.35 0.8 25.65 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 30.79 0.8 31.09 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 49.83 0.8 50.13 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.23 0.8 36.53 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.55 0.8 52.85 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 17.19 0.8 17.49 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 86.55 0.8 86.85 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.59 0.8 37.89 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 28.07 0.8 28.37 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 14.47 0.8 14.77 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 51.19 0.8 51.49 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 32.15 0.8 32.45 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 26.71 0.8 27.01 ;
    END
  END chanx_left_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.43 0.8 29.73 ;
    END
  END ccff_tail[0]
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 37.42 108.315 37.56 108.8 ;
    END
  END prog_clk_0_N_in
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 25.76 2.48 26.24 2.96 ;
        RECT 91.52 2.48 92 2.96 ;
        RECT 25.76 7.92 26.24 8.4 ;
        RECT 91.52 7.92 92 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 91.52 13.36 92 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 91.52 18.8 92 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 91.52 24.24 92 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 91.52 29.68 92 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 91.52 35.12 92 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 91.52 40.56 92 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 91.52 46 92 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 91.52 51.44 92 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 91.52 56.88 92 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 91.52 62.32 92 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 91.52 67.76 92 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 91.52 73.2 92 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 91.52 78.64 92 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 91.52 84.08 92 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 91.52 89.52 92 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 91.52 94.96 92 95.44 ;
        RECT 25.76 100.4 26.24 100.88 ;
        RECT 91.52 100.4 92 100.88 ;
        RECT 25.76 105.84 26.24 106.32 ;
        RECT 91.52 105.84 92 106.32 ;
      LAYER met5 ;
        RECT 0 22.2 3.2 25.4 ;
        RECT 88.8 22.2 92 25.4 ;
        RECT 0 63 3.2 66.2 ;
        RECT 88.8 63 92 66.2 ;
      LAYER met4 ;
        RECT 36.5 0 37.1 0.6 ;
        RECT 65.94 0 66.54 0.6 ;
        RECT 36.5 108.2 37.1 108.8 ;
        RECT 65.94 108.2 66.54 108.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 25.76 0 45.4 0.24 ;
        RECT 46.6 0 92 0.24 ;
        RECT 25.76 5.2 26.24 5.68 ;
        RECT 91.52 5.2 92 5.68 ;
        RECT 0 10.64 45.4 11.12 ;
        RECT 91.52 10.64 92 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 91.52 16.08 92 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 91.52 21.52 92 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 91.52 26.96 92 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 91.52 32.4 92 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 91.52 37.84 92 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 91.52 43.28 92 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 91.52 48.72 92 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 91.52 54.16 92 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 91.52 59.6 92 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 91.52 65.04 92 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 91.52 70.48 92 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 91.52 75.92 92 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 91.52 81.36 92 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 91.52 86.8 92 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 91.52 92.24 92 92.72 ;
        RECT 0 97.68 45.4 98.16 ;
        RECT 91.52 97.68 92 98.16 ;
        RECT 25.76 103.12 26.24 103.6 ;
        RECT 91.52 103.12 92 103.6 ;
        RECT 25.76 108.56 45.4 108.8 ;
        RECT 46.6 108.56 92 108.8 ;
      LAYER met5 ;
        RECT 0 42.6 3.2 45.8 ;
        RECT 88.8 42.6 92 45.8 ;
        RECT 0 83.4 3.2 86.6 ;
        RECT 88.8 83.4 92 86.6 ;
      LAYER met4 ;
        RECT 51.22 0 51.82 0.6 ;
        RECT 80.66 0 81.26 0.6 ;
        RECT 10.74 10.88 11.34 11.48 ;
        RECT 10.74 97.32 11.34 97.92 ;
        RECT 51.22 108.2 51.82 108.8 ;
        RECT 80.66 108.2 81.26 108.8 ;
    END
  END VSS
  OBS
    LAYER met2 ;
      RECT 80.82 108.615 81.1 108.985 ;
      RECT 51.38 108.615 51.66 108.985 ;
      POLYGON 75.28 108.7 75.28 70.14 75.14 70.14 75.14 108.56 75.1 108.56 75.1 108.7 ;
      RECT 63.58 107.79 63.84 108.11 ;
      RECT 10.9 97.735 11.18 98.105 ;
      RECT 9.76 96.91 10.02 97.23 ;
      POLYGON 20.08 23.02 20.08 11.405 20.15 11.405 20.15 11.035 19.87 11.035 19.87 11.405 19.94 11.405 19.94 23.02 ;
      RECT 10.9 10.695 11.18 11.065 ;
      RECT 64.96 0.69 65.22 1.01 ;
      RECT 80.82 -0.185 81.1 0.185 ;
      RECT 51.38 -0.185 51.66 0.185 ;
      POLYGON 91.72 108.52 91.72 0.28 82.92 0.28 82.92 0.765 82.22 0.765 82.22 0.28 82 0.28 82 0.765 81.3 0.765 81.3 0.28 80.62 0.28 80.62 0.765 79.92 0.765 79.92 0.28 79.7 0.28 79.7 0.765 79 0.765 79 0.28 78.78 0.28 78.78 0.765 78.08 0.765 78.08 0.28 77.86 0.28 77.86 0.765 77.16 0.765 77.16 0.28 76.94 0.28 76.94 0.765 76.24 0.765 76.24 0.28 76.02 0.28 76.02 0.765 75.32 0.765 75.32 0.28 75.1 0.28 75.1 0.765 74.4 0.765 74.4 0.28 74.18 0.28 74.18 0.765 73.48 0.765 73.48 0.28 73.26 0.28 73.26 0.765 72.56 0.765 72.56 0.28 72.34 0.28 72.34 0.765 71.64 0.765 71.64 0.28 71.42 0.28 71.42 0.765 70.72 0.765 70.72 0.28 70.5 0.28 70.5 0.765 69.8 0.765 69.8 0.28 69.58 0.28 69.58 0.765 68.88 0.765 68.88 0.28 68.66 0.28 68.66 0.765 67.96 0.765 67.96 0.28 67.74 0.28 67.74 0.765 67.04 0.765 67.04 0.28 66.82 0.28 66.82 0.765 66.12 0.765 66.12 0.28 65.9 0.28 65.9 0.765 65.2 0.765 65.2 0.28 64.98 0.28 64.98 0.765 64.28 0.765 64.28 0.28 64.06 0.28 64.06 0.765 63.36 0.765 63.36 0.28 62.68 0.28 62.68 0.765 61.98 0.765 61.98 0.28 61.76 0.28 61.76 0.765 61.06 0.765 61.06 0.28 60.38 0.28 60.38 0.765 59.68 0.765 59.68 0.28 59.46 0.28 59.46 0.765 58.76 0.765 58.76 0.28 58.54 0.28 58.54 0.765 57.84 0.765 57.84 0.28 57.62 0.28 57.62 0.765 56.92 0.765 56.92 0.28 56.7 0.28 56.7 0.765 56 0.765 56 0.28 55.78 0.28 55.78 0.765 55.08 0.765 55.08 0.28 54.86 0.28 54.86 0.765 54.16 0.765 54.16 0.28 53.48 0.28 53.48 0.765 52.78 0.765 52.78 0.28 52.56 0.28 52.56 0.765 51.86 0.765 51.86 0.28 50.72 0.28 50.72 0.765 50.02 0.765 50.02 0.28 49.8 0.28 49.8 0.765 49.1 0.765 49.1 0.28 48.42 0.28 48.42 0.765 47.72 0.765 47.72 0.28 47.5 0.28 47.5 0.765 46.8 0.765 46.8 0.28 38.76 0.28 38.76 0.765 38.06 0.765 38.06 0.28 35.54 0.28 35.54 0.765 34.84 0.765 34.84 0.28 34.16 0.28 34.16 0.765 33.46 0.765 33.46 0.28 32.78 0.28 32.78 0.765 32.08 0.765 32.08 0.28 31.86 0.28 31.86 0.765 31.16 0.765 31.16 0.28 26.04 0.28 26.04 11.16 18.98 11.16 18.98 11.645 18.28 11.645 18.28 11.16 15.76 11.16 15.76 11.645 15.06 11.645 15.06 11.16 14.84 11.16 14.84 11.645 14.14 11.645 14.14 11.16 13.92 11.16 13.92 11.645 13.22 11.645 13.22 11.16 13 11.16 13 11.645 12.3 11.645 12.3 11.16 12.08 11.16 12.08 11.645 11.38 11.645 11.38 11.16 10.7 11.16 10.7 11.645 10 11.645 10 11.16 9.32 11.16 9.32 11.645 8.62 11.645 8.62 11.16 8.4 11.16 8.4 11.645 7.7 11.645 7.7 11.16 7.48 11.16 7.48 11.645 6.78 11.645 6.78 11.16 6.56 11.16 6.56 11.645 5.86 11.645 5.86 11.16 5.64 11.16 5.64 11.645 4.94 11.645 4.94 11.16 4.72 11.16 4.72 11.645 4.02 11.645 4.02 11.16 3.34 11.16 3.34 11.645 2.64 11.645 2.64 11.16 0.28 11.16 0.28 97.64 4.02 97.64 4.02 97.155 4.72 97.155 4.72 97.64 6.78 97.64 6.78 97.155 7.48 97.155 7.48 97.64 8.16 97.64 8.16 97.155 8.86 97.155 8.86 97.64 9.08 97.64 9.08 97.155 9.78 97.155 9.78 97.64 10 97.64 10 97.155 10.7 97.155 10.7 97.64 11.38 97.64 11.38 97.155 12.08 97.155 12.08 97.64 12.3 97.64 12.3 97.155 13 97.155 13 97.64 13.22 97.64 13.22 97.155 13.92 97.155 13.92 97.64 26.04 97.64 26.04 108.52 30.24 108.52 30.24 108.035 30.94 108.035 30.94 108.52 31.16 108.52 31.16 108.035 31.86 108.035 31.86 108.52 32.08 108.52 32.08 108.035 32.78 108.035 32.78 108.52 33 108.52 33 108.035 33.7 108.035 33.7 108.52 37.14 108.52 37.14 108.035 37.84 108.035 37.84 108.52 38.06 108.52 38.06 108.035 38.76 108.035 38.76 108.52 43.58 108.52 43.58 108.035 44.28 108.035 44.28 108.52 44.5 108.52 44.5 108.035 45.2 108.035 45.2 108.52 45.42 108.52 45.42 108.035 46.12 108.035 46.12 108.52 46.34 108.52 46.34 108.035 47.04 108.035 47.04 108.52 47.26 108.52 47.26 108.035 47.96 108.035 47.96 108.52 48.18 108.52 48.18 108.035 48.88 108.035 48.88 108.52 49.56 108.52 49.56 108.035 50.26 108.035 50.26 108.52 50.48 108.52 50.48 108.035 51.18 108.035 51.18 108.52 51.86 108.52 51.86 108.035 52.56 108.035 52.56 108.52 52.78 108.52 52.78 108.035 53.48 108.035 53.48 108.52 53.7 108.52 53.7 108.035 54.4 108.035 54.4 108.52 54.62 108.52 54.62 108.035 55.32 108.035 55.32 108.52 55.54 108.52 55.54 108.035 56.24 108.035 56.24 108.52 56.46 108.52 56.46 108.035 57.16 108.035 57.16 108.52 57.84 108.52 57.84 108.035 58.54 108.035 58.54 108.52 58.76 108.52 58.76 108.035 59.46 108.035 59.46 108.52 59.68 108.52 59.68 108.035 60.38 108.035 60.38 108.52 61.06 108.52 61.06 108.035 61.76 108.035 61.76 108.52 61.98 108.52 61.98 108.035 62.68 108.035 62.68 108.52 62.9 108.52 62.9 108.035 63.6 108.035 63.6 108.52 63.82 108.52 63.82 108.035 64.52 108.035 64.52 108.52 64.74 108.52 64.74 108.035 65.44 108.035 65.44 108.52 65.66 108.52 65.66 108.035 66.36 108.035 66.36 108.52 66.58 108.52 66.58 108.035 67.28 108.035 67.28 108.52 67.5 108.52 67.5 108.035 68.2 108.035 68.2 108.52 68.88 108.52 68.88 108.035 69.58 108.035 69.58 108.52 69.8 108.52 69.8 108.035 70.5 108.035 70.5 108.52 70.72 108.52 70.72 108.035 71.42 108.035 71.42 108.52 71.64 108.52 71.64 108.035 72.34 108.035 72.34 108.52 72.56 108.52 72.56 108.035 73.26 108.035 73.26 108.52 73.48 108.52 73.48 108.035 74.18 108.035 74.18 108.52 74.4 108.52 74.4 108.035 75.1 108.035 75.1 108.52 75.32 108.52 75.32 108.035 76.02 108.035 76.02 108.52 76.24 108.52 76.24 108.035 76.94 108.035 76.94 108.52 77.16 108.52 77.16 108.035 77.86 108.035 77.86 108.52 78.08 108.52 78.08 108.035 78.78 108.035 78.78 108.52 79 108.52 79 108.035 79.7 108.035 79.7 108.52 ;
    LAYER met3 ;
      POLYGON 81.125 108.965 81.125 108.96 81.34 108.96 81.34 108.64 81.125 108.64 81.125 108.635 80.795 108.635 80.795 108.64 80.58 108.64 80.58 108.96 80.795 108.96 80.795 108.965 ;
      POLYGON 51.685 108.965 51.685 108.96 51.9 108.96 51.9 108.64 51.685 108.64 51.685 108.635 51.355 108.635 51.355 108.64 51.14 108.64 51.14 108.96 51.355 108.96 51.355 108.965 ;
      POLYGON 55.135 108.625 55.135 108.295 54.805 108.295 54.805 108.3 54.395 108.3 54.395 108.62 54.805 108.62 54.805 108.625 ;
      POLYGON 11.205 98.085 11.205 98.08 11.42 98.08 11.42 97.76 11.205 97.76 11.205 97.755 10.875 97.755 10.875 97.76 10.66 97.76 10.66 98.08 10.875 98.08 10.875 98.085 ;
      POLYGON 8.89 13.41 8.89 11.38 8.93 11.38 8.93 11.06 8.55 11.06 8.55 11.38 8.59 11.38 8.59 13.41 ;
      POLYGON 20.175 11.385 20.175 11.055 19.845 11.055 19.845 11.07 15.575 11.07 15.575 11.055 15.245 11.055 15.245 11.385 15.575 11.385 15.575 11.37 19.845 11.37 19.845 11.385 ;
      POLYGON 11.205 11.045 11.205 11.04 11.42 11.04 11.42 10.72 11.205 10.72 11.205 10.715 10.875 10.715 10.875 10.72 10.66 10.72 10.66 11.04 10.875 11.04 10.875 11.045 ;
      POLYGON 81.125 0.165 81.125 0.16 81.34 0.16 81.34 -0.16 81.125 -0.16 81.125 -0.165 80.795 -0.165 80.795 -0.16 80.58 -0.16 80.58 0.16 80.795 0.16 80.795 0.165 ;
      POLYGON 51.685 0.165 51.685 0.16 51.9 0.16 51.9 -0.16 51.685 -0.16 51.685 -0.165 51.355 -0.165 51.355 -0.16 51.14 -0.16 51.14 0.16 51.355 0.16 51.355 0.165 ;
      POLYGON 91.6 108.4 91.6 0.4 26.16 0.4 26.16 11.28 0.4 11.28 0.4 14.07 1.2 14.07 1.2 15.17 0.4 15.17 0.4 15.43 1.2 15.43 1.2 16.53 0.4 16.53 0.4 16.79 1.2 16.79 1.2 17.89 0.4 17.89 0.4 22.23 1.2 22.23 1.2 23.33 0.4 23.33 0.4 23.59 1.2 23.59 1.2 24.69 0.4 24.69 0.4 24.95 1.2 24.95 1.2 26.05 0.4 26.05 0.4 26.31 1.2 26.31 1.2 27.41 0.4 27.41 0.4 27.67 1.2 27.67 1.2 28.77 0.4 28.77 0.4 29.03 1.2 29.03 1.2 30.13 0.4 30.13 0.4 30.39 1.2 30.39 1.2 31.49 0.4 31.49 0.4 31.75 1.2 31.75 1.2 32.85 0.4 32.85 0.4 33.11 1.2 33.11 1.2 34.21 0.4 34.21 0.4 34.47 1.2 34.47 1.2 35.57 0.4 35.57 0.4 35.83 1.2 35.83 1.2 36.93 0.4 36.93 0.4 37.19 1.2 37.19 1.2 38.29 0.4 38.29 0.4 41.27 1.2 41.27 1.2 42.37 0.4 42.37 0.4 42.63 1.2 42.63 1.2 43.73 0.4 43.73 0.4 43.99 1.2 43.99 1.2 45.09 0.4 45.09 0.4 45.35 1.2 45.35 1.2 46.45 0.4 46.45 0.4 46.71 1.2 46.71 1.2 47.81 0.4 47.81 0.4 48.07 1.2 48.07 1.2 49.17 0.4 49.17 0.4 49.43 1.2 49.43 1.2 50.53 0.4 50.53 0.4 50.79 1.2 50.79 1.2 51.89 0.4 51.89 0.4 52.15 1.2 52.15 1.2 53.25 0.4 53.25 0.4 53.51 1.2 53.51 1.2 54.61 0.4 54.61 0.4 54.87 1.2 54.87 1.2 55.97 0.4 55.97 0.4 56.23 1.2 56.23 1.2 57.33 0.4 57.33 0.4 57.59 1.2 57.59 1.2 58.69 0.4 58.69 0.4 58.95 1.2 58.95 1.2 60.05 0.4 60.05 0.4 60.31 1.2 60.31 1.2 61.41 0.4 61.41 0.4 61.67 1.2 61.67 1.2 62.77 0.4 62.77 0.4 63.03 1.2 63.03 1.2 64.13 0.4 64.13 0.4 64.39 1.2 64.39 1.2 65.49 0.4 65.49 0.4 66.43 1.2 66.43 1.2 67.53 0.4 67.53 0.4 67.79 1.2 67.79 1.2 68.89 0.4 68.89 0.4 69.15 1.2 69.15 1.2 70.25 0.4 70.25 0.4 70.51 1.2 70.51 1.2 71.61 0.4 71.61 0.4 71.87 1.2 71.87 1.2 72.97 0.4 72.97 0.4 84.79 1.2 84.79 1.2 85.89 0.4 85.89 0.4 86.15 1.2 86.15 1.2 87.25 0.4 87.25 0.4 87.51 1.2 87.51 1.2 88.61 0.4 88.61 0.4 97.52 26.16 97.52 26.16 108.4 ;
    LAYER met4 ;
      POLYGON 54.905 108.625 54.905 108.295 54.89 108.295 54.89 77.03 54.59 77.03 54.59 108.295 54.575 108.295 54.575 108.625 ;
      POLYGON 91.6 108.4 91.6 0.4 81.66 0.4 81.66 1 80.26 1 80.26 0.4 66.94 0.4 66.94 1 65.54 1 65.54 0.4 52.22 0.4 52.22 1 50.82 1 50.82 0.4 37.5 0.4 37.5 1 36.1 1 36.1 0.4 26.16 0.4 26.16 11.28 11.74 11.28 11.74 11.88 10.34 11.88 10.34 11.28 9.29 11.28 9.29 12.08 8.19 12.08 8.19 11.28 7.45 11.28 7.45 12.08 6.35 12.08 6.35 11.28 0.4 11.28 0.4 97.52 10.34 97.52 10.34 96.92 11.74 96.92 11.74 97.52 26.16 97.52 26.16 108.4 36.1 108.4 36.1 107.8 37.5 107.8 37.5 108.4 50.82 108.4 50.82 107.8 52.22 107.8 52.22 108.4 65.54 108.4 65.54 107.8 66.94 107.8 66.94 108.4 80.26 108.4 80.26 107.8 81.66 107.8 81.66 108.4 ;
    LAYER met5 ;
      POLYGON 90.4 107.2 90.4 88.2 87.2 88.2 87.2 81.8 90.4 81.8 90.4 67.8 87.2 67.8 87.2 61.4 90.4 61.4 90.4 47.4 87.2 47.4 87.2 41 90.4 41 90.4 27 87.2 27 87.2 20.6 90.4 20.6 90.4 1.6 27.36 1.6 27.36 12.48 1.6 12.48 1.6 20.6 4.8 20.6 4.8 27 1.6 27 1.6 41 4.8 41 4.8 47.4 1.6 47.4 1.6 61.4 4.8 61.4 4.8 67.8 1.6 67.8 1.6 81.8 4.8 81.8 4.8 88.2 1.6 88.2 1.6 96.32 27.36 96.32 27.36 107.2 ;
    LAYER met1 ;
      RECT 45.68 108.56 46.32 109.04 ;
      POLYGON 36.64 98.84 36.64 98.5 40.105 98.5 40.105 98.545 40.395 98.545 40.395 98.315 40.105 98.315 40.105 98.36 36.5 98.36 36.5 98.84 ;
      POLYGON 34.34 98.84 34.34 98.545 34.415 98.545 34.415 98.315 34.125 98.315 34.125 98.545 34.2 98.545 34.2 98.84 ;
      RECT 42.39 98.3 42.71 98.56 ;
      RECT 35.49 98.3 35.81 98.56 ;
      RECT 31.81 98.3 32.13 98.56 ;
      POLYGON 34.43 97.54 34.43 97.48 59.18 97.48 59.18 97.34 34.43 97.34 34.43 97.28 34.11 97.28 34.11 97.54 ;
      POLYGON 28.45 97.54 28.45 97.28 28.13 97.28 28.13 97.34 12.81 97.34 12.81 97.28 12.49 97.28 12.49 97.54 12.81 97.54 12.81 97.48 28.13 97.48 28.13 97.54 ;
      POLYGON 9.5 11.8 9.5 11.32 1.31 11.32 1.31 11.26 0.99 11.26 0.99 11.52 1.31 11.52 1.31 11.46 9.36 11.46 9.36 11.8 ;
      POLYGON 34.43 11.52 34.43 11.46 44.705 11.46 44.705 11.505 44.995 11.505 44.995 11.275 44.705 11.275 44.705 11.32 34.43 11.32 34.43 11.26 34.11 11.26 34.11 11.52 ;
      POLYGON 28.45 11.52 28.45 11.26 28.13 11.26 28.13 11.275 27.775 11.275 27.775 11.505 28.13 11.505 28.13 11.52 ;
      POLYGON 76.2 1.26 76.2 0.58 77.35 0.58 77.35 0.64 77.67 0.64 77.67 0.38 77.35 0.38 77.35 0.44 76.06 0.44 76.06 1.26 ;
      RECT 45.68 -0.24 46.32 0.24 ;
      POLYGON 46.32 108.52 46.32 108.28 91.72 108.28 91.72 106.6 91.24 106.6 91.24 105.56 91.72 105.56 91.72 103.88 91.24 103.88 91.24 102.84 91.72 102.84 91.72 101.16 91.24 101.16 91.24 100.12 91.72 100.12 91.72 98.44 91.24 98.44 91.24 97.4 91.72 97.4 91.72 95.72 91.24 95.72 91.24 94.68 91.72 94.68 91.72 93 91.24 93 91.24 91.96 91.72 91.96 91.72 90.28 91.24 90.28 91.24 89.24 91.72 89.24 91.72 87.56 91.24 87.56 91.24 86.52 91.72 86.52 91.72 84.84 91.24 84.84 91.24 83.8 91.72 83.8 91.72 82.12 91.24 82.12 91.24 81.08 91.72 81.08 91.72 79.4 91.24 79.4 91.24 78.36 91.72 78.36 91.72 76.68 91.24 76.68 91.24 75.64 91.72 75.64 91.72 73.96 91.24 73.96 91.24 72.92 91.72 72.92 91.72 71.24 91.24 71.24 91.24 70.2 91.72 70.2 91.72 68.52 91.24 68.52 91.24 67.48 91.72 67.48 91.72 65.8 91.24 65.8 91.24 64.76 91.72 64.76 91.72 63.08 91.24 63.08 91.24 62.04 91.72 62.04 91.72 60.36 91.24 60.36 91.24 59.32 91.72 59.32 91.72 57.64 91.24 57.64 91.24 56.6 91.72 56.6 91.72 54.92 91.24 54.92 91.24 53.88 91.72 53.88 91.72 52.2 91.24 52.2 91.24 51.16 91.72 51.16 91.72 49.48 91.24 49.48 91.24 48.44 91.72 48.44 91.72 46.76 91.24 46.76 91.24 45.72 91.72 45.72 91.72 44.04 91.24 44.04 91.24 43 91.72 43 91.72 41.32 91.24 41.32 91.24 40.28 91.72 40.28 91.72 38.6 91.24 38.6 91.24 37.56 91.72 37.56 91.72 35.88 91.24 35.88 91.24 34.84 91.72 34.84 91.72 33.16 91.24 33.16 91.24 32.12 91.72 32.12 91.72 30.44 91.24 30.44 91.24 29.4 91.72 29.4 91.72 27.72 91.24 27.72 91.24 26.68 91.72 26.68 91.72 25 91.24 25 91.24 23.96 91.72 23.96 91.72 22.28 91.24 22.28 91.24 21.24 91.72 21.24 91.72 19.56 91.24 19.56 91.24 18.52 91.72 18.52 91.72 16.84 91.24 16.84 91.24 15.8 91.72 15.8 91.72 14.12 91.24 14.12 91.24 13.08 91.72 13.08 91.72 11.4 91.24 11.4 91.24 10.36 91.72 10.36 91.72 8.68 91.24 8.68 91.24 7.64 91.72 7.64 91.72 5.96 91.24 5.96 91.24 4.92 91.72 4.92 91.72 3.24 91.24 3.24 91.24 2.2 91.72 2.2 91.72 0.52 46.32 0.52 46.32 0.28 45.68 0.28 45.68 0.52 26.04 0.52 26.04 2.2 26.52 2.2 26.52 3.24 26.04 3.24 26.04 4.92 26.52 4.92 26.52 5.96 26.04 5.96 26.04 7.64 26.52 7.64 26.52 8.68 26.04 8.68 26.04 10.36 45.68 10.36 45.68 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 45.68 97.4 45.68 98.44 26.04 98.44 26.04 100.12 26.52 100.12 26.52 101.16 26.04 101.16 26.04 102.84 26.52 102.84 26.52 103.88 26.04 103.88 26.04 105.56 26.52 105.56 26.52 106.6 26.04 106.6 26.04 108.28 45.68 108.28 45.68 108.52 ;
    LAYER li1 ;
      POLYGON 92 108.885 92 108.715 89.615 108.715 89.615 107.99 89.325 107.99 89.325 108.715 82.255 108.715 82.255 107.99 81.965 107.99 81.965 108.715 74.005 108.715 74.005 108.235 73.675 108.235 73.675 108.715 73.165 108.715 73.165 108.235 72.835 108.235 72.835 108.715 72.325 108.715 72.325 108.235 71.995 108.235 71.995 108.715 71.485 108.715 71.485 108.235 71.155 108.235 71.155 108.715 70.645 108.715 70.645 108.235 70.315 108.235 70.315 108.715 69.805 108.715 69.805 107.915 69.475 107.915 69.475 108.715 67.535 108.715 67.535 107.99 67.245 107.99 67.245 108.715 65.725 108.715 65.725 108.235 65.395 108.235 65.395 108.715 64.885 108.715 64.885 108.235 64.555 108.235 64.555 108.715 64.045 108.715 64.045 108.235 63.715 108.235 63.715 108.715 63.205 108.715 63.205 108.235 62.875 108.235 62.875 108.715 62.365 108.715 62.365 108.235 62.035 108.235 62.035 108.715 61.525 108.715 61.525 107.915 61.195 107.915 61.195 108.715 57.485 108.715 57.485 107.915 57.155 107.915 57.155 108.715 56.645 108.715 56.645 108.235 56.315 108.235 56.315 108.715 55.805 108.715 55.805 108.235 55.475 108.235 55.475 108.715 54.965 108.715 54.965 108.235 54.635 108.235 54.635 108.715 54.125 108.715 54.125 108.235 53.795 108.235 53.795 108.715 53.285 108.715 53.285 108.235 52.955 108.235 52.955 108.715 52.355 108.715 52.355 107.99 52.065 107.99 52.065 108.715 48.205 108.715 48.205 107.915 47.875 107.915 47.875 108.715 47.365 108.715 47.365 108.235 47.035 108.235 47.035 108.715 46.525 108.715 46.525 108.235 46.195 108.235 46.195 108.715 45.605 108.715 45.605 108.235 45.435 108.235 45.435 108.715 44.765 108.715 44.765 108.235 44.595 108.235 44.595 108.715 37.635 108.715 37.635 107.99 37.345 107.99 37.345 108.715 36.625 108.715 36.625 108.105 36.455 108.105 36.455 108.715 35.695 108.715 35.695 108.185 35.485 108.185 35.485 108.715 33.67 108.715 33.67 108.215 33.3 108.215 33.3 108.715 31.605 108.715 31.605 108.255 31.355 108.255 31.355 108.715 30.745 108.715 30.745 108.335 30.415 108.335 30.415 108.715 29.815 108.715 29.815 107.99 29.525 107.99 29.525 108.715 25.76 108.715 25.76 108.885 ;
      RECT 91.54 105.995 92 106.165 ;
      RECT 25.76 105.995 29.44 106.165 ;
      RECT 91.54 103.275 92 103.445 ;
      RECT 25.76 103.275 29.44 103.445 ;
      RECT 91.54 100.555 92 100.725 ;
      RECT 25.76 100.555 29.44 100.725 ;
      RECT 91.54 97.835 92 98.005 ;
      POLYGON 29.44 98.005 29.44 97.835 26.155 97.835 26.155 97.455 25.825 97.455 25.825 97.835 22.455 97.835 22.455 97.11 22.165 97.11 22.165 97.835 20.645 97.835 20.645 97.435 20.315 97.435 20.315 97.835 18.355 97.835 18.355 97.3 17.845 97.3 17.845 97.835 14.545 97.835 14.545 97.225 14.375 97.225 14.375 97.835 13.615 97.835 13.615 97.305 13.405 97.305 13.405 97.835 11.59 97.835 11.59 97.335 11.22 97.335 11.22 97.835 9.525 97.835 9.525 97.375 9.275 97.375 9.275 97.835 8.665 97.835 8.665 97.455 8.335 97.455 8.335 97.835 7.735 97.835 7.735 97.11 7.445 97.11 7.445 97.835 0 97.835 0 98.005 ;
      RECT 91.54 95.115 92 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 91.54 92.395 92 92.565 ;
      RECT 0 92.395 1.84 92.565 ;
      RECT 91.54 89.675 92 89.845 ;
      RECT 0 89.675 1.84 89.845 ;
      RECT 91.54 86.955 92 87.125 ;
      RECT 0 86.955 1.84 87.125 ;
      RECT 91.54 84.235 92 84.405 ;
      RECT 0 84.235 1.84 84.405 ;
      RECT 91.54 81.515 92 81.685 ;
      RECT 0 81.515 1.84 81.685 ;
      RECT 91.54 78.795 92 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 91.54 76.075 92 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 91.54 73.355 92 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 91.54 70.635 92 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 91.54 67.915 92 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 91.08 65.195 92 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 91.08 62.475 92 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 91.54 59.755 92 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 91.54 57.035 92 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 91.54 54.315 92 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 91.54 51.595 92 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 91.54 48.875 92 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 91.54 46.155 92 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 90.16 43.435 92 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 90.16 40.715 92 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 91.54 37.995 92 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 91.54 35.275 92 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 91.54 32.555 92 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 91.54 29.835 92 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 91.54 27.115 92 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 91.54 24.395 92 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 91.54 21.675 92 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 91.54 18.955 92 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 91.54 16.235 92 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 91.54 13.515 92 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      POLYGON 5.66 11.785 5.66 10.965 7.445 10.965 7.445 11.69 7.735 11.69 7.735 10.965 8.835 10.965 8.835 11.765 9.165 11.765 9.165 10.965 9.675 10.965 9.675 11.445 10.005 11.445 10.005 10.965 10.515 10.965 10.515 11.445 10.845 11.445 10.845 10.965 11.435 10.965 11.435 11.445 11.605 11.445 11.605 10.965 12.275 10.965 12.275 11.445 12.445 11.445 12.445 10.965 15.235 10.965 15.235 11.345 15.565 11.345 15.565 10.965 16.175 10.965 16.175 11.425 16.425 11.425 16.425 10.965 18.12 10.965 18.12 11.465 18.49 11.465 18.49 10.965 20.305 10.965 20.305 11.495 20.515 11.495 20.515 10.965 21.275 10.965 21.275 11.575 21.445 11.575 21.445 10.965 22.165 10.965 22.165 11.69 22.455 11.69 22.455 10.965 25.735 10.965 25.735 11.445 25.905 11.445 25.905 10.965 26.575 10.965 26.575 11.445 26.745 11.445 26.745 10.965 27.335 10.965 27.335 11.445 27.665 11.445 27.665 10.965 28.175 10.965 28.175 11.445 28.505 11.445 28.505 10.965 29.015 10.965 29.015 11.765 29.345 11.765 29.345 10.965 29.44 10.965 29.44 10.795 0 10.795 0 10.965 5.43 10.965 5.43 11.785 ;
      RECT 88.32 10.795 92 10.965 ;
      RECT 88.32 8.075 92 8.245 ;
      RECT 25.76 8.075 29.44 8.245 ;
      RECT 91.54 5.355 92 5.525 ;
      RECT 25.76 5.355 29.44 5.525 ;
      RECT 91.54 2.635 92 2.805 ;
      RECT 25.76 2.635 29.44 2.805 ;
      POLYGON 87.845 0.885 87.845 0.085 89.325 0.085 89.325 0.81 89.615 0.81 89.615 0.085 92 0.085 92 -0.085 25.76 -0.085 25.76 0.085 29.525 0.085 29.525 0.81 29.815 0.81 29.815 0.085 30.335 0.085 30.335 0.565 30.505 0.565 30.505 0.085 31.175 0.085 31.175 0.565 31.345 0.565 31.345 0.085 31.935 0.085 31.935 0.565 32.265 0.565 32.265 0.085 32.775 0.085 32.775 0.565 33.105 0.565 33.105 0.085 33.615 0.085 33.615 0.885 33.945 0.885 33.945 0.085 37.345 0.085 37.345 0.81 37.635 0.81 37.635 0.085 41.415 0.085 41.415 0.885 41.745 0.885 41.745 0.085 42.255 0.085 42.255 0.565 42.585 0.565 42.585 0.085 43.095 0.085 43.095 0.565 43.425 0.565 43.425 0.085 43.935 0.085 43.935 0.565 44.265 0.565 44.265 0.085 44.775 0.085 44.775 0.565 45.105 0.565 45.105 0.085 45.615 0.085 45.615 0.565 45.945 0.565 45.945 0.085 46.935 0.085 46.935 0.885 47.265 0.885 47.265 0.085 47.775 0.085 47.775 0.565 48.105 0.565 48.105 0.085 48.615 0.085 48.615 0.565 48.945 0.565 48.945 0.085 49.455 0.085 49.455 0.565 49.785 0.565 49.785 0.085 50.295 0.085 50.295 0.565 50.625 0.565 50.625 0.085 51.135 0.085 51.135 0.565 51.465 0.565 51.465 0.085 52.065 0.085 52.065 0.81 52.355 0.81 52.355 0.085 53.875 0.085 53.875 0.565 54.205 0.565 54.205 0.085 54.715 0.085 54.715 0.565 55.045 0.565 55.045 0.085 55.555 0.085 55.555 0.565 55.885 0.565 55.885 0.085 56.395 0.085 56.395 0.565 56.725 0.565 56.725 0.085 57.235 0.085 57.235 0.565 57.565 0.565 57.565 0.085 58.075 0.085 58.075 0.885 58.405 0.885 58.405 0.085 60.735 0.085 60.735 0.885 61.065 0.885 61.065 0.085 61.575 0.085 61.575 0.565 61.905 0.565 61.905 0.085 62.415 0.085 62.415 0.565 62.745 0.565 62.745 0.085 63.255 0.085 63.255 0.565 63.585 0.565 63.585 0.085 64.095 0.085 64.095 0.565 64.425 0.565 64.425 0.085 64.935 0.085 64.935 0.565 65.265 0.565 65.265 0.085 67.245 0.085 67.245 0.81 67.535 0.81 67.535 0.085 71.315 0.085 71.315 0.885 71.645 0.885 71.645 0.085 72.155 0.085 72.155 0.565 72.485 0.565 72.485 0.085 72.995 0.085 72.995 0.565 73.325 0.565 73.325 0.085 73.835 0.085 73.835 0.565 74.165 0.565 74.165 0.085 74.675 0.085 74.675 0.565 75.005 0.565 75.005 0.085 75.515 0.085 75.515 0.565 75.845 0.565 75.845 0.085 76.875 0.085 76.875 0.565 77.205 0.565 77.205 0.085 77.715 0.085 77.715 0.565 78.045 0.565 78.045 0.085 78.555 0.085 78.555 0.565 78.885 0.565 78.885 0.085 79.395 0.085 79.395 0.565 79.725 0.565 79.725 0.085 80.235 0.085 80.235 0.565 80.565 0.565 80.565 0.085 81.075 0.085 81.075 0.885 81.405 0.885 81.405 0.085 81.965 0.085 81.965 0.81 82.255 0.81 82.255 0.085 83.315 0.085 83.315 0.565 83.645 0.565 83.645 0.085 84.155 0.085 84.155 0.565 84.485 0.565 84.485 0.085 84.995 0.085 84.995 0.565 85.325 0.565 85.325 0.085 85.835 0.085 85.835 0.565 86.165 0.565 86.165 0.085 86.675 0.085 86.675 0.565 87.005 0.565 87.005 0.085 87.515 0.085 87.515 0.885 ;
      POLYGON 91.83 108.63 91.83 0.17 25.93 0.17 25.93 11.05 0.17 11.05 0.17 97.75 25.93 97.75 25.93 108.63 ;
    LAYER mcon ;
      RECT 42.465 98.345 42.635 98.515 ;
      RECT 40.165 98.345 40.335 98.515 ;
      RECT 35.565 98.345 35.735 98.515 ;
      RECT 34.185 98.345 34.355 98.515 ;
      RECT 31.885 98.345 32.055 98.515 ;
      RECT 44.765 11.305 44.935 11.475 ;
      RECT 27.835 11.305 28.005 11.475 ;
    LAYER via ;
      RECT 80.885 108.725 81.035 108.875 ;
      RECT 51.445 108.725 51.595 108.875 ;
      RECT 42.475 98.355 42.625 98.505 ;
      RECT 35.575 98.355 35.725 98.505 ;
      RECT 31.895 98.355 32.045 98.505 ;
      RECT 10.965 97.845 11.115 97.995 ;
      RECT 34.195 97.335 34.345 97.485 ;
      RECT 28.215 97.335 28.365 97.485 ;
      RECT 12.575 97.335 12.725 97.485 ;
      RECT 34.195 11.315 34.345 11.465 ;
      RECT 28.215 11.315 28.365 11.465 ;
      RECT 1.075 11.315 1.225 11.465 ;
      RECT 10.965 10.805 11.115 10.955 ;
      RECT 77.435 0.435 77.585 0.585 ;
      RECT 80.885 -0.075 81.035 0.075 ;
      RECT 51.445 -0.075 51.595 0.075 ;
    LAYER via2 ;
      RECT 80.86 108.7 81.06 108.9 ;
      RECT 51.42 108.7 51.62 108.9 ;
      RECT 54.87 108.36 55.07 108.56 ;
      RECT 10.94 97.82 11.14 98.02 ;
      RECT 1.05 62.12 1.25 62.32 ;
      RECT 1.05 15.88 1.25 16.08 ;
      RECT 19.91 11.12 20.11 11.32 ;
      RECT 15.31 11.12 15.51 11.32 ;
      RECT 10.94 10.78 11.14 10.98 ;
      RECT 80.86 -0.1 81.06 0.1 ;
      RECT 51.42 -0.1 51.62 0.1 ;
    LAYER via3 ;
      RECT 80.86 108.7 81.06 108.9 ;
      RECT 51.42 108.7 51.62 108.9 ;
      RECT 54.64 108.36 54.84 108.56 ;
      RECT 10.94 97.82 11.14 98.02 ;
      RECT 8.64 11.12 8.84 11.32 ;
      RECT 10.94 10.78 11.14 10.98 ;
      RECT 80.86 -0.1 81.06 0.1 ;
      RECT 51.42 -0.1 51.62 0.1 ;
    LAYER OVERLAP ;
      POLYGON 25.76 0 25.76 10.88 0 10.88 0 97.92 25.76 97.92 25.76 108.8 92 108.8 92 0 ;
  END
END sb_2__1_

END LIBRARY
