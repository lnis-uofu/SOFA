VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_2__0_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 84.64 BY 81.6 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 2.23 63.92 2.37 65.28 ;
    END
  END prog_clk[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.51 80.24 56.65 81.6 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.05 80.24 33.19 81.6 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.89 80.24 57.19 81.6 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.13 80.24 32.27 81.6 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.93 80.24 23.07 81.6 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.15 80.24 49.29 81.6 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.87 80.24 64.01 81.6 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 80.24 57.57 81.6 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.03 80.24 62.17 81.6 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.85 80.24 46.15 81.6 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.61 80.24 48.91 81.6 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 80.24 48.37 81.6 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 80.24 52.97 81.6 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.79 80.24 64.93 81.6 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.11 80.24 61.25 81.6 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.27 80.24 59.41 81.6 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 80.24 50.21 81.6 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.95 80.24 63.09 81.6 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.35 80.24 58.49 81.6 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.19 80.24 60.33 81.6 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.69 80.24 24.99 81.6 ;
    END
  END top_left_grid_pin_42_[0]
  PIN top_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.97 63.92 11.11 65.28 ;
    END
  END top_left_grid_pin_43_[0]
  PIN top_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.85 80.24 23.15 81.6 ;
    END
  END top_left_grid_pin_44_[0]
  PIN top_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.27 63.92 13.41 65.28 ;
    END
  END top_left_grid_pin_45_[0]
  PIN top_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.63 80.24 20.77 81.6 ;
    END
  END top_left_grid_pin_46_[0]
  PIN top_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.67 63.92 8.81 65.28 ;
    END
  END top_left_grid_pin_47_[0]
  PIN top_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.55 80.24 21.69 81.6 ;
    END
  END top_left_grid_pin_48_[0]
  PIN top_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.53 80.24 26.83 81.6 ;
    END
  END top_left_grid_pin_49_[0]
  PIN top_right_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.85 80.24 23.99 81.6 ;
    END
  END top_right_grid_pin_1_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 3.93 1.38 4.23 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 55.61 1.38 55.91 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 38.61 1.38 38.91 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 12.09 1.38 12.39 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.89 1.38 53.19 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 16.17 1.38 16.47 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 20.25 1.38 20.55 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 6.65 1.38 6.95 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 9.37 1.38 9.67 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 21.61 1.38 21.91 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 41.33 1.38 41.63 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.53 63.92 4.67 65.28 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 5.29 1.38 5.59 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 4.45 63.92 4.75 65.28 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.61 63.92 3.75 65.28 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.17 1.38 50.47 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 47.45 1.38 47.75 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 51.53 1.38 51.83 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.97 1.38 23.27 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 24.33 1.38 24.63 ;
    END
  END chanx_left_in[19]
  PIN left_bottom_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.05 1.38 44.35 ;
    END
  END left_bottom_grid_pin_1_[0]
  PIN left_bottom_grid_pin_3_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.81 1.38 49.11 ;
    END
  END left_bottom_grid_pin_3_[0]
  PIN left_bottom_grid_pin_5_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.57 1.38 36.87 ;
    END
  END left_bottom_grid_pin_5_[0]
  PIN left_bottom_grid_pin_7_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 30.45 1.38 30.75 ;
    END
  END left_bottom_grid_pin_7_[0]
  PIN left_bottom_grid_pin_9_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.69 1.38 42.99 ;
    END
  END left_bottom_grid_pin_9_[0]
  PIN left_bottom_grid_pin_11_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 46.09 1.38 46.39 ;
    END
  END left_bottom_grid_pin_11_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.03 80.24 39.17 81.6 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.87 80.24 41.01 81.6 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.97 80.24 34.11 81.6 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 80.24 46.53 81.6 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 80.24 52.05 81.6 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.17 80.24 43.31 81.6 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.69 80.24 25.83 81.6 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.35 80.24 35.49 81.6 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 80.24 47.45 81.6 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.65 80.24 37.79 81.6 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 80.24 51.13 81.6 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.73 80.24 36.87 81.6 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.75 80.24 53.89 81.6 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.37 80.24 29.51 81.6 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.95 80.24 40.09 81.6 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.61 80.24 26.75 81.6 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 80.24 45.61 81.6 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.77 80.24 24.91 81.6 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.45 80.24 28.59 81.6 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.25 80.24 42.39 81.6 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.53 80.24 27.67 81.6 ;
    END
  END chany_top_out[19]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 58.33 1.38 58.63 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.97 1.38 57.27 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.97 1.38 40.27 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.45 63.92 5.59 65.28 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 54.25 1.38 54.55 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 61.05 1.38 61.35 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.15 0 3.29 1.36 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.69 1.38 59.99 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.81 1.38 32.11 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.23 0 2.37 1.36 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 18.89 1.38 19.19 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 34.53 1.38 34.83 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.09 1.38 29.39 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 8.01 1.38 8.31 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.69 1.38 25.99 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 17.53 1.38 17.83 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.17 1.38 33.47 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 14.81 1.38 15.11 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 27.05 1.38 27.35 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 10.73 1.38 11.03 ;
    END
  END chanx_left_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 13.45 1.38 13.75 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 84.16 2.48 84.64 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 84.16 7.92 84.64 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 84.16 13.36 84.64 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 84.16 18.8 84.64 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 84.16 24.24 84.64 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 84.16 29.68 84.64 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 84.16 35.12 84.64 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 84.16 40.56 84.64 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 84.16 46 84.64 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 84.16 51.44 84.64 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 84.16 56.88 84.64 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 84.16 62.32 84.64 62.8 ;
        RECT 18.4 67.76 18.88 68.24 ;
        RECT 84.16 67.76 84.64 68.24 ;
        RECT 18.4 73.2 18.88 73.68 ;
        RECT 84.16 73.2 84.64 73.68 ;
        RECT 18.4 78.64 18.88 79.12 ;
        RECT 84.16 78.64 84.64 79.12 ;
      LAYER met4 ;
        RECT 29.14 0 29.74 0.6 ;
        RECT 58.58 0 59.18 0.6 ;
        RECT 29.14 81 29.74 81.6 ;
        RECT 58.58 81 59.18 81.6 ;
      LAYER met5 ;
        RECT 0 10.64 3.2 13.84 ;
        RECT 81.44 10.64 84.64 13.84 ;
        RECT 0 51.44 3.2 54.64 ;
        RECT 81.44 51.44 84.64 54.64 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 0 84.64 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 84.16 5.2 84.64 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 84.16 10.64 84.64 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 84.16 16.08 84.64 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 84.16 21.52 84.64 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 84.16 26.96 84.64 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 84.16 32.4 84.64 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 84.16 37.84 84.64 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 84.16 43.28 84.64 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 84.16 48.72 84.64 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 84.16 54.16 84.64 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 84.16 59.6 84.64 60.08 ;
        RECT 0 65.04 84.64 65.52 ;
        RECT 18.4 70.48 18.88 70.96 ;
        RECT 84.16 70.48 84.64 70.96 ;
        RECT 18.4 75.92 18.88 76.4 ;
        RECT 84.16 75.92 84.64 76.4 ;
        RECT 18.4 81.36 84.64 81.6 ;
      LAYER met4 ;
        RECT 43.86 0 44.46 0.6 ;
        RECT 73.3 0 73.9 0.6 ;
        RECT 43.86 81 44.46 81.6 ;
        RECT 73.3 81 73.9 81.6 ;
      LAYER met5 ;
        RECT 0 31.04 3.2 34.24 ;
        RECT 81.44 31.04 84.64 34.24 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 18.4 81.515 84.64 81.685 ;
      RECT 80.96 78.795 84.64 78.965 ;
      RECT 18.4 78.795 22.08 78.965 ;
      RECT 80.96 76.075 84.64 76.245 ;
      RECT 18.4 76.075 22.08 76.245 ;
      RECT 80.96 73.355 84.64 73.525 ;
      RECT 18.4 73.355 22.08 73.525 ;
      RECT 80.96 70.635 84.64 70.805 ;
      RECT 18.4 70.635 20.24 70.805 ;
      RECT 80.96 67.915 84.64 68.085 ;
      RECT 18.4 67.915 22.08 68.085 ;
      RECT 80.96 65.195 84.64 65.365 ;
      RECT 0 65.195 22.08 65.365 ;
      RECT 84.18 62.475 84.64 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 84.18 59.755 84.64 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 80.96 57.035 84.64 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 80.96 54.315 84.64 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 80.96 51.595 84.64 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 80.96 48.875 84.64 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 80.96 46.155 84.64 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 83.72 43.435 84.64 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 84.18 40.715 84.64 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 84.18 37.995 84.64 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 84.18 35.275 84.64 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 83.72 32.555 84.64 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 83.72 29.835 84.64 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 83.72 27.115 84.64 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 80.96 24.395 84.64 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 80.96 21.675 84.64 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 82.8 18.955 84.64 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 80.96 16.235 84.64 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 80.96 13.515 84.64 13.685 ;
      RECT 0 13.515 1.84 13.685 ;
      RECT 83.72 10.795 84.64 10.965 ;
      RECT 0 10.795 1.84 10.965 ;
      RECT 83.72 8.075 84.64 8.245 ;
      RECT 0 8.075 1.84 8.245 ;
      RECT 83.72 5.355 84.64 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 84.18 2.635 84.64 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 84.64 0.085 ;
    LAYER met2 ;
      RECT 73.46 81.415 73.74 81.785 ;
      RECT 44.02 81.415 44.3 81.785 ;
      RECT 34.37 79.74 34.63 80.06 ;
      RECT 73.46 -0.185 73.74 0.185 ;
      RECT 44.02 -0.185 44.3 0.185 ;
      POLYGON 84.36 81.32 84.36 0.28 3.57 0.28 3.57 1.64 2.87 1.64 2.87 0.28 2.65 0.28 2.65 1.64 1.95 1.64 1.95 0.28 0.28 0.28 0.28 65 1.95 65 1.95 63.64 2.65 63.64 2.65 65 3.33 65 3.33 63.64 4.03 63.64 4.03 65 4.25 65 4.25 63.64 4.95 63.64 4.95 65 5.17 65 5.17 63.64 5.87 63.64 5.87 65 8.39 65 8.39 63.64 9.09 63.64 9.09 65 10.69 65 10.69 63.64 11.39 63.64 11.39 65 12.99 65 12.99 63.64 13.69 63.64 13.69 65 18.68 65 18.68 81.32 20.35 81.32 20.35 79.96 21.05 79.96 21.05 81.32 21.27 81.32 21.27 79.96 21.97 79.96 21.97 81.32 22.65 81.32 22.65 79.96 23.35 79.96 23.35 81.32 23.57 81.32 23.57 79.96 24.27 79.96 24.27 81.32 24.49 81.32 24.49 79.96 25.19 79.96 25.19 81.32 25.41 81.32 25.41 79.96 26.11 79.96 26.11 81.32 26.33 81.32 26.33 79.96 27.03 79.96 27.03 81.32 27.25 81.32 27.25 79.96 27.95 79.96 27.95 81.32 28.17 81.32 28.17 79.96 28.87 79.96 28.87 81.32 29.09 81.32 29.09 79.96 29.79 79.96 29.79 81.32 31.85 81.32 31.85 79.96 32.55 79.96 32.55 81.32 32.77 81.32 32.77 79.96 33.47 79.96 33.47 81.32 33.69 81.32 33.69 79.96 34.39 79.96 34.39 81.32 35.07 81.32 35.07 79.96 35.77 79.96 35.77 81.32 36.45 81.32 36.45 79.96 37.15 79.96 37.15 81.32 37.37 81.32 37.37 79.96 38.07 79.96 38.07 81.32 38.75 81.32 38.75 79.96 39.45 79.96 39.45 81.32 39.67 81.32 39.67 79.96 40.37 79.96 40.37 81.32 40.59 81.32 40.59 79.96 41.29 79.96 41.29 81.32 41.97 81.32 41.97 79.96 42.67 79.96 42.67 81.32 42.89 81.32 42.89 79.96 43.59 79.96 43.59 81.32 45.19 81.32 45.19 79.96 45.89 79.96 45.89 81.32 46.11 81.32 46.11 79.96 46.81 79.96 46.81 81.32 47.03 81.32 47.03 79.96 47.73 79.96 47.73 81.32 47.95 81.32 47.95 79.96 48.65 79.96 48.65 81.32 48.87 81.32 48.87 79.96 49.57 79.96 49.57 81.32 49.79 81.32 49.79 79.96 50.49 79.96 50.49 81.32 50.71 81.32 50.71 79.96 51.41 79.96 51.41 81.32 51.63 81.32 51.63 79.96 52.33 79.96 52.33 81.32 52.55 81.32 52.55 79.96 53.25 79.96 53.25 81.32 53.47 81.32 53.47 79.96 54.17 79.96 54.17 81.32 56.23 81.32 56.23 79.96 56.93 79.96 56.93 81.32 57.15 81.32 57.15 79.96 57.85 79.96 57.85 81.32 58.07 81.32 58.07 79.96 58.77 79.96 58.77 81.32 58.99 81.32 58.99 79.96 59.69 79.96 59.69 81.32 59.91 81.32 59.91 79.96 60.61 79.96 60.61 81.32 60.83 81.32 60.83 79.96 61.53 79.96 61.53 81.32 61.75 81.32 61.75 79.96 62.45 79.96 62.45 81.32 62.67 81.32 62.67 79.96 63.37 79.96 63.37 81.32 63.59 81.32 63.59 79.96 64.29 79.96 64.29 81.32 64.51 81.32 64.51 79.96 65.21 79.96 65.21 81.32 ;
    LAYER met4 ;
      POLYGON 84.24 81.2 84.24 0.4 74.3 0.4 74.3 1 72.9 1 72.9 0.4 59.58 0.4 59.58 1 58.18 1 58.18 0.4 44.86 0.4 44.86 1 43.46 1 43.46 0.4 30.14 0.4 30.14 1 28.74 1 28.74 0.4 0.4 0.4 0.4 64.88 4.05 64.88 4.05 63.52 5.15 63.52 5.15 64.88 18.8 64.88 18.8 81.2 22.45 81.2 22.45 79.84 23.55 79.84 23.55 81.2 24.29 81.2 24.29 79.84 25.39 79.84 25.39 81.2 26.13 81.2 26.13 79.84 27.23 79.84 27.23 81.2 28.74 81.2 28.74 80.6 30.14 80.6 30.14 81.2 43.46 81.2 43.46 80.6 44.86 80.6 44.86 81.2 45.45 81.2 45.45 79.84 46.55 79.84 46.55 81.2 48.21 81.2 48.21 79.84 49.31 79.84 49.31 81.2 56.49 81.2 56.49 79.84 57.59 79.84 57.59 81.2 58.18 81.2 58.18 80.6 59.58 80.6 59.58 81.2 72.9 81.2 72.9 80.6 74.3 80.6 74.3 81.2 ;
    LAYER met3 ;
      POLYGON 73.765 81.765 73.765 81.76 73.98 81.76 73.98 81.44 73.765 81.44 73.765 81.435 73.435 81.435 73.435 81.44 73.22 81.44 73.22 81.76 73.435 81.76 73.435 81.765 ;
      POLYGON 44.325 81.765 44.325 81.76 44.54 81.76 44.54 81.44 44.325 81.44 44.325 81.435 43.995 81.435 43.995 81.44 43.78 81.44 43.78 81.76 43.995 81.76 43.995 81.765 ;
      POLYGON 73.765 0.165 73.765 0.16 73.98 0.16 73.98 -0.16 73.765 -0.16 73.765 -0.165 73.435 -0.165 73.435 -0.16 73.22 -0.16 73.22 0.16 73.435 0.16 73.435 0.165 ;
      POLYGON 44.325 0.165 44.325 0.16 44.54 0.16 44.54 -0.16 44.325 -0.16 44.325 -0.165 43.995 -0.165 43.995 -0.16 43.78 -0.16 43.78 0.16 43.995 0.16 43.995 0.165 ;
      POLYGON 84.24 81.2 84.24 0.4 0.4 0.4 0.4 3.53 1.78 3.53 1.78 4.63 0.4 4.63 0.4 4.89 1.78 4.89 1.78 5.99 0.4 5.99 0.4 6.25 1.78 6.25 1.78 7.35 0.4 7.35 0.4 7.61 1.78 7.61 1.78 8.71 0.4 8.71 0.4 8.97 1.78 8.97 1.78 10.07 0.4 10.07 0.4 10.33 1.78 10.33 1.78 11.43 0.4 11.43 0.4 11.69 1.78 11.69 1.78 12.79 0.4 12.79 0.4 13.05 1.78 13.05 1.78 14.15 0.4 14.15 0.4 14.41 1.78 14.41 1.78 15.51 0.4 15.51 0.4 15.77 1.78 15.77 1.78 16.87 0.4 16.87 0.4 17.13 1.78 17.13 1.78 18.23 0.4 18.23 0.4 18.49 1.78 18.49 1.78 19.59 0.4 19.59 0.4 19.85 1.78 19.85 1.78 20.95 0.4 20.95 0.4 21.21 1.78 21.21 1.78 22.31 0.4 22.31 0.4 22.57 1.78 22.57 1.78 23.67 0.4 23.67 0.4 23.93 1.78 23.93 1.78 25.03 0.4 25.03 0.4 25.29 1.78 25.29 1.78 26.39 0.4 26.39 0.4 26.65 1.78 26.65 1.78 27.75 0.4 27.75 0.4 28.69 1.78 28.69 1.78 29.79 0.4 29.79 0.4 30.05 1.78 30.05 1.78 31.15 0.4 31.15 0.4 31.41 1.78 31.41 1.78 32.51 0.4 32.51 0.4 32.77 1.78 32.77 1.78 33.87 0.4 33.87 0.4 34.13 1.78 34.13 1.78 35.23 0.4 35.23 0.4 36.17 1.78 36.17 1.78 37.27 0.4 37.27 0.4 38.21 1.78 38.21 1.78 39.31 0.4 39.31 0.4 39.57 1.78 39.57 1.78 40.67 0.4 40.67 0.4 40.93 1.78 40.93 1.78 42.03 0.4 42.03 0.4 42.29 1.78 42.29 1.78 43.39 0.4 43.39 0.4 43.65 1.78 43.65 1.78 44.75 0.4 44.75 0.4 45.69 1.78 45.69 1.78 46.79 0.4 46.79 0.4 47.05 1.78 47.05 1.78 48.15 0.4 48.15 0.4 48.41 1.78 48.41 1.78 49.51 0.4 49.51 0.4 49.77 1.78 49.77 1.78 50.87 0.4 50.87 0.4 51.13 1.78 51.13 1.78 52.23 0.4 52.23 0.4 52.49 1.78 52.49 1.78 53.59 0.4 53.59 0.4 53.85 1.78 53.85 1.78 54.95 0.4 54.95 0.4 55.21 1.78 55.21 1.78 56.31 0.4 56.31 0.4 56.57 1.78 56.57 1.78 57.67 0.4 57.67 0.4 57.93 1.78 57.93 1.78 59.03 0.4 59.03 0.4 59.29 1.78 59.29 1.78 60.39 0.4 60.39 0.4 60.65 1.78 60.65 1.78 61.75 0.4 61.75 0.4 64.88 18.8 64.88 18.8 81.2 ;
    LAYER met5 ;
      POLYGON 83.04 80 83.04 56.24 79.84 56.24 79.84 49.84 83.04 49.84 83.04 35.84 79.84 35.84 79.84 29.44 83.04 29.44 83.04 15.44 79.84 15.44 79.84 9.04 83.04 9.04 83.04 1.6 1.6 1.6 1.6 9.04 4.8 9.04 4.8 15.44 1.6 15.44 1.6 29.44 4.8 29.44 4.8 35.84 1.6 35.84 1.6 49.84 4.8 49.84 4.8 56.24 1.6 56.24 1.6 63.68 20 63.68 20 80 ;
    LAYER met1 ;
      POLYGON 84.36 81.08 84.36 79.4 83.88 79.4 83.88 78.36 84.36 78.36 84.36 76.68 83.88 76.68 83.88 75.64 84.36 75.64 84.36 73.96 83.88 73.96 83.88 72.92 84.36 72.92 84.36 71.24 83.88 71.24 83.88 70.2 84.36 70.2 84.36 68.52 83.88 68.52 83.88 67.48 84.36 67.48 84.36 65.8 18.68 65.8 18.68 67.48 19.16 67.48 19.16 68.52 18.68 68.52 18.68 70.2 19.16 70.2 19.16 71.24 18.68 71.24 18.68 72.92 19.16 72.92 19.16 73.96 18.68 73.96 18.68 75.64 19.16 75.64 19.16 76.68 18.68 76.68 18.68 78.36 19.16 78.36 19.16 79.4 18.68 79.4 18.68 81.08 ;
      POLYGON 84.36 64.76 84.36 63.08 83.88 63.08 83.88 62.04 84.36 62.04 84.36 60.36 83.88 60.36 83.88 59.32 84.36 59.32 84.36 57.64 83.88 57.64 83.88 56.6 84.36 56.6 84.36 54.92 83.88 54.92 83.88 53.88 84.36 53.88 84.36 52.2 83.88 52.2 83.88 51.16 84.36 51.16 84.36 49.48 83.88 49.48 83.88 48.44 84.36 48.44 84.36 46.76 83.88 46.76 83.88 45.72 84.36 45.72 84.36 44.04 83.88 44.04 83.88 43 84.36 43 84.36 41.32 83.88 41.32 83.88 40.28 84.36 40.28 84.36 38.6 83.88 38.6 83.88 37.56 84.36 37.56 84.36 35.88 83.88 35.88 83.88 34.84 84.36 34.84 84.36 33.16 83.88 33.16 83.88 32.12 84.36 32.12 84.36 30.44 83.88 30.44 83.88 29.4 84.36 29.4 84.36 27.72 83.88 27.72 83.88 26.68 84.36 26.68 84.36 25 83.88 25 83.88 23.96 84.36 23.96 84.36 22.28 83.88 22.28 83.88 21.24 84.36 21.24 84.36 19.56 83.88 19.56 83.88 18.52 84.36 18.52 84.36 16.84 83.88 16.84 83.88 15.8 84.36 15.8 84.36 14.12 83.88 14.12 83.88 13.08 84.36 13.08 84.36 11.4 83.88 11.4 83.88 10.36 84.36 10.36 84.36 8.68 83.88 8.68 83.88 7.64 84.36 7.64 84.36 5.96 83.88 5.96 83.88 4.92 84.36 4.92 84.36 3.24 83.88 3.24 83.88 2.2 84.36 2.2 84.36 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 ;
    LAYER li1 ;
      POLYGON 84.47 81.43 84.47 0.17 0.17 0.17 0.17 65.11 18.57 65.11 18.57 81.43 ;
    LAYER mcon ;
      RECT 84.325 81.515 84.495 81.685 ;
      RECT 83.865 81.515 84.035 81.685 ;
      RECT 83.405 81.515 83.575 81.685 ;
      RECT 82.945 81.515 83.115 81.685 ;
      RECT 82.485 81.515 82.655 81.685 ;
      RECT 82.025 81.515 82.195 81.685 ;
      RECT 81.565 81.515 81.735 81.685 ;
      RECT 81.105 81.515 81.275 81.685 ;
      RECT 80.645 81.515 80.815 81.685 ;
      RECT 80.185 81.515 80.355 81.685 ;
      RECT 79.725 81.515 79.895 81.685 ;
      RECT 79.265 81.515 79.435 81.685 ;
      RECT 78.805 81.515 78.975 81.685 ;
      RECT 78.345 81.515 78.515 81.685 ;
      RECT 77.885 81.515 78.055 81.685 ;
      RECT 77.425 81.515 77.595 81.685 ;
      RECT 76.965 81.515 77.135 81.685 ;
      RECT 76.505 81.515 76.675 81.685 ;
      RECT 76.045 81.515 76.215 81.685 ;
      RECT 75.585 81.515 75.755 81.685 ;
      RECT 75.125 81.515 75.295 81.685 ;
      RECT 74.665 81.515 74.835 81.685 ;
      RECT 74.205 81.515 74.375 81.685 ;
      RECT 73.745 81.515 73.915 81.685 ;
      RECT 73.285 81.515 73.455 81.685 ;
      RECT 72.825 81.515 72.995 81.685 ;
      RECT 72.365 81.515 72.535 81.685 ;
      RECT 71.905 81.515 72.075 81.685 ;
      RECT 71.445 81.515 71.615 81.685 ;
      RECT 70.985 81.515 71.155 81.685 ;
      RECT 70.525 81.515 70.695 81.685 ;
      RECT 70.065 81.515 70.235 81.685 ;
      RECT 69.605 81.515 69.775 81.685 ;
      RECT 69.145 81.515 69.315 81.685 ;
      RECT 68.685 81.515 68.855 81.685 ;
      RECT 68.225 81.515 68.395 81.685 ;
      RECT 67.765 81.515 67.935 81.685 ;
      RECT 67.305 81.515 67.475 81.685 ;
      RECT 66.845 81.515 67.015 81.685 ;
      RECT 66.385 81.515 66.555 81.685 ;
      RECT 65.925 81.515 66.095 81.685 ;
      RECT 65.465 81.515 65.635 81.685 ;
      RECT 65.005 81.515 65.175 81.685 ;
      RECT 64.545 81.515 64.715 81.685 ;
      RECT 64.085 81.515 64.255 81.685 ;
      RECT 63.625 81.515 63.795 81.685 ;
      RECT 63.165 81.515 63.335 81.685 ;
      RECT 62.705 81.515 62.875 81.685 ;
      RECT 62.245 81.515 62.415 81.685 ;
      RECT 61.785 81.515 61.955 81.685 ;
      RECT 61.325 81.515 61.495 81.685 ;
      RECT 60.865 81.515 61.035 81.685 ;
      RECT 60.405 81.515 60.575 81.685 ;
      RECT 59.945 81.515 60.115 81.685 ;
      RECT 59.485 81.515 59.655 81.685 ;
      RECT 59.025 81.515 59.195 81.685 ;
      RECT 58.565 81.515 58.735 81.685 ;
      RECT 58.105 81.515 58.275 81.685 ;
      RECT 57.645 81.515 57.815 81.685 ;
      RECT 57.185 81.515 57.355 81.685 ;
      RECT 56.725 81.515 56.895 81.685 ;
      RECT 56.265 81.515 56.435 81.685 ;
      RECT 55.805 81.515 55.975 81.685 ;
      RECT 55.345 81.515 55.515 81.685 ;
      RECT 54.885 81.515 55.055 81.685 ;
      RECT 54.425 81.515 54.595 81.685 ;
      RECT 53.965 81.515 54.135 81.685 ;
      RECT 53.505 81.515 53.675 81.685 ;
      RECT 53.045 81.515 53.215 81.685 ;
      RECT 52.585 81.515 52.755 81.685 ;
      RECT 52.125 81.515 52.295 81.685 ;
      RECT 51.665 81.515 51.835 81.685 ;
      RECT 51.205 81.515 51.375 81.685 ;
      RECT 50.745 81.515 50.915 81.685 ;
      RECT 50.285 81.515 50.455 81.685 ;
      RECT 49.825 81.515 49.995 81.685 ;
      RECT 49.365 81.515 49.535 81.685 ;
      RECT 48.905 81.515 49.075 81.685 ;
      RECT 48.445 81.515 48.615 81.685 ;
      RECT 47.985 81.515 48.155 81.685 ;
      RECT 47.525 81.515 47.695 81.685 ;
      RECT 47.065 81.515 47.235 81.685 ;
      RECT 46.605 81.515 46.775 81.685 ;
      RECT 46.145 81.515 46.315 81.685 ;
      RECT 45.685 81.515 45.855 81.685 ;
      RECT 45.225 81.515 45.395 81.685 ;
      RECT 44.765 81.515 44.935 81.685 ;
      RECT 44.305 81.515 44.475 81.685 ;
      RECT 43.845 81.515 44.015 81.685 ;
      RECT 43.385 81.515 43.555 81.685 ;
      RECT 42.925 81.515 43.095 81.685 ;
      RECT 42.465 81.515 42.635 81.685 ;
      RECT 42.005 81.515 42.175 81.685 ;
      RECT 41.545 81.515 41.715 81.685 ;
      RECT 41.085 81.515 41.255 81.685 ;
      RECT 40.625 81.515 40.795 81.685 ;
      RECT 40.165 81.515 40.335 81.685 ;
      RECT 39.705 81.515 39.875 81.685 ;
      RECT 39.245 81.515 39.415 81.685 ;
      RECT 38.785 81.515 38.955 81.685 ;
      RECT 38.325 81.515 38.495 81.685 ;
      RECT 37.865 81.515 38.035 81.685 ;
      RECT 37.405 81.515 37.575 81.685 ;
      RECT 36.945 81.515 37.115 81.685 ;
      RECT 36.485 81.515 36.655 81.685 ;
      RECT 36.025 81.515 36.195 81.685 ;
      RECT 35.565 81.515 35.735 81.685 ;
      RECT 35.105 81.515 35.275 81.685 ;
      RECT 34.645 81.515 34.815 81.685 ;
      RECT 34.185 81.515 34.355 81.685 ;
      RECT 33.725 81.515 33.895 81.685 ;
      RECT 33.265 81.515 33.435 81.685 ;
      RECT 32.805 81.515 32.975 81.685 ;
      RECT 32.345 81.515 32.515 81.685 ;
      RECT 31.885 81.515 32.055 81.685 ;
      RECT 31.425 81.515 31.595 81.685 ;
      RECT 30.965 81.515 31.135 81.685 ;
      RECT 30.505 81.515 30.675 81.685 ;
      RECT 30.045 81.515 30.215 81.685 ;
      RECT 29.585 81.515 29.755 81.685 ;
      RECT 29.125 81.515 29.295 81.685 ;
      RECT 28.665 81.515 28.835 81.685 ;
      RECT 28.205 81.515 28.375 81.685 ;
      RECT 27.745 81.515 27.915 81.685 ;
      RECT 27.285 81.515 27.455 81.685 ;
      RECT 26.825 81.515 26.995 81.685 ;
      RECT 26.365 81.515 26.535 81.685 ;
      RECT 25.905 81.515 26.075 81.685 ;
      RECT 25.445 81.515 25.615 81.685 ;
      RECT 24.985 81.515 25.155 81.685 ;
      RECT 24.525 81.515 24.695 81.685 ;
      RECT 24.065 81.515 24.235 81.685 ;
      RECT 23.605 81.515 23.775 81.685 ;
      RECT 23.145 81.515 23.315 81.685 ;
      RECT 22.685 81.515 22.855 81.685 ;
      RECT 22.225 81.515 22.395 81.685 ;
      RECT 21.765 81.515 21.935 81.685 ;
      RECT 21.305 81.515 21.475 81.685 ;
      RECT 20.845 81.515 21.015 81.685 ;
      RECT 20.385 81.515 20.555 81.685 ;
      RECT 19.925 81.515 20.095 81.685 ;
      RECT 19.465 81.515 19.635 81.685 ;
      RECT 19.005 81.515 19.175 81.685 ;
      RECT 18.545 81.515 18.715 81.685 ;
      RECT 84.325 78.795 84.495 78.965 ;
      RECT 83.865 78.795 84.035 78.965 ;
      RECT 19.005 78.795 19.175 78.965 ;
      RECT 18.545 78.795 18.715 78.965 ;
      RECT 84.325 76.075 84.495 76.245 ;
      RECT 83.865 76.075 84.035 76.245 ;
      RECT 19.005 76.075 19.175 76.245 ;
      RECT 18.545 76.075 18.715 76.245 ;
      RECT 84.325 73.355 84.495 73.525 ;
      RECT 83.865 73.355 84.035 73.525 ;
      RECT 19.005 73.355 19.175 73.525 ;
      RECT 18.545 73.355 18.715 73.525 ;
      RECT 84.325 70.635 84.495 70.805 ;
      RECT 83.865 70.635 84.035 70.805 ;
      RECT 19.005 70.635 19.175 70.805 ;
      RECT 18.545 70.635 18.715 70.805 ;
      RECT 84.325 67.915 84.495 68.085 ;
      RECT 83.865 67.915 84.035 68.085 ;
      RECT 19.005 67.915 19.175 68.085 ;
      RECT 18.545 67.915 18.715 68.085 ;
      RECT 84.325 65.195 84.495 65.365 ;
      RECT 83.865 65.195 84.035 65.365 ;
      RECT 83.405 65.195 83.575 65.365 ;
      RECT 82.945 65.195 83.115 65.365 ;
      RECT 82.485 65.195 82.655 65.365 ;
      RECT 82.025 65.195 82.195 65.365 ;
      RECT 81.565 65.195 81.735 65.365 ;
      RECT 81.105 65.195 81.275 65.365 ;
      RECT 80.645 65.195 80.815 65.365 ;
      RECT 80.185 65.195 80.355 65.365 ;
      RECT 79.725 65.195 79.895 65.365 ;
      RECT 79.265 65.195 79.435 65.365 ;
      RECT 78.805 65.195 78.975 65.365 ;
      RECT 78.345 65.195 78.515 65.365 ;
      RECT 77.885 65.195 78.055 65.365 ;
      RECT 77.425 65.195 77.595 65.365 ;
      RECT 76.965 65.195 77.135 65.365 ;
      RECT 76.505 65.195 76.675 65.365 ;
      RECT 76.045 65.195 76.215 65.365 ;
      RECT 75.585 65.195 75.755 65.365 ;
      RECT 75.125 65.195 75.295 65.365 ;
      RECT 74.665 65.195 74.835 65.365 ;
      RECT 74.205 65.195 74.375 65.365 ;
      RECT 73.745 65.195 73.915 65.365 ;
      RECT 73.285 65.195 73.455 65.365 ;
      RECT 72.825 65.195 72.995 65.365 ;
      RECT 72.365 65.195 72.535 65.365 ;
      RECT 71.905 65.195 72.075 65.365 ;
      RECT 71.445 65.195 71.615 65.365 ;
      RECT 70.985 65.195 71.155 65.365 ;
      RECT 70.525 65.195 70.695 65.365 ;
      RECT 70.065 65.195 70.235 65.365 ;
      RECT 69.605 65.195 69.775 65.365 ;
      RECT 69.145 65.195 69.315 65.365 ;
      RECT 68.685 65.195 68.855 65.365 ;
      RECT 68.225 65.195 68.395 65.365 ;
      RECT 67.765 65.195 67.935 65.365 ;
      RECT 67.305 65.195 67.475 65.365 ;
      RECT 66.845 65.195 67.015 65.365 ;
      RECT 66.385 65.195 66.555 65.365 ;
      RECT 65.925 65.195 66.095 65.365 ;
      RECT 65.465 65.195 65.635 65.365 ;
      RECT 65.005 65.195 65.175 65.365 ;
      RECT 64.545 65.195 64.715 65.365 ;
      RECT 64.085 65.195 64.255 65.365 ;
      RECT 63.625 65.195 63.795 65.365 ;
      RECT 63.165 65.195 63.335 65.365 ;
      RECT 62.705 65.195 62.875 65.365 ;
      RECT 62.245 65.195 62.415 65.365 ;
      RECT 61.785 65.195 61.955 65.365 ;
      RECT 61.325 65.195 61.495 65.365 ;
      RECT 60.865 65.195 61.035 65.365 ;
      RECT 60.405 65.195 60.575 65.365 ;
      RECT 59.945 65.195 60.115 65.365 ;
      RECT 59.485 65.195 59.655 65.365 ;
      RECT 59.025 65.195 59.195 65.365 ;
      RECT 58.565 65.195 58.735 65.365 ;
      RECT 58.105 65.195 58.275 65.365 ;
      RECT 57.645 65.195 57.815 65.365 ;
      RECT 57.185 65.195 57.355 65.365 ;
      RECT 56.725 65.195 56.895 65.365 ;
      RECT 56.265 65.195 56.435 65.365 ;
      RECT 55.805 65.195 55.975 65.365 ;
      RECT 55.345 65.195 55.515 65.365 ;
      RECT 54.885 65.195 55.055 65.365 ;
      RECT 54.425 65.195 54.595 65.365 ;
      RECT 53.965 65.195 54.135 65.365 ;
      RECT 53.505 65.195 53.675 65.365 ;
      RECT 53.045 65.195 53.215 65.365 ;
      RECT 52.585 65.195 52.755 65.365 ;
      RECT 52.125 65.195 52.295 65.365 ;
      RECT 51.665 65.195 51.835 65.365 ;
      RECT 51.205 65.195 51.375 65.365 ;
      RECT 50.745 65.195 50.915 65.365 ;
      RECT 50.285 65.195 50.455 65.365 ;
      RECT 49.825 65.195 49.995 65.365 ;
      RECT 49.365 65.195 49.535 65.365 ;
      RECT 48.905 65.195 49.075 65.365 ;
      RECT 48.445 65.195 48.615 65.365 ;
      RECT 47.985 65.195 48.155 65.365 ;
      RECT 47.525 65.195 47.695 65.365 ;
      RECT 47.065 65.195 47.235 65.365 ;
      RECT 46.605 65.195 46.775 65.365 ;
      RECT 46.145 65.195 46.315 65.365 ;
      RECT 45.685 65.195 45.855 65.365 ;
      RECT 45.225 65.195 45.395 65.365 ;
      RECT 44.765 65.195 44.935 65.365 ;
      RECT 44.305 65.195 44.475 65.365 ;
      RECT 43.845 65.195 44.015 65.365 ;
      RECT 43.385 65.195 43.555 65.365 ;
      RECT 42.925 65.195 43.095 65.365 ;
      RECT 42.465 65.195 42.635 65.365 ;
      RECT 42.005 65.195 42.175 65.365 ;
      RECT 41.545 65.195 41.715 65.365 ;
      RECT 41.085 65.195 41.255 65.365 ;
      RECT 40.625 65.195 40.795 65.365 ;
      RECT 40.165 65.195 40.335 65.365 ;
      RECT 39.705 65.195 39.875 65.365 ;
      RECT 39.245 65.195 39.415 65.365 ;
      RECT 38.785 65.195 38.955 65.365 ;
      RECT 38.325 65.195 38.495 65.365 ;
      RECT 37.865 65.195 38.035 65.365 ;
      RECT 37.405 65.195 37.575 65.365 ;
      RECT 36.945 65.195 37.115 65.365 ;
      RECT 36.485 65.195 36.655 65.365 ;
      RECT 36.025 65.195 36.195 65.365 ;
      RECT 35.565 65.195 35.735 65.365 ;
      RECT 35.105 65.195 35.275 65.365 ;
      RECT 34.645 65.195 34.815 65.365 ;
      RECT 34.185 65.195 34.355 65.365 ;
      RECT 33.725 65.195 33.895 65.365 ;
      RECT 33.265 65.195 33.435 65.365 ;
      RECT 32.805 65.195 32.975 65.365 ;
      RECT 32.345 65.195 32.515 65.365 ;
      RECT 31.885 65.195 32.055 65.365 ;
      RECT 31.425 65.195 31.595 65.365 ;
      RECT 30.965 65.195 31.135 65.365 ;
      RECT 30.505 65.195 30.675 65.365 ;
      RECT 30.045 65.195 30.215 65.365 ;
      RECT 29.585 65.195 29.755 65.365 ;
      RECT 29.125 65.195 29.295 65.365 ;
      RECT 28.665 65.195 28.835 65.365 ;
      RECT 28.205 65.195 28.375 65.365 ;
      RECT 27.745 65.195 27.915 65.365 ;
      RECT 27.285 65.195 27.455 65.365 ;
      RECT 26.825 65.195 26.995 65.365 ;
      RECT 26.365 65.195 26.535 65.365 ;
      RECT 25.905 65.195 26.075 65.365 ;
      RECT 25.445 65.195 25.615 65.365 ;
      RECT 24.985 65.195 25.155 65.365 ;
      RECT 24.525 65.195 24.695 65.365 ;
      RECT 24.065 65.195 24.235 65.365 ;
      RECT 23.605 65.195 23.775 65.365 ;
      RECT 23.145 65.195 23.315 65.365 ;
      RECT 22.685 65.195 22.855 65.365 ;
      RECT 22.225 65.195 22.395 65.365 ;
      RECT 21.765 65.195 21.935 65.365 ;
      RECT 21.305 65.195 21.475 65.365 ;
      RECT 20.845 65.195 21.015 65.365 ;
      RECT 20.385 65.195 20.555 65.365 ;
      RECT 19.925 65.195 20.095 65.365 ;
      RECT 19.465 65.195 19.635 65.365 ;
      RECT 19.005 65.195 19.175 65.365 ;
      RECT 18.545 65.195 18.715 65.365 ;
      RECT 18.085 65.195 18.255 65.365 ;
      RECT 17.625 65.195 17.795 65.365 ;
      RECT 17.165 65.195 17.335 65.365 ;
      RECT 16.705 65.195 16.875 65.365 ;
      RECT 16.245 65.195 16.415 65.365 ;
      RECT 15.785 65.195 15.955 65.365 ;
      RECT 15.325 65.195 15.495 65.365 ;
      RECT 14.865 65.195 15.035 65.365 ;
      RECT 14.405 65.195 14.575 65.365 ;
      RECT 13.945 65.195 14.115 65.365 ;
      RECT 13.485 65.195 13.655 65.365 ;
      RECT 13.025 65.195 13.195 65.365 ;
      RECT 12.565 65.195 12.735 65.365 ;
      RECT 12.105 65.195 12.275 65.365 ;
      RECT 11.645 65.195 11.815 65.365 ;
      RECT 11.185 65.195 11.355 65.365 ;
      RECT 10.725 65.195 10.895 65.365 ;
      RECT 10.265 65.195 10.435 65.365 ;
      RECT 9.805 65.195 9.975 65.365 ;
      RECT 9.345 65.195 9.515 65.365 ;
      RECT 8.885 65.195 9.055 65.365 ;
      RECT 8.425 65.195 8.595 65.365 ;
      RECT 7.965 65.195 8.135 65.365 ;
      RECT 7.505 65.195 7.675 65.365 ;
      RECT 7.045 65.195 7.215 65.365 ;
      RECT 6.585 65.195 6.755 65.365 ;
      RECT 6.125 65.195 6.295 65.365 ;
      RECT 5.665 65.195 5.835 65.365 ;
      RECT 5.205 65.195 5.375 65.365 ;
      RECT 4.745 65.195 4.915 65.365 ;
      RECT 4.285 65.195 4.455 65.365 ;
      RECT 3.825 65.195 3.995 65.365 ;
      RECT 3.365 65.195 3.535 65.365 ;
      RECT 2.905 65.195 3.075 65.365 ;
      RECT 2.445 65.195 2.615 65.365 ;
      RECT 1.985 65.195 2.155 65.365 ;
      RECT 1.525 65.195 1.695 65.365 ;
      RECT 1.065 65.195 1.235 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 84.325 62.475 84.495 62.645 ;
      RECT 83.865 62.475 84.035 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 84.325 59.755 84.495 59.925 ;
      RECT 83.865 59.755 84.035 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 84.325 57.035 84.495 57.205 ;
      RECT 83.865 57.035 84.035 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 84.325 54.315 84.495 54.485 ;
      RECT 83.865 54.315 84.035 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 84.325 51.595 84.495 51.765 ;
      RECT 83.865 51.595 84.035 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 84.325 48.875 84.495 49.045 ;
      RECT 83.865 48.875 84.035 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 84.325 46.155 84.495 46.325 ;
      RECT 83.865 46.155 84.035 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 84.325 43.435 84.495 43.605 ;
      RECT 83.865 43.435 84.035 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 84.325 40.715 84.495 40.885 ;
      RECT 83.865 40.715 84.035 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 84.325 37.995 84.495 38.165 ;
      RECT 83.865 37.995 84.035 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 84.325 35.275 84.495 35.445 ;
      RECT 83.865 35.275 84.035 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 84.325 32.555 84.495 32.725 ;
      RECT 83.865 32.555 84.035 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 84.325 29.835 84.495 30.005 ;
      RECT 83.865 29.835 84.035 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 84.325 27.115 84.495 27.285 ;
      RECT 83.865 27.115 84.035 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 84.325 24.395 84.495 24.565 ;
      RECT 83.865 24.395 84.035 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 84.325 21.675 84.495 21.845 ;
      RECT 83.865 21.675 84.035 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 84.325 18.955 84.495 19.125 ;
      RECT 83.865 18.955 84.035 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 84.325 16.235 84.495 16.405 ;
      RECT 83.865 16.235 84.035 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 84.325 13.515 84.495 13.685 ;
      RECT 83.865 13.515 84.035 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 84.325 10.795 84.495 10.965 ;
      RECT 83.865 10.795 84.035 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 84.325 8.075 84.495 8.245 ;
      RECT 83.865 8.075 84.035 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 84.325 5.355 84.495 5.525 ;
      RECT 83.865 5.355 84.035 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 84.325 2.635 84.495 2.805 ;
      RECT 83.865 2.635 84.035 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 73.525 81.525 73.675 81.675 ;
      RECT 44.085 81.525 44.235 81.675 ;
      RECT 49.145 79.825 49.295 79.975 ;
      RECT 73.525 65.205 73.675 65.355 ;
      RECT 44.085 65.205 44.235 65.355 ;
      RECT 4.525 63.505 4.675 63.655 ;
      RECT 3.605 63.505 3.755 63.655 ;
      RECT 2.225 1.625 2.375 1.775 ;
      RECT 73.525 -0.075 73.675 0.075 ;
      RECT 44.085 -0.075 44.235 0.075 ;
    LAYER via2 ;
      RECT 73.5 81.5 73.7 81.7 ;
      RECT 44.06 81.5 44.26 81.7 ;
      RECT 1.28 57.02 1.48 57.22 ;
      RECT 1.28 41.38 1.48 41.58 ;
      RECT 1.74 24.38 1.94 24.58 ;
      RECT 1.74 8.06 1.94 8.26 ;
      RECT 73.5 -0.1 73.7 0.1 ;
      RECT 44.06 -0.1 44.26 0.1 ;
    LAYER via3 ;
      RECT 73.5 81.5 73.7 81.7 ;
      RECT 44.06 81.5 44.26 81.7 ;
      RECT 73.5 -0.1 73.7 0.1 ;
      RECT 44.06 -0.1 44.26 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 65.28 18.4 65.28 18.4 81.6 84.64 81.6 84.64 0 ;
  END
END sb_2__0_

END LIBRARY
