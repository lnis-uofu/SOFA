VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_1__2_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 123.28 BY 97.92 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 55.59 0 55.73 1.36 ;
    END
  END prog_clk[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 71.25 123.28 71.55 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 34.53 123.28 34.83 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 73.97 123.28 74.27 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 81.45 123.28 81.75 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 35.89 123.28 36.19 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 17.53 123.28 17.83 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 40.65 123.28 40.95 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 50.17 123.28 50.47 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 76.69 123.28 76.99 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 61.05 123.28 61.35 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 72.61 123.28 72.91 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 80.09 123.28 80.39 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 57.65 123.28 57.95 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 67.85 123.28 68.15 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 54.93 123.28 55.23 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 52.89 123.28 53.19 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 59.69 123.28 59.99 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 84.17 123.28 84.47 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 75.33 123.28 75.63 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 62.41 123.28 62.71 ;
    END
  END chanx_right_in[19]
  PIN right_top_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 37.25 123.28 37.55 ;
    END
  END right_top_grid_pin_1_[0]
  PIN right_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.93 10.88 115.07 12.24 ;
    END
  END right_bottom_grid_pin_34_[0]
  PIN right_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.85 10.88 115.99 12.24 ;
    END
  END right_bottom_grid_pin_35_[0]
  PIN right_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.87 10.88 110.01 12.24 ;
    END
  END right_bottom_grid_pin_36_[0]
  PIN right_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.63 10.88 112.77 12.24 ;
    END
  END right_bottom_grid_pin_37_[0]
  PIN right_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.61 10.88 118.75 12.24 ;
    END
  END right_bottom_grid_pin_38_[0]
  PIN right_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.77 10.88 116.91 12.24 ;
    END
  END right_bottom_grid_pin_39_[0]
  PIN right_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.69 10.88 117.83 12.24 ;
    END
  END right_bottom_grid_pin_40_[0]
  PIN right_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.01 10.88 114.15 12.24 ;
    END
  END right_bottom_grid_pin_41_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.47 0 68.61 1.36 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.39 0 69.53 1.36 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.43 0 80.57 1.36 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.31 0 70.45 1.36 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.65 0 60.79 1.36 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.33 0 64.47 1.36 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.57 0 61.71 1.36 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.45 0 74.59 1.36 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.55 0 67.69 1.36 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.73 0 82.87 1.36 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.23 0 71.37 1.36 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.37 0 75.51 1.36 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.63 0 66.77 1.36 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 0 48.37 1.36 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.35 0 81.49 1.36 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.15 0 49.29 1.36 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.73 0 59.87 1.36 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.41 0 63.55 1.36 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.71 0 65.85 1.36 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.59 0 78.73 1.36 ;
    END
  END chany_bottom_in[19]
  PIN bottom_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.43 10.88 11.57 12.24 ;
    END
  END bottom_left_grid_pin_42_[0]
  PIN bottom_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.13 10.88 9.27 12.24 ;
    END
  END bottom_left_grid_pin_43_[0]
  PIN bottom_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.35 10.88 12.49 12.24 ;
    END
  END bottom_left_grid_pin_44_[0]
  PIN bottom_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.19 10.88 14.33 12.24 ;
    END
  END bottom_left_grid_pin_45_[0]
  PIN bottom_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.03 10.88 16.17 12.24 ;
    END
  END bottom_left_grid_pin_46_[0]
  PIN bottom_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.87 10.88 18.01 12.24 ;
    END
  END bottom_left_grid_pin_47_[0]
  PIN bottom_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 5.37 10.88 5.67 12.24 ;
    END
  END bottom_left_grid_pin_48_[0]
  PIN bottom_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.81 10.88 12.11 12.24 ;
    END
  END bottom_left_grid_pin_49_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.73 1.38 45.03 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 61.05 1.38 61.35 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.97 1.38 40.27 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 23.65 1.38 23.95 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.09 1.38 29.39 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.01 1.38 25.31 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 41.33 1.38 41.63 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 35.89 1.38 36.19 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.17 1.38 33.47 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 65.13 1.38 65.43 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 47.45 1.38 47.75 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 20.25 1.38 20.55 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 17.53 1.38 17.83 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.29 1.38 22.59 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 18.89 1.38 19.19 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 34.53 1.38 34.83 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 58.33 1.38 58.63 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 63.77 1.38 64.07 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.97 1.38 57.27 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 38.61 1.38 38.91 ;
    END
  END chanx_left_in[19]
  PIN left_top_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 55.61 1.38 55.91 ;
    END
  END left_top_grid_pin_1_[0]
  PIN left_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.11 10.88 15.25 12.24 ;
    END
  END left_bottom_grid_pin_34_[0]
  PIN left_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.27 10.88 13.41 12.24 ;
    END
  END left_bottom_grid_pin_35_[0]
  PIN left_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.99 10.88 5.13 12.24 ;
    END
  END left_bottom_grid_pin_36_[0]
  PIN left_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.91 10.88 6.05 12.24 ;
    END
  END left_bottom_grid_pin_37_[0]
  PIN left_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.75 10.88 7.89 12.24 ;
    END
  END left_bottom_grid_pin_38_[0]
  PIN left_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.07 10.88 4.21 12.24 ;
    END
  END left_bottom_grid_pin_39_[0]
  PIN left_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.15 10.88 3.29 12.24 ;
    END
  END left_bottom_grid_pin_40_[0]
  PIN left_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.83 10.88 6.97 12.24 ;
    END
  END left_bottom_grid_pin_41_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 42.69 123.28 42.99 ;
    END
  END ccff_head[0]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 31.81 123.28 32.11 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 33.17 123.28 33.47 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 29.09 123.28 29.39 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 30.45 123.28 30.75 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 63.77 123.28 64.07 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 19.57 123.28 19.87 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 46.09 123.28 46.39 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 27.73 123.28 28.03 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 48.13 123.28 48.43 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 24.33 123.28 24.63 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 51.53 123.28 51.83 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 22.97 123.28 23.27 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 56.29 123.28 56.59 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 26.37 123.28 26.67 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 44.05 123.28 44.35 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 38.61 123.28 38.91 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 69.89 123.28 70.19 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 82.81 123.28 83.11 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 65.81 123.28 66.11 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 21.61 123.28 21.91 ;
    END
  END chanx_right_out[19]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.89 0 58.03 1.36 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.49 0 62.63 1.36 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.81 0 58.95 1.36 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.51 0 79.65 1.36 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 0 52.97 1.36 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.79 0 87.93 1.36 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 0 50.21 1.36 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.67 0 77.81 1.36 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.49 0 85.63 1.36 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.07 0 73.21 1.36 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 0 52.05 1.36 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.75 0 76.89 1.36 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.63 0 43.77 1.36 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.71 0 88.85 1.36 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 0 51.13 1.36 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.63 0 89.77 1.36 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.57 0 84.71 1.36 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.15 0 72.29 1.36 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.97 0 57.11 1.36 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.55 0 90.69 1.36 ;
    END
  END chany_bottom_out[19]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 71.25 1.38 71.55 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 89.61 1.38 89.91 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 68.53 1.38 68.83 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 51.53 1.38 51.83 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 75.33 1.38 75.63 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 46.09 1.38 46.39 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 54.25 1.38 54.55 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.17 1.38 50.47 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 73.97 1.38 74.27 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.25 1.38 37.55 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 72.61 1.38 72.91 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 30.45 1.38 30.75 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.89 1.38 70.19 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.81 1.38 49.11 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.89 1.38 53.19 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 62.41 1.38 62.71 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.37 1.38 43.67 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 26.37 1.38 26.67 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.69 1.38 59.99 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 27.73 1.38 28.03 ;
    END
  END chanx_left_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.81 1.38 32.11 ;
    END
  END ccff_tail[0]
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.33 96.56 64.47 97.92 ;
    END
  END SC_IN_TOP
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.41 96.56 63.55 97.92 ;
    END
  END SC_IN_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.49 96.56 62.63 97.92 ;
    END
  END SC_OUT_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.57 96.56 61.71 97.92 ;
    END
  END SC_OUT_BOT
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 27.6 2.48 28.08 2.96 ;
        RECT 95.2 2.48 95.68 2.96 ;
        RECT 27.6 7.92 28.08 8.4 ;
        RECT 95.2 7.92 95.68 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 122.8 13.36 123.28 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 122.8 18.8 123.28 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 122.8 24.24 123.28 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 122.8 29.68 123.28 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 122.8 35.12 123.28 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 122.8 40.56 123.28 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 122.8 46 123.28 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 122.8 51.44 123.28 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 122.8 56.88 123.28 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 122.8 62.32 123.28 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 122.8 67.76 123.28 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 122.8 73.2 123.28 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 122.8 78.64 123.28 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 122.8 84.08 123.28 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 122.8 89.52 123.28 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 122.8 94.96 123.28 95.44 ;
      LAYER met4 ;
        RECT 39.26 0 39.86 0.6 ;
        RECT 68.7 0 69.3 0.6 ;
        RECT 112.86 10.88 113.46 11.48 ;
        RECT 39.26 97.32 39.86 97.92 ;
        RECT 68.7 97.32 69.3 97.92 ;
        RECT 112.86 97.32 113.46 97.92 ;
      LAYER met5 ;
        RECT 0 22.2 3.2 25.4 ;
        RECT 120.08 22.2 123.28 25.4 ;
        RECT 0 63 3.2 66.2 ;
        RECT 120.08 63 123.28 66.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 27.6 0 95.68 0.24 ;
        RECT 27.6 5.2 28.08 5.68 ;
        RECT 95.2 5.2 95.68 5.68 ;
        RECT 0 10.64 123.28 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 122.8 16.08 123.28 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 122.8 21.52 123.28 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 122.8 26.96 123.28 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 122.8 32.4 123.28 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 122.8 37.84 123.28 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 122.8 43.28 123.28 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 122.8 48.72 123.28 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 122.8 54.16 123.28 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 122.8 59.6 123.28 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 122.8 65.04 123.28 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 122.8 70.48 123.28 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 122.8 75.92 123.28 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 122.8 81.36 123.28 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 122.8 86.8 123.28 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 122.8 92.24 123.28 92.72 ;
        RECT 0 97.68 123.28 97.92 ;
      LAYER met4 ;
        RECT 53.98 0 54.58 0.6 ;
        RECT 83.42 0 84.02 0.6 ;
        RECT 9.82 10.88 10.42 11.48 ;
        RECT 9.82 97.32 10.42 97.92 ;
        RECT 53.98 97.32 54.58 97.92 ;
        RECT 83.42 97.32 84.02 97.92 ;
      LAYER met5 ;
        RECT 0 42.6 3.2 45.8 ;
        RECT 120.08 42.6 123.28 45.8 ;
        RECT 0 83.4 3.2 86.6 ;
        RECT 120.08 83.4 123.28 86.6 ;
    END
  END VSS
  PIN grid_clb_0_bottom_width_0_height_0__pin_50___FEEDTHRU_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.81 0 35.95 1.36 ;
    END
  END grid_clb_0_bottom_width_0_height_0__pin_50___FEEDTHRU_0[0]
  PIN grid_clb_0_bottom_width_0_height_0__pin_50___FEEDTHRU_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.9 14.13 123.28 14.43 ;
    END
  END grid_clb_0_bottom_width_0_height_0__pin_50___FEEDTHRU_1[0]
  OBS
    LAYER li1 ;
      RECT 0 97.835 123.28 98.005 ;
      RECT 122.82 95.115 123.28 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 122.82 92.395 123.28 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 122.82 89.675 123.28 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 122.82 86.955 123.28 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 122.36 84.235 123.28 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 122.36 81.515 123.28 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 122.82 78.795 123.28 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 121.44 76.075 123.28 76.245 ;
      RECT 0 76.075 1.84 76.245 ;
      RECT 119.6 73.355 123.28 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 119.6 70.635 123.28 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 122.36 67.915 123.28 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 119.6 65.195 123.28 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 119.6 62.475 123.28 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 122.36 59.755 123.28 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 122.36 57.035 123.28 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 122.36 54.315 123.28 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 122.36 51.595 123.28 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 122.36 48.875 123.28 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 122.36 46.155 123.28 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 122.36 43.435 123.28 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 122.36 40.715 123.28 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 122.36 37.995 123.28 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 122.36 35.275 123.28 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 122.36 32.555 123.28 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 122.36 29.835 123.28 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 122.36 27.115 123.28 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 122.36 24.395 123.28 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 122.36 21.675 123.28 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 122.36 18.955 123.28 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 122.36 16.235 123.28 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 122.36 13.515 123.28 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 92.92 10.795 123.28 10.965 ;
      RECT 0 10.795 29.44 10.965 ;
      RECT 94.76 8.075 95.68 8.245 ;
      RECT 27.6 8.075 29.44 8.245 ;
      RECT 94.76 5.355 95.68 5.525 ;
      RECT 27.6 5.355 31.28 5.525 ;
      RECT 95.22 2.635 95.68 2.805 ;
      RECT 27.6 2.635 31.28 2.805 ;
      RECT 27.6 -0.085 95.68 0.085 ;
    LAYER met2 ;
      RECT 83.58 97.735 83.86 98.105 ;
      RECT 54.14 97.735 54.42 98.105 ;
      RECT 9.98 97.735 10.26 98.105 ;
      RECT 9.98 10.695 10.26 11.065 ;
      RECT 62.89 1.54 63.15 1.86 ;
      RECT 61.05 1.54 61.31 1.86 ;
      RECT 83.58 -0.185 83.86 0.185 ;
      RECT 54.14 -0.185 54.42 0.185 ;
      POLYGON 123 97.64 123 11.16 119.03 11.16 119.03 12.52 118.33 12.52 118.33 11.16 118.11 11.16 118.11 12.52 117.41 12.52 117.41 11.16 117.19 11.16 117.19 12.52 116.49 12.52 116.49 11.16 116.27 11.16 116.27 12.52 115.57 12.52 115.57 11.16 115.35 11.16 115.35 12.52 114.65 12.52 114.65 11.16 114.43 11.16 114.43 12.52 113.73 12.52 113.73 11.16 113.05 11.16 113.05 12.52 112.35 12.52 112.35 11.16 110.29 11.16 110.29 12.52 109.59 12.52 109.59 11.16 95.4 11.16 95.4 0.28 90.97 0.28 90.97 1.64 90.27 1.64 90.27 0.28 90.05 0.28 90.05 1.64 89.35 1.64 89.35 0.28 89.13 0.28 89.13 1.64 88.43 1.64 88.43 0.28 88.21 0.28 88.21 1.64 87.51 1.64 87.51 0.28 85.91 0.28 85.91 1.64 85.21 1.64 85.21 0.28 84.99 0.28 84.99 1.64 84.29 1.64 84.29 0.28 83.15 0.28 83.15 1.64 82.45 1.64 82.45 0.28 81.77 0.28 81.77 1.64 81.07 1.64 81.07 0.28 80.85 0.28 80.85 1.64 80.15 1.64 80.15 0.28 79.93 0.28 79.93 1.64 79.23 1.64 79.23 0.28 79.01 0.28 79.01 1.64 78.31 1.64 78.31 0.28 78.09 0.28 78.09 1.64 77.39 1.64 77.39 0.28 77.17 0.28 77.17 1.64 76.47 1.64 76.47 0.28 75.79 0.28 75.79 1.64 75.09 1.64 75.09 0.28 74.87 0.28 74.87 1.64 74.17 1.64 74.17 0.28 73.49 0.28 73.49 1.64 72.79 1.64 72.79 0.28 72.57 0.28 72.57 1.64 71.87 1.64 71.87 0.28 71.65 0.28 71.65 1.64 70.95 1.64 70.95 0.28 70.73 0.28 70.73 1.64 70.03 1.64 70.03 0.28 69.81 0.28 69.81 1.64 69.11 1.64 69.11 0.28 68.89 0.28 68.89 1.64 68.19 1.64 68.19 0.28 67.97 0.28 67.97 1.64 67.27 1.64 67.27 0.28 67.05 0.28 67.05 1.64 66.35 1.64 66.35 0.28 66.13 0.28 66.13 1.64 65.43 1.64 65.43 0.28 64.75 0.28 64.75 1.64 64.05 1.64 64.05 0.28 63.83 0.28 63.83 1.64 63.13 1.64 63.13 0.28 62.91 0.28 62.91 1.64 62.21 1.64 62.21 0.28 61.99 0.28 61.99 1.64 61.29 1.64 61.29 0.28 61.07 0.28 61.07 1.64 60.37 1.64 60.37 0.28 60.15 0.28 60.15 1.64 59.45 1.64 59.45 0.28 59.23 0.28 59.23 1.64 58.53 1.64 58.53 0.28 58.31 0.28 58.31 1.64 57.61 1.64 57.61 0.28 57.39 0.28 57.39 1.64 56.69 1.64 56.69 0.28 56.01 0.28 56.01 1.64 55.31 1.64 55.31 0.28 53.25 0.28 53.25 1.64 52.55 1.64 52.55 0.28 52.33 0.28 52.33 1.64 51.63 1.64 51.63 0.28 51.41 0.28 51.41 1.64 50.71 1.64 50.71 0.28 50.49 0.28 50.49 1.64 49.79 1.64 49.79 0.28 49.57 0.28 49.57 1.64 48.87 1.64 48.87 0.28 48.65 0.28 48.65 1.64 47.95 1.64 47.95 0.28 44.05 0.28 44.05 1.64 43.35 1.64 43.35 0.28 36.23 0.28 36.23 1.64 35.53 1.64 35.53 0.28 27.88 0.28 27.88 11.16 18.29 11.16 18.29 12.52 17.59 12.52 17.59 11.16 16.45 11.16 16.45 12.52 15.75 12.52 15.75 11.16 15.53 11.16 15.53 12.52 14.83 12.52 14.83 11.16 14.61 11.16 14.61 12.52 13.91 12.52 13.91 11.16 13.69 11.16 13.69 12.52 12.99 12.52 12.99 11.16 12.77 11.16 12.77 12.52 12.07 12.52 12.07 11.16 11.85 11.16 11.85 12.52 11.15 12.52 11.15 11.16 9.55 11.16 9.55 12.52 8.85 12.52 8.85 11.16 8.17 11.16 8.17 12.52 7.47 12.52 7.47 11.16 7.25 11.16 7.25 12.52 6.55 12.52 6.55 11.16 6.33 11.16 6.33 12.52 5.63 12.52 5.63 11.16 5.41 11.16 5.41 12.52 4.71 12.52 4.71 11.16 4.49 11.16 4.49 12.52 3.79 12.52 3.79 11.16 3.57 11.16 3.57 12.52 2.87 12.52 2.87 11.16 0.28 11.16 0.28 97.64 61.29 97.64 61.29 96.28 61.99 96.28 61.99 97.64 62.21 97.64 62.21 96.28 62.91 96.28 62.91 97.64 63.13 97.64 63.13 96.28 63.83 96.28 63.83 97.64 64.05 97.64 64.05 96.28 64.75 96.28 64.75 97.64 ;
    LAYER met3 ;
      POLYGON 83.885 98.085 83.885 98.08 84.1 98.08 84.1 97.76 83.885 97.76 83.885 97.755 83.555 97.755 83.555 97.76 83.34 97.76 83.34 98.08 83.555 98.08 83.555 98.085 ;
      POLYGON 54.445 98.085 54.445 98.08 54.66 98.08 54.66 97.76 54.445 97.76 54.445 97.755 54.115 97.755 54.115 97.76 53.9 97.76 53.9 98.08 54.115 98.08 54.115 98.085 ;
      POLYGON 10.285 98.085 10.285 98.08 10.5 98.08 10.5 97.76 10.285 97.76 10.285 97.755 9.955 97.755 9.955 97.76 9.74 97.76 9.74 98.08 9.955 98.08 9.955 98.085 ;
      POLYGON 2.91 60.67 2.91 60.37 1.99 60.37 1.99 59.69 1.78 59.69 1.78 60.39 1.69 60.39 1.69 60.67 ;
      POLYGON 70.99 59.31 70.99 59.01 1.78 59.01 1.78 59.03 1.23 59.03 1.23 59.31 ;
      POLYGON 2.005 53.885 2.005 53.88 2.03 53.88 2.03 53.56 2.005 53.56 2.005 53.555 1.275 53.555 1.275 53.885 ;
      POLYGON 121.5 43.67 121.5 43.65 122.97 43.65 122.97 43.37 118.99 43.37 118.99 43.67 ;
      POLYGON 1.545 17.165 1.545 17.15 30.51 17.15 30.51 16.85 1.545 16.85 1.545 16.835 1.215 16.835 1.215 17.165 ;
      POLYGON 121.63 17.16 121.63 16.84 121.25 16.84 121.25 16.85 91.39 16.85 91.39 17.15 121.25 17.15 121.25 17.16 ;
      POLYGON 10.285 11.045 10.285 11.04 10.5 11.04 10.5 10.72 10.285 10.72 10.285 10.715 9.955 10.715 9.955 10.72 9.74 10.72 9.74 11.04 9.955 11.04 9.955 11.045 ;
      POLYGON 83.885 0.165 83.885 0.16 84.1 0.16 84.1 -0.16 83.885 -0.16 83.885 -0.165 83.555 -0.165 83.555 -0.16 83.34 -0.16 83.34 0.16 83.555 0.16 83.555 0.165 ;
      POLYGON 54.445 0.165 54.445 0.16 54.66 0.16 54.66 -0.16 54.445 -0.16 54.445 -0.165 54.115 -0.165 54.115 -0.16 53.9 -0.16 53.9 0.16 54.115 0.16 54.115 0.165 ;
      POLYGON 122.88 97.52 122.88 84.87 121.5 84.87 121.5 83.77 122.88 83.77 122.88 83.51 121.5 83.51 121.5 82.41 122.88 82.41 122.88 82.15 121.5 82.15 121.5 81.05 122.88 81.05 122.88 80.79 121.5 80.79 121.5 79.69 122.88 79.69 122.88 77.39 121.5 77.39 121.5 76.29 122.88 76.29 122.88 76.03 121.5 76.03 121.5 74.93 122.88 74.93 122.88 74.67 121.5 74.67 121.5 73.57 122.88 73.57 122.88 73.31 121.5 73.31 121.5 72.21 122.88 72.21 122.88 71.95 121.5 71.95 121.5 70.85 122.88 70.85 122.88 70.59 121.5 70.59 121.5 69.49 122.88 69.49 122.88 68.55 121.5 68.55 121.5 67.45 122.88 67.45 122.88 66.51 121.5 66.51 121.5 65.41 122.88 65.41 122.88 64.47 121.5 64.47 121.5 63.37 122.88 63.37 122.88 63.11 121.5 63.11 121.5 62.01 122.88 62.01 122.88 61.75 121.5 61.75 121.5 60.65 122.88 60.65 122.88 60.39 121.5 60.39 121.5 59.29 122.88 59.29 122.88 58.35 121.5 58.35 121.5 57.25 122.88 57.25 122.88 56.99 121.5 56.99 121.5 55.89 122.88 55.89 122.88 55.63 121.5 55.63 121.5 54.53 122.88 54.53 122.88 53.59 121.5 53.59 121.5 52.49 122.88 52.49 122.88 52.23 121.5 52.23 121.5 51.13 122.88 51.13 122.88 50.87 121.5 50.87 121.5 49.77 122.88 49.77 122.88 48.83 121.5 48.83 121.5 47.73 122.88 47.73 122.88 46.79 121.5 46.79 121.5 45.69 122.88 45.69 122.88 44.75 121.5 44.75 121.5 43.65 122.88 43.65 122.88 43.39 121.5 43.39 121.5 42.29 122.88 42.29 122.88 41.35 121.5 41.35 121.5 40.25 122.88 40.25 122.88 39.31 121.5 39.31 121.5 38.21 122.88 38.21 122.88 37.95 121.5 37.95 121.5 36.85 122.88 36.85 122.88 36.59 121.5 36.59 121.5 35.49 122.88 35.49 122.88 35.23 121.5 35.23 121.5 34.13 122.88 34.13 122.88 33.87 121.5 33.87 121.5 32.77 122.88 32.77 122.88 32.51 121.5 32.51 121.5 31.41 122.88 31.41 122.88 31.15 121.5 31.15 121.5 30.05 122.88 30.05 122.88 29.79 121.5 29.79 121.5 28.69 122.88 28.69 122.88 28.43 121.5 28.43 121.5 27.33 122.88 27.33 122.88 27.07 121.5 27.07 121.5 25.97 122.88 25.97 122.88 25.03 121.5 25.03 121.5 23.93 122.88 23.93 122.88 23.67 121.5 23.67 121.5 22.57 122.88 22.57 122.88 22.31 121.5 22.31 121.5 21.21 122.88 21.21 122.88 20.27 121.5 20.27 121.5 19.17 122.88 19.17 122.88 18.23 121.5 18.23 121.5 17.13 122.88 17.13 122.88 14.83 121.5 14.83 121.5 13.73 122.88 13.73 122.88 11.28 95.28 11.28 95.28 0.4 28 0.4 28 11.28 0.4 11.28 0.4 17.13 1.78 17.13 1.78 18.23 0.4 18.23 0.4 18.49 1.78 18.49 1.78 19.59 0.4 19.59 0.4 19.85 1.78 19.85 1.78 20.95 0.4 20.95 0.4 21.89 1.78 21.89 1.78 22.99 0.4 22.99 0.4 23.25 1.78 23.25 1.78 24.35 0.4 24.35 0.4 24.61 1.78 24.61 1.78 25.71 0.4 25.71 0.4 25.97 1.78 25.97 1.78 27.07 0.4 27.07 0.4 27.33 1.78 27.33 1.78 28.43 0.4 28.43 0.4 28.69 1.78 28.69 1.78 29.79 0.4 29.79 0.4 30.05 1.78 30.05 1.78 31.15 0.4 31.15 0.4 31.41 1.78 31.41 1.78 32.51 0.4 32.51 0.4 32.77 1.78 32.77 1.78 33.87 0.4 33.87 0.4 34.13 1.78 34.13 1.78 35.23 0.4 35.23 0.4 35.49 1.78 35.49 1.78 36.59 0.4 36.59 0.4 36.85 1.78 36.85 1.78 37.95 0.4 37.95 0.4 38.21 1.78 38.21 1.78 39.31 0.4 39.31 0.4 39.57 1.78 39.57 1.78 40.67 0.4 40.67 0.4 40.93 1.78 40.93 1.78 42.03 0.4 42.03 0.4 42.97 1.78 42.97 1.78 44.07 0.4 44.07 0.4 44.33 1.78 44.33 1.78 45.43 0.4 45.43 0.4 45.69 1.78 45.69 1.78 46.79 0.4 46.79 0.4 47.05 1.78 47.05 1.78 48.15 0.4 48.15 0.4 48.41 1.78 48.41 1.78 49.51 0.4 49.51 0.4 49.77 1.78 49.77 1.78 50.87 0.4 50.87 0.4 51.13 1.78 51.13 1.78 52.23 0.4 52.23 0.4 52.49 1.78 52.49 1.78 53.59 0.4 53.59 0.4 53.85 1.78 53.85 1.78 54.95 0.4 54.95 0.4 55.21 1.78 55.21 1.78 56.31 0.4 56.31 0.4 56.57 1.78 56.57 1.78 57.67 0.4 57.67 0.4 57.93 1.78 57.93 1.78 59.03 0.4 59.03 0.4 59.29 1.78 59.29 1.78 60.39 0.4 60.39 0.4 60.65 1.78 60.65 1.78 61.75 0.4 61.75 0.4 62.01 1.78 62.01 1.78 63.11 0.4 63.11 0.4 63.37 1.78 63.37 1.78 64.47 0.4 64.47 0.4 64.73 1.78 64.73 1.78 65.83 0.4 65.83 0.4 68.13 1.78 68.13 1.78 69.23 0.4 69.23 0.4 69.49 1.78 69.49 1.78 70.59 0.4 70.59 0.4 70.85 1.78 70.85 1.78 71.95 0.4 71.95 0.4 72.21 1.78 72.21 1.78 73.31 0.4 73.31 0.4 73.57 1.78 73.57 1.78 74.67 0.4 74.67 0.4 74.93 1.78 74.93 1.78 76.03 0.4 76.03 0.4 89.21 1.78 89.21 1.78 90.31 0.4 90.31 0.4 97.52 ;
    LAYER met4 ;
      POLYGON 122.88 97.52 122.88 11.28 113.86 11.28 113.86 11.88 112.46 11.88 112.46 11.28 95.28 11.28 95.28 0.4 84.42 0.4 84.42 1 83.02 1 83.02 0.4 69.7 0.4 69.7 1 68.3 1 68.3 0.4 54.98 0.4 54.98 1 53.58 1 53.58 0.4 40.26 0.4 40.26 1 38.86 1 38.86 0.4 28 0.4 28 11.28 12.51 11.28 12.51 12.64 11.41 12.64 11.41 11.28 10.82 11.28 10.82 11.88 9.42 11.88 9.42 11.28 6.07 11.28 6.07 12.64 4.97 12.64 4.97 11.28 0.4 11.28 0.4 97.52 9.42 97.52 9.42 96.92 10.82 96.92 10.82 97.52 38.86 97.52 38.86 96.92 40.26 96.92 40.26 97.52 53.58 97.52 53.58 96.92 54.98 96.92 54.98 97.52 68.3 97.52 68.3 96.92 69.7 96.92 69.7 97.52 83.02 97.52 83.02 96.92 84.42 96.92 84.42 97.52 112.46 97.52 112.46 96.92 113.86 96.92 113.86 97.52 ;
    LAYER met5 ;
      POLYGON 121.68 96.32 121.68 88.2 118.48 88.2 118.48 81.8 121.68 81.8 121.68 67.8 118.48 67.8 118.48 61.4 121.68 61.4 121.68 47.4 118.48 47.4 118.48 41 121.68 41 121.68 27 118.48 27 118.48 20.6 121.68 20.6 121.68 12.48 94.08 12.48 94.08 1.6 29.2 1.6 29.2 12.48 1.6 12.48 1.6 20.6 4.8 20.6 4.8 27 1.6 27 1.6 41 4.8 41 4.8 47.4 1.6 47.4 1.6 61.4 4.8 61.4 4.8 67.8 1.6 67.8 1.6 81.8 4.8 81.8 4.8 88.2 1.6 88.2 1.6 96.32 ;
    LAYER met1 ;
      POLYGON 123 97.4 123 95.72 122.52 95.72 122.52 94.68 123 94.68 123 93 122.52 93 122.52 91.96 123 91.96 123 90.28 122.52 90.28 122.52 89.24 123 89.24 123 87.56 122.52 87.56 122.52 86.52 123 86.52 123 84.84 122.52 84.84 122.52 83.8 123 83.8 123 82.12 122.52 82.12 122.52 81.08 123 81.08 123 79.4 122.52 79.4 122.52 78.36 123 78.36 123 76.68 122.52 76.68 122.52 75.64 123 75.64 123 73.96 122.52 73.96 122.52 72.92 123 72.92 123 71.24 122.52 71.24 122.52 70.2 123 70.2 123 68.52 122.52 68.52 122.52 67.48 123 67.48 123 65.8 122.52 65.8 122.52 64.76 123 64.76 123 63.08 122.52 63.08 122.52 62.04 123 62.04 123 60.36 122.52 60.36 122.52 59.32 123 59.32 123 57.64 122.52 57.64 122.52 56.6 123 56.6 123 54.92 122.52 54.92 122.52 53.88 123 53.88 123 52.2 122.52 52.2 122.52 51.16 123 51.16 123 49.48 122.52 49.48 122.52 48.44 123 48.44 123 46.76 122.52 46.76 122.52 45.72 123 45.72 123 44.04 122.52 44.04 122.52 43 123 43 123 41.32 122.52 41.32 122.52 40.28 123 40.28 123 38.6 122.52 38.6 122.52 37.56 123 37.56 123 35.88 122.52 35.88 122.52 34.84 123 34.84 123 33.16 122.52 33.16 122.52 32.12 123 32.12 123 30.44 122.52 30.44 122.52 29.4 123 29.4 123 27.72 122.52 27.72 122.52 26.68 123 26.68 123 25 122.52 25 122.52 23.96 123 23.96 123 22.28 122.52 22.28 122.52 21.24 123 21.24 123 19.56 122.52 19.56 122.52 18.52 123 18.52 123 16.84 122.52 16.84 122.52 15.8 123 15.8 123 14.12 122.52 14.12 122.52 13.08 123 13.08 123 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 ;
      POLYGON 95.4 10.36 95.4 8.68 94.92 8.68 94.92 7.64 95.4 7.64 95.4 5.96 94.92 5.96 94.92 4.92 95.4 4.92 95.4 3.24 94.92 3.24 94.92 2.2 95.4 2.2 95.4 0.52 27.88 0.52 27.88 2.2 28.36 2.2 28.36 3.24 27.88 3.24 27.88 4.92 28.36 4.92 28.36 5.96 27.88 5.96 27.88 7.64 28.36 7.64 28.36 8.68 27.88 8.68 27.88 10.36 ;
    LAYER li1 ;
      POLYGON 123.11 97.75 123.11 11.05 95.51 11.05 95.51 0.17 27.77 0.17 27.77 11.05 0.17 11.05 0.17 97.75 ;
    LAYER mcon ;
      RECT 122.965 97.835 123.135 98.005 ;
      RECT 122.505 97.835 122.675 98.005 ;
      RECT 122.045 97.835 122.215 98.005 ;
      RECT 121.585 97.835 121.755 98.005 ;
      RECT 121.125 97.835 121.295 98.005 ;
      RECT 120.665 97.835 120.835 98.005 ;
      RECT 120.205 97.835 120.375 98.005 ;
      RECT 119.745 97.835 119.915 98.005 ;
      RECT 119.285 97.835 119.455 98.005 ;
      RECT 118.825 97.835 118.995 98.005 ;
      RECT 118.365 97.835 118.535 98.005 ;
      RECT 117.905 97.835 118.075 98.005 ;
      RECT 117.445 97.835 117.615 98.005 ;
      RECT 116.985 97.835 117.155 98.005 ;
      RECT 116.525 97.835 116.695 98.005 ;
      RECT 116.065 97.835 116.235 98.005 ;
      RECT 115.605 97.835 115.775 98.005 ;
      RECT 115.145 97.835 115.315 98.005 ;
      RECT 114.685 97.835 114.855 98.005 ;
      RECT 114.225 97.835 114.395 98.005 ;
      RECT 113.765 97.835 113.935 98.005 ;
      RECT 113.305 97.835 113.475 98.005 ;
      RECT 112.845 97.835 113.015 98.005 ;
      RECT 112.385 97.835 112.555 98.005 ;
      RECT 111.925 97.835 112.095 98.005 ;
      RECT 111.465 97.835 111.635 98.005 ;
      RECT 111.005 97.835 111.175 98.005 ;
      RECT 110.545 97.835 110.715 98.005 ;
      RECT 110.085 97.835 110.255 98.005 ;
      RECT 109.625 97.835 109.795 98.005 ;
      RECT 109.165 97.835 109.335 98.005 ;
      RECT 108.705 97.835 108.875 98.005 ;
      RECT 108.245 97.835 108.415 98.005 ;
      RECT 107.785 97.835 107.955 98.005 ;
      RECT 107.325 97.835 107.495 98.005 ;
      RECT 106.865 97.835 107.035 98.005 ;
      RECT 106.405 97.835 106.575 98.005 ;
      RECT 105.945 97.835 106.115 98.005 ;
      RECT 105.485 97.835 105.655 98.005 ;
      RECT 105.025 97.835 105.195 98.005 ;
      RECT 104.565 97.835 104.735 98.005 ;
      RECT 104.105 97.835 104.275 98.005 ;
      RECT 103.645 97.835 103.815 98.005 ;
      RECT 103.185 97.835 103.355 98.005 ;
      RECT 102.725 97.835 102.895 98.005 ;
      RECT 102.265 97.835 102.435 98.005 ;
      RECT 101.805 97.835 101.975 98.005 ;
      RECT 101.345 97.835 101.515 98.005 ;
      RECT 100.885 97.835 101.055 98.005 ;
      RECT 100.425 97.835 100.595 98.005 ;
      RECT 99.965 97.835 100.135 98.005 ;
      RECT 99.505 97.835 99.675 98.005 ;
      RECT 99.045 97.835 99.215 98.005 ;
      RECT 98.585 97.835 98.755 98.005 ;
      RECT 98.125 97.835 98.295 98.005 ;
      RECT 97.665 97.835 97.835 98.005 ;
      RECT 97.205 97.835 97.375 98.005 ;
      RECT 96.745 97.835 96.915 98.005 ;
      RECT 96.285 97.835 96.455 98.005 ;
      RECT 95.825 97.835 95.995 98.005 ;
      RECT 95.365 97.835 95.535 98.005 ;
      RECT 94.905 97.835 95.075 98.005 ;
      RECT 94.445 97.835 94.615 98.005 ;
      RECT 93.985 97.835 94.155 98.005 ;
      RECT 93.525 97.835 93.695 98.005 ;
      RECT 93.065 97.835 93.235 98.005 ;
      RECT 92.605 97.835 92.775 98.005 ;
      RECT 92.145 97.835 92.315 98.005 ;
      RECT 91.685 97.835 91.855 98.005 ;
      RECT 91.225 97.835 91.395 98.005 ;
      RECT 90.765 97.835 90.935 98.005 ;
      RECT 90.305 97.835 90.475 98.005 ;
      RECT 89.845 97.835 90.015 98.005 ;
      RECT 89.385 97.835 89.555 98.005 ;
      RECT 88.925 97.835 89.095 98.005 ;
      RECT 88.465 97.835 88.635 98.005 ;
      RECT 88.005 97.835 88.175 98.005 ;
      RECT 87.545 97.835 87.715 98.005 ;
      RECT 87.085 97.835 87.255 98.005 ;
      RECT 86.625 97.835 86.795 98.005 ;
      RECT 86.165 97.835 86.335 98.005 ;
      RECT 85.705 97.835 85.875 98.005 ;
      RECT 85.245 97.835 85.415 98.005 ;
      RECT 84.785 97.835 84.955 98.005 ;
      RECT 84.325 97.835 84.495 98.005 ;
      RECT 83.865 97.835 84.035 98.005 ;
      RECT 83.405 97.835 83.575 98.005 ;
      RECT 82.945 97.835 83.115 98.005 ;
      RECT 82.485 97.835 82.655 98.005 ;
      RECT 82.025 97.835 82.195 98.005 ;
      RECT 81.565 97.835 81.735 98.005 ;
      RECT 81.105 97.835 81.275 98.005 ;
      RECT 80.645 97.835 80.815 98.005 ;
      RECT 80.185 97.835 80.355 98.005 ;
      RECT 79.725 97.835 79.895 98.005 ;
      RECT 79.265 97.835 79.435 98.005 ;
      RECT 78.805 97.835 78.975 98.005 ;
      RECT 78.345 97.835 78.515 98.005 ;
      RECT 77.885 97.835 78.055 98.005 ;
      RECT 77.425 97.835 77.595 98.005 ;
      RECT 76.965 97.835 77.135 98.005 ;
      RECT 76.505 97.835 76.675 98.005 ;
      RECT 76.045 97.835 76.215 98.005 ;
      RECT 75.585 97.835 75.755 98.005 ;
      RECT 75.125 97.835 75.295 98.005 ;
      RECT 74.665 97.835 74.835 98.005 ;
      RECT 74.205 97.835 74.375 98.005 ;
      RECT 73.745 97.835 73.915 98.005 ;
      RECT 73.285 97.835 73.455 98.005 ;
      RECT 72.825 97.835 72.995 98.005 ;
      RECT 72.365 97.835 72.535 98.005 ;
      RECT 71.905 97.835 72.075 98.005 ;
      RECT 71.445 97.835 71.615 98.005 ;
      RECT 70.985 97.835 71.155 98.005 ;
      RECT 70.525 97.835 70.695 98.005 ;
      RECT 70.065 97.835 70.235 98.005 ;
      RECT 69.605 97.835 69.775 98.005 ;
      RECT 69.145 97.835 69.315 98.005 ;
      RECT 68.685 97.835 68.855 98.005 ;
      RECT 68.225 97.835 68.395 98.005 ;
      RECT 67.765 97.835 67.935 98.005 ;
      RECT 67.305 97.835 67.475 98.005 ;
      RECT 66.845 97.835 67.015 98.005 ;
      RECT 66.385 97.835 66.555 98.005 ;
      RECT 65.925 97.835 66.095 98.005 ;
      RECT 65.465 97.835 65.635 98.005 ;
      RECT 65.005 97.835 65.175 98.005 ;
      RECT 64.545 97.835 64.715 98.005 ;
      RECT 64.085 97.835 64.255 98.005 ;
      RECT 63.625 97.835 63.795 98.005 ;
      RECT 63.165 97.835 63.335 98.005 ;
      RECT 62.705 97.835 62.875 98.005 ;
      RECT 62.245 97.835 62.415 98.005 ;
      RECT 61.785 97.835 61.955 98.005 ;
      RECT 61.325 97.835 61.495 98.005 ;
      RECT 60.865 97.835 61.035 98.005 ;
      RECT 60.405 97.835 60.575 98.005 ;
      RECT 59.945 97.835 60.115 98.005 ;
      RECT 59.485 97.835 59.655 98.005 ;
      RECT 59.025 97.835 59.195 98.005 ;
      RECT 58.565 97.835 58.735 98.005 ;
      RECT 58.105 97.835 58.275 98.005 ;
      RECT 57.645 97.835 57.815 98.005 ;
      RECT 57.185 97.835 57.355 98.005 ;
      RECT 56.725 97.835 56.895 98.005 ;
      RECT 56.265 97.835 56.435 98.005 ;
      RECT 55.805 97.835 55.975 98.005 ;
      RECT 55.345 97.835 55.515 98.005 ;
      RECT 54.885 97.835 55.055 98.005 ;
      RECT 54.425 97.835 54.595 98.005 ;
      RECT 53.965 97.835 54.135 98.005 ;
      RECT 53.505 97.835 53.675 98.005 ;
      RECT 53.045 97.835 53.215 98.005 ;
      RECT 52.585 97.835 52.755 98.005 ;
      RECT 52.125 97.835 52.295 98.005 ;
      RECT 51.665 97.835 51.835 98.005 ;
      RECT 51.205 97.835 51.375 98.005 ;
      RECT 50.745 97.835 50.915 98.005 ;
      RECT 50.285 97.835 50.455 98.005 ;
      RECT 49.825 97.835 49.995 98.005 ;
      RECT 49.365 97.835 49.535 98.005 ;
      RECT 48.905 97.835 49.075 98.005 ;
      RECT 48.445 97.835 48.615 98.005 ;
      RECT 47.985 97.835 48.155 98.005 ;
      RECT 47.525 97.835 47.695 98.005 ;
      RECT 47.065 97.835 47.235 98.005 ;
      RECT 46.605 97.835 46.775 98.005 ;
      RECT 46.145 97.835 46.315 98.005 ;
      RECT 45.685 97.835 45.855 98.005 ;
      RECT 45.225 97.835 45.395 98.005 ;
      RECT 44.765 97.835 44.935 98.005 ;
      RECT 44.305 97.835 44.475 98.005 ;
      RECT 43.845 97.835 44.015 98.005 ;
      RECT 43.385 97.835 43.555 98.005 ;
      RECT 42.925 97.835 43.095 98.005 ;
      RECT 42.465 97.835 42.635 98.005 ;
      RECT 42.005 97.835 42.175 98.005 ;
      RECT 41.545 97.835 41.715 98.005 ;
      RECT 41.085 97.835 41.255 98.005 ;
      RECT 40.625 97.835 40.795 98.005 ;
      RECT 40.165 97.835 40.335 98.005 ;
      RECT 39.705 97.835 39.875 98.005 ;
      RECT 39.245 97.835 39.415 98.005 ;
      RECT 38.785 97.835 38.955 98.005 ;
      RECT 38.325 97.835 38.495 98.005 ;
      RECT 37.865 97.835 38.035 98.005 ;
      RECT 37.405 97.835 37.575 98.005 ;
      RECT 36.945 97.835 37.115 98.005 ;
      RECT 36.485 97.835 36.655 98.005 ;
      RECT 36.025 97.835 36.195 98.005 ;
      RECT 35.565 97.835 35.735 98.005 ;
      RECT 35.105 97.835 35.275 98.005 ;
      RECT 34.645 97.835 34.815 98.005 ;
      RECT 34.185 97.835 34.355 98.005 ;
      RECT 33.725 97.835 33.895 98.005 ;
      RECT 33.265 97.835 33.435 98.005 ;
      RECT 32.805 97.835 32.975 98.005 ;
      RECT 32.345 97.835 32.515 98.005 ;
      RECT 31.885 97.835 32.055 98.005 ;
      RECT 31.425 97.835 31.595 98.005 ;
      RECT 30.965 97.835 31.135 98.005 ;
      RECT 30.505 97.835 30.675 98.005 ;
      RECT 30.045 97.835 30.215 98.005 ;
      RECT 29.585 97.835 29.755 98.005 ;
      RECT 29.125 97.835 29.295 98.005 ;
      RECT 28.665 97.835 28.835 98.005 ;
      RECT 28.205 97.835 28.375 98.005 ;
      RECT 27.745 97.835 27.915 98.005 ;
      RECT 27.285 97.835 27.455 98.005 ;
      RECT 26.825 97.835 26.995 98.005 ;
      RECT 26.365 97.835 26.535 98.005 ;
      RECT 25.905 97.835 26.075 98.005 ;
      RECT 25.445 97.835 25.615 98.005 ;
      RECT 24.985 97.835 25.155 98.005 ;
      RECT 24.525 97.835 24.695 98.005 ;
      RECT 24.065 97.835 24.235 98.005 ;
      RECT 23.605 97.835 23.775 98.005 ;
      RECT 23.145 97.835 23.315 98.005 ;
      RECT 22.685 97.835 22.855 98.005 ;
      RECT 22.225 97.835 22.395 98.005 ;
      RECT 21.765 97.835 21.935 98.005 ;
      RECT 21.305 97.835 21.475 98.005 ;
      RECT 20.845 97.835 21.015 98.005 ;
      RECT 20.385 97.835 20.555 98.005 ;
      RECT 19.925 97.835 20.095 98.005 ;
      RECT 19.465 97.835 19.635 98.005 ;
      RECT 19.005 97.835 19.175 98.005 ;
      RECT 18.545 97.835 18.715 98.005 ;
      RECT 18.085 97.835 18.255 98.005 ;
      RECT 17.625 97.835 17.795 98.005 ;
      RECT 17.165 97.835 17.335 98.005 ;
      RECT 16.705 97.835 16.875 98.005 ;
      RECT 16.245 97.835 16.415 98.005 ;
      RECT 15.785 97.835 15.955 98.005 ;
      RECT 15.325 97.835 15.495 98.005 ;
      RECT 14.865 97.835 15.035 98.005 ;
      RECT 14.405 97.835 14.575 98.005 ;
      RECT 13.945 97.835 14.115 98.005 ;
      RECT 13.485 97.835 13.655 98.005 ;
      RECT 13.025 97.835 13.195 98.005 ;
      RECT 12.565 97.835 12.735 98.005 ;
      RECT 12.105 97.835 12.275 98.005 ;
      RECT 11.645 97.835 11.815 98.005 ;
      RECT 11.185 97.835 11.355 98.005 ;
      RECT 10.725 97.835 10.895 98.005 ;
      RECT 10.265 97.835 10.435 98.005 ;
      RECT 9.805 97.835 9.975 98.005 ;
      RECT 9.345 97.835 9.515 98.005 ;
      RECT 8.885 97.835 9.055 98.005 ;
      RECT 8.425 97.835 8.595 98.005 ;
      RECT 7.965 97.835 8.135 98.005 ;
      RECT 7.505 97.835 7.675 98.005 ;
      RECT 7.045 97.835 7.215 98.005 ;
      RECT 6.585 97.835 6.755 98.005 ;
      RECT 6.125 97.835 6.295 98.005 ;
      RECT 5.665 97.835 5.835 98.005 ;
      RECT 5.205 97.835 5.375 98.005 ;
      RECT 4.745 97.835 4.915 98.005 ;
      RECT 4.285 97.835 4.455 98.005 ;
      RECT 3.825 97.835 3.995 98.005 ;
      RECT 3.365 97.835 3.535 98.005 ;
      RECT 2.905 97.835 3.075 98.005 ;
      RECT 2.445 97.835 2.615 98.005 ;
      RECT 1.985 97.835 2.155 98.005 ;
      RECT 1.525 97.835 1.695 98.005 ;
      RECT 1.065 97.835 1.235 98.005 ;
      RECT 0.605 97.835 0.775 98.005 ;
      RECT 0.145 97.835 0.315 98.005 ;
      RECT 122.965 95.115 123.135 95.285 ;
      RECT 122.505 95.115 122.675 95.285 ;
      RECT 0.605 95.115 0.775 95.285 ;
      RECT 0.145 95.115 0.315 95.285 ;
      RECT 122.965 92.395 123.135 92.565 ;
      RECT 122.505 92.395 122.675 92.565 ;
      RECT 0.605 92.395 0.775 92.565 ;
      RECT 0.145 92.395 0.315 92.565 ;
      RECT 122.965 89.675 123.135 89.845 ;
      RECT 122.505 89.675 122.675 89.845 ;
      RECT 0.605 89.675 0.775 89.845 ;
      RECT 0.145 89.675 0.315 89.845 ;
      RECT 122.965 86.955 123.135 87.125 ;
      RECT 122.505 86.955 122.675 87.125 ;
      RECT 0.605 86.955 0.775 87.125 ;
      RECT 0.145 86.955 0.315 87.125 ;
      RECT 122.965 84.235 123.135 84.405 ;
      RECT 122.505 84.235 122.675 84.405 ;
      RECT 0.605 84.235 0.775 84.405 ;
      RECT 0.145 84.235 0.315 84.405 ;
      RECT 122.965 81.515 123.135 81.685 ;
      RECT 122.505 81.515 122.675 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 122.965 78.795 123.135 78.965 ;
      RECT 122.505 78.795 122.675 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 122.965 76.075 123.135 76.245 ;
      RECT 122.505 76.075 122.675 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 122.965 73.355 123.135 73.525 ;
      RECT 122.505 73.355 122.675 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 122.965 70.635 123.135 70.805 ;
      RECT 122.505 70.635 122.675 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 122.965 67.915 123.135 68.085 ;
      RECT 122.505 67.915 122.675 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 122.965 65.195 123.135 65.365 ;
      RECT 122.505 65.195 122.675 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 122.965 62.475 123.135 62.645 ;
      RECT 122.505 62.475 122.675 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 122.965 59.755 123.135 59.925 ;
      RECT 122.505 59.755 122.675 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 122.965 57.035 123.135 57.205 ;
      RECT 122.505 57.035 122.675 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 122.965 54.315 123.135 54.485 ;
      RECT 122.505 54.315 122.675 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 122.965 51.595 123.135 51.765 ;
      RECT 122.505 51.595 122.675 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 122.965 48.875 123.135 49.045 ;
      RECT 122.505 48.875 122.675 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 122.965 46.155 123.135 46.325 ;
      RECT 122.505 46.155 122.675 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 122.965 43.435 123.135 43.605 ;
      RECT 122.505 43.435 122.675 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 122.965 40.715 123.135 40.885 ;
      RECT 122.505 40.715 122.675 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 122.965 37.995 123.135 38.165 ;
      RECT 122.505 37.995 122.675 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 122.965 35.275 123.135 35.445 ;
      RECT 122.505 35.275 122.675 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 122.965 32.555 123.135 32.725 ;
      RECT 122.505 32.555 122.675 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 122.965 29.835 123.135 30.005 ;
      RECT 122.505 29.835 122.675 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 122.965 27.115 123.135 27.285 ;
      RECT 122.505 27.115 122.675 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 122.965 24.395 123.135 24.565 ;
      RECT 122.505 24.395 122.675 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 122.965 21.675 123.135 21.845 ;
      RECT 122.505 21.675 122.675 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 122.965 18.955 123.135 19.125 ;
      RECT 122.505 18.955 122.675 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 122.965 16.235 123.135 16.405 ;
      RECT 122.505 16.235 122.675 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 122.965 13.515 123.135 13.685 ;
      RECT 122.505 13.515 122.675 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 122.965 10.795 123.135 10.965 ;
      RECT 122.505 10.795 122.675 10.965 ;
      RECT 122.045 10.795 122.215 10.965 ;
      RECT 121.585 10.795 121.755 10.965 ;
      RECT 121.125 10.795 121.295 10.965 ;
      RECT 120.665 10.795 120.835 10.965 ;
      RECT 120.205 10.795 120.375 10.965 ;
      RECT 119.745 10.795 119.915 10.965 ;
      RECT 119.285 10.795 119.455 10.965 ;
      RECT 118.825 10.795 118.995 10.965 ;
      RECT 118.365 10.795 118.535 10.965 ;
      RECT 117.905 10.795 118.075 10.965 ;
      RECT 117.445 10.795 117.615 10.965 ;
      RECT 116.985 10.795 117.155 10.965 ;
      RECT 116.525 10.795 116.695 10.965 ;
      RECT 116.065 10.795 116.235 10.965 ;
      RECT 115.605 10.795 115.775 10.965 ;
      RECT 115.145 10.795 115.315 10.965 ;
      RECT 114.685 10.795 114.855 10.965 ;
      RECT 114.225 10.795 114.395 10.965 ;
      RECT 113.765 10.795 113.935 10.965 ;
      RECT 113.305 10.795 113.475 10.965 ;
      RECT 112.845 10.795 113.015 10.965 ;
      RECT 112.385 10.795 112.555 10.965 ;
      RECT 111.925 10.795 112.095 10.965 ;
      RECT 111.465 10.795 111.635 10.965 ;
      RECT 111.005 10.795 111.175 10.965 ;
      RECT 110.545 10.795 110.715 10.965 ;
      RECT 110.085 10.795 110.255 10.965 ;
      RECT 109.625 10.795 109.795 10.965 ;
      RECT 109.165 10.795 109.335 10.965 ;
      RECT 108.705 10.795 108.875 10.965 ;
      RECT 108.245 10.795 108.415 10.965 ;
      RECT 107.785 10.795 107.955 10.965 ;
      RECT 107.325 10.795 107.495 10.965 ;
      RECT 106.865 10.795 107.035 10.965 ;
      RECT 106.405 10.795 106.575 10.965 ;
      RECT 105.945 10.795 106.115 10.965 ;
      RECT 105.485 10.795 105.655 10.965 ;
      RECT 105.025 10.795 105.195 10.965 ;
      RECT 104.565 10.795 104.735 10.965 ;
      RECT 104.105 10.795 104.275 10.965 ;
      RECT 103.645 10.795 103.815 10.965 ;
      RECT 103.185 10.795 103.355 10.965 ;
      RECT 102.725 10.795 102.895 10.965 ;
      RECT 102.265 10.795 102.435 10.965 ;
      RECT 101.805 10.795 101.975 10.965 ;
      RECT 101.345 10.795 101.515 10.965 ;
      RECT 100.885 10.795 101.055 10.965 ;
      RECT 100.425 10.795 100.595 10.965 ;
      RECT 99.965 10.795 100.135 10.965 ;
      RECT 99.505 10.795 99.675 10.965 ;
      RECT 99.045 10.795 99.215 10.965 ;
      RECT 98.585 10.795 98.755 10.965 ;
      RECT 98.125 10.795 98.295 10.965 ;
      RECT 97.665 10.795 97.835 10.965 ;
      RECT 97.205 10.795 97.375 10.965 ;
      RECT 96.745 10.795 96.915 10.965 ;
      RECT 96.285 10.795 96.455 10.965 ;
      RECT 95.825 10.795 95.995 10.965 ;
      RECT 95.365 10.795 95.535 10.965 ;
      RECT 94.905 10.795 95.075 10.965 ;
      RECT 94.445 10.795 94.615 10.965 ;
      RECT 93.985 10.795 94.155 10.965 ;
      RECT 93.525 10.795 93.695 10.965 ;
      RECT 93.065 10.795 93.235 10.965 ;
      RECT 92.605 10.795 92.775 10.965 ;
      RECT 92.145 10.795 92.315 10.965 ;
      RECT 91.685 10.795 91.855 10.965 ;
      RECT 91.225 10.795 91.395 10.965 ;
      RECT 90.765 10.795 90.935 10.965 ;
      RECT 90.305 10.795 90.475 10.965 ;
      RECT 89.845 10.795 90.015 10.965 ;
      RECT 89.385 10.795 89.555 10.965 ;
      RECT 88.925 10.795 89.095 10.965 ;
      RECT 88.465 10.795 88.635 10.965 ;
      RECT 88.005 10.795 88.175 10.965 ;
      RECT 87.545 10.795 87.715 10.965 ;
      RECT 87.085 10.795 87.255 10.965 ;
      RECT 86.625 10.795 86.795 10.965 ;
      RECT 86.165 10.795 86.335 10.965 ;
      RECT 85.705 10.795 85.875 10.965 ;
      RECT 85.245 10.795 85.415 10.965 ;
      RECT 84.785 10.795 84.955 10.965 ;
      RECT 84.325 10.795 84.495 10.965 ;
      RECT 83.865 10.795 84.035 10.965 ;
      RECT 83.405 10.795 83.575 10.965 ;
      RECT 82.945 10.795 83.115 10.965 ;
      RECT 82.485 10.795 82.655 10.965 ;
      RECT 82.025 10.795 82.195 10.965 ;
      RECT 81.565 10.795 81.735 10.965 ;
      RECT 81.105 10.795 81.275 10.965 ;
      RECT 80.645 10.795 80.815 10.965 ;
      RECT 80.185 10.795 80.355 10.965 ;
      RECT 79.725 10.795 79.895 10.965 ;
      RECT 79.265 10.795 79.435 10.965 ;
      RECT 78.805 10.795 78.975 10.965 ;
      RECT 78.345 10.795 78.515 10.965 ;
      RECT 77.885 10.795 78.055 10.965 ;
      RECT 77.425 10.795 77.595 10.965 ;
      RECT 76.965 10.795 77.135 10.965 ;
      RECT 76.505 10.795 76.675 10.965 ;
      RECT 76.045 10.795 76.215 10.965 ;
      RECT 75.585 10.795 75.755 10.965 ;
      RECT 75.125 10.795 75.295 10.965 ;
      RECT 74.665 10.795 74.835 10.965 ;
      RECT 74.205 10.795 74.375 10.965 ;
      RECT 73.745 10.795 73.915 10.965 ;
      RECT 73.285 10.795 73.455 10.965 ;
      RECT 72.825 10.795 72.995 10.965 ;
      RECT 72.365 10.795 72.535 10.965 ;
      RECT 71.905 10.795 72.075 10.965 ;
      RECT 71.445 10.795 71.615 10.965 ;
      RECT 70.985 10.795 71.155 10.965 ;
      RECT 70.525 10.795 70.695 10.965 ;
      RECT 70.065 10.795 70.235 10.965 ;
      RECT 69.605 10.795 69.775 10.965 ;
      RECT 69.145 10.795 69.315 10.965 ;
      RECT 68.685 10.795 68.855 10.965 ;
      RECT 68.225 10.795 68.395 10.965 ;
      RECT 67.765 10.795 67.935 10.965 ;
      RECT 67.305 10.795 67.475 10.965 ;
      RECT 66.845 10.795 67.015 10.965 ;
      RECT 66.385 10.795 66.555 10.965 ;
      RECT 65.925 10.795 66.095 10.965 ;
      RECT 65.465 10.795 65.635 10.965 ;
      RECT 65.005 10.795 65.175 10.965 ;
      RECT 64.545 10.795 64.715 10.965 ;
      RECT 64.085 10.795 64.255 10.965 ;
      RECT 63.625 10.795 63.795 10.965 ;
      RECT 63.165 10.795 63.335 10.965 ;
      RECT 62.705 10.795 62.875 10.965 ;
      RECT 62.245 10.795 62.415 10.965 ;
      RECT 61.785 10.795 61.955 10.965 ;
      RECT 61.325 10.795 61.495 10.965 ;
      RECT 60.865 10.795 61.035 10.965 ;
      RECT 60.405 10.795 60.575 10.965 ;
      RECT 59.945 10.795 60.115 10.965 ;
      RECT 59.485 10.795 59.655 10.965 ;
      RECT 59.025 10.795 59.195 10.965 ;
      RECT 58.565 10.795 58.735 10.965 ;
      RECT 58.105 10.795 58.275 10.965 ;
      RECT 57.645 10.795 57.815 10.965 ;
      RECT 57.185 10.795 57.355 10.965 ;
      RECT 56.725 10.795 56.895 10.965 ;
      RECT 56.265 10.795 56.435 10.965 ;
      RECT 55.805 10.795 55.975 10.965 ;
      RECT 55.345 10.795 55.515 10.965 ;
      RECT 54.885 10.795 55.055 10.965 ;
      RECT 54.425 10.795 54.595 10.965 ;
      RECT 53.965 10.795 54.135 10.965 ;
      RECT 53.505 10.795 53.675 10.965 ;
      RECT 53.045 10.795 53.215 10.965 ;
      RECT 52.585 10.795 52.755 10.965 ;
      RECT 52.125 10.795 52.295 10.965 ;
      RECT 51.665 10.795 51.835 10.965 ;
      RECT 51.205 10.795 51.375 10.965 ;
      RECT 50.745 10.795 50.915 10.965 ;
      RECT 50.285 10.795 50.455 10.965 ;
      RECT 49.825 10.795 49.995 10.965 ;
      RECT 49.365 10.795 49.535 10.965 ;
      RECT 48.905 10.795 49.075 10.965 ;
      RECT 48.445 10.795 48.615 10.965 ;
      RECT 47.985 10.795 48.155 10.965 ;
      RECT 47.525 10.795 47.695 10.965 ;
      RECT 47.065 10.795 47.235 10.965 ;
      RECT 46.605 10.795 46.775 10.965 ;
      RECT 46.145 10.795 46.315 10.965 ;
      RECT 45.685 10.795 45.855 10.965 ;
      RECT 45.225 10.795 45.395 10.965 ;
      RECT 44.765 10.795 44.935 10.965 ;
      RECT 44.305 10.795 44.475 10.965 ;
      RECT 43.845 10.795 44.015 10.965 ;
      RECT 43.385 10.795 43.555 10.965 ;
      RECT 42.925 10.795 43.095 10.965 ;
      RECT 42.465 10.795 42.635 10.965 ;
      RECT 42.005 10.795 42.175 10.965 ;
      RECT 41.545 10.795 41.715 10.965 ;
      RECT 41.085 10.795 41.255 10.965 ;
      RECT 40.625 10.795 40.795 10.965 ;
      RECT 40.165 10.795 40.335 10.965 ;
      RECT 39.705 10.795 39.875 10.965 ;
      RECT 39.245 10.795 39.415 10.965 ;
      RECT 38.785 10.795 38.955 10.965 ;
      RECT 38.325 10.795 38.495 10.965 ;
      RECT 37.865 10.795 38.035 10.965 ;
      RECT 37.405 10.795 37.575 10.965 ;
      RECT 36.945 10.795 37.115 10.965 ;
      RECT 36.485 10.795 36.655 10.965 ;
      RECT 36.025 10.795 36.195 10.965 ;
      RECT 35.565 10.795 35.735 10.965 ;
      RECT 35.105 10.795 35.275 10.965 ;
      RECT 34.645 10.795 34.815 10.965 ;
      RECT 34.185 10.795 34.355 10.965 ;
      RECT 33.725 10.795 33.895 10.965 ;
      RECT 33.265 10.795 33.435 10.965 ;
      RECT 32.805 10.795 32.975 10.965 ;
      RECT 32.345 10.795 32.515 10.965 ;
      RECT 31.885 10.795 32.055 10.965 ;
      RECT 31.425 10.795 31.595 10.965 ;
      RECT 30.965 10.795 31.135 10.965 ;
      RECT 30.505 10.795 30.675 10.965 ;
      RECT 30.045 10.795 30.215 10.965 ;
      RECT 29.585 10.795 29.755 10.965 ;
      RECT 29.125 10.795 29.295 10.965 ;
      RECT 28.665 10.795 28.835 10.965 ;
      RECT 28.205 10.795 28.375 10.965 ;
      RECT 27.745 10.795 27.915 10.965 ;
      RECT 27.285 10.795 27.455 10.965 ;
      RECT 26.825 10.795 26.995 10.965 ;
      RECT 26.365 10.795 26.535 10.965 ;
      RECT 25.905 10.795 26.075 10.965 ;
      RECT 25.445 10.795 25.615 10.965 ;
      RECT 24.985 10.795 25.155 10.965 ;
      RECT 24.525 10.795 24.695 10.965 ;
      RECT 24.065 10.795 24.235 10.965 ;
      RECT 23.605 10.795 23.775 10.965 ;
      RECT 23.145 10.795 23.315 10.965 ;
      RECT 22.685 10.795 22.855 10.965 ;
      RECT 22.225 10.795 22.395 10.965 ;
      RECT 21.765 10.795 21.935 10.965 ;
      RECT 21.305 10.795 21.475 10.965 ;
      RECT 20.845 10.795 21.015 10.965 ;
      RECT 20.385 10.795 20.555 10.965 ;
      RECT 19.925 10.795 20.095 10.965 ;
      RECT 19.465 10.795 19.635 10.965 ;
      RECT 19.005 10.795 19.175 10.965 ;
      RECT 18.545 10.795 18.715 10.965 ;
      RECT 18.085 10.795 18.255 10.965 ;
      RECT 17.625 10.795 17.795 10.965 ;
      RECT 17.165 10.795 17.335 10.965 ;
      RECT 16.705 10.795 16.875 10.965 ;
      RECT 16.245 10.795 16.415 10.965 ;
      RECT 15.785 10.795 15.955 10.965 ;
      RECT 15.325 10.795 15.495 10.965 ;
      RECT 14.865 10.795 15.035 10.965 ;
      RECT 14.405 10.795 14.575 10.965 ;
      RECT 13.945 10.795 14.115 10.965 ;
      RECT 13.485 10.795 13.655 10.965 ;
      RECT 13.025 10.795 13.195 10.965 ;
      RECT 12.565 10.795 12.735 10.965 ;
      RECT 12.105 10.795 12.275 10.965 ;
      RECT 11.645 10.795 11.815 10.965 ;
      RECT 11.185 10.795 11.355 10.965 ;
      RECT 10.725 10.795 10.895 10.965 ;
      RECT 10.265 10.795 10.435 10.965 ;
      RECT 9.805 10.795 9.975 10.965 ;
      RECT 9.345 10.795 9.515 10.965 ;
      RECT 8.885 10.795 9.055 10.965 ;
      RECT 8.425 10.795 8.595 10.965 ;
      RECT 7.965 10.795 8.135 10.965 ;
      RECT 7.505 10.795 7.675 10.965 ;
      RECT 7.045 10.795 7.215 10.965 ;
      RECT 6.585 10.795 6.755 10.965 ;
      RECT 6.125 10.795 6.295 10.965 ;
      RECT 5.665 10.795 5.835 10.965 ;
      RECT 5.205 10.795 5.375 10.965 ;
      RECT 4.745 10.795 4.915 10.965 ;
      RECT 4.285 10.795 4.455 10.965 ;
      RECT 3.825 10.795 3.995 10.965 ;
      RECT 3.365 10.795 3.535 10.965 ;
      RECT 2.905 10.795 3.075 10.965 ;
      RECT 2.445 10.795 2.615 10.965 ;
      RECT 1.985 10.795 2.155 10.965 ;
      RECT 1.525 10.795 1.695 10.965 ;
      RECT 1.065 10.795 1.235 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 95.365 8.075 95.535 8.245 ;
      RECT 94.905 8.075 95.075 8.245 ;
      RECT 28.205 8.075 28.375 8.245 ;
      RECT 27.745 8.075 27.915 8.245 ;
      RECT 95.365 5.355 95.535 5.525 ;
      RECT 94.905 5.355 95.075 5.525 ;
      RECT 28.205 5.355 28.375 5.525 ;
      RECT 27.745 5.355 27.915 5.525 ;
      RECT 95.365 2.635 95.535 2.805 ;
      RECT 94.905 2.635 95.075 2.805 ;
      RECT 28.205 2.635 28.375 2.805 ;
      RECT 27.745 2.635 27.915 2.805 ;
      RECT 95.365 -0.085 95.535 0.085 ;
      RECT 94.905 -0.085 95.075 0.085 ;
      RECT 94.445 -0.085 94.615 0.085 ;
      RECT 93.985 -0.085 94.155 0.085 ;
      RECT 93.525 -0.085 93.695 0.085 ;
      RECT 93.065 -0.085 93.235 0.085 ;
      RECT 92.605 -0.085 92.775 0.085 ;
      RECT 92.145 -0.085 92.315 0.085 ;
      RECT 91.685 -0.085 91.855 0.085 ;
      RECT 91.225 -0.085 91.395 0.085 ;
      RECT 90.765 -0.085 90.935 0.085 ;
      RECT 90.305 -0.085 90.475 0.085 ;
      RECT 89.845 -0.085 90.015 0.085 ;
      RECT 89.385 -0.085 89.555 0.085 ;
      RECT 88.925 -0.085 89.095 0.085 ;
      RECT 88.465 -0.085 88.635 0.085 ;
      RECT 88.005 -0.085 88.175 0.085 ;
      RECT 87.545 -0.085 87.715 0.085 ;
      RECT 87.085 -0.085 87.255 0.085 ;
      RECT 86.625 -0.085 86.795 0.085 ;
      RECT 86.165 -0.085 86.335 0.085 ;
      RECT 85.705 -0.085 85.875 0.085 ;
      RECT 85.245 -0.085 85.415 0.085 ;
      RECT 84.785 -0.085 84.955 0.085 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
    LAYER via ;
      RECT 83.645 97.845 83.795 97.995 ;
      RECT 54.205 97.845 54.355 97.995 ;
      RECT 10.045 97.845 10.195 97.995 ;
      RECT 115.845 12.505 115.995 12.655 ;
      RECT 14.185 12.505 14.335 12.655 ;
      RECT 83.645 10.805 83.795 10.955 ;
      RECT 54.205 10.805 54.355 10.955 ;
      RECT 10.045 10.805 10.195 10.955 ;
      RECT 77.665 1.625 77.815 1.775 ;
      RECT 58.805 1.625 58.955 1.775 ;
      RECT 52.825 1.625 52.975 1.775 ;
      RECT 83.645 -0.075 83.795 0.075 ;
      RECT 54.205 -0.075 54.355 0.075 ;
    LAYER via2 ;
      RECT 83.62 97.82 83.82 98.02 ;
      RECT 54.18 97.82 54.38 98.02 ;
      RECT 10.02 97.82 10.22 98.02 ;
      RECT 1.28 89.66 1.48 89.86 ;
      RECT 121.8 74.02 122 74.22 ;
      RECT 1.74 72.66 1.94 72.86 ;
      RECT 121.8 61.1 122 61.3 ;
      RECT 121.8 56.34 122 56.54 ;
      RECT 1.28 54.3 1.48 54.5 ;
      RECT 1.28 51.58 1.48 51.78 ;
      RECT 1.74 48.86 1.94 49.06 ;
      RECT 1.28 44.78 1.48 44.98 ;
      RECT 121.8 42.74 122 42.94 ;
      RECT 121.8 38.66 122 38.86 ;
      RECT 1.74 37.3 1.94 37.5 ;
      RECT 1.28 34.58 1.48 34.78 ;
      RECT 121.8 29.14 122 29.34 ;
      RECT 121.34 27.78 121.54 27.98 ;
      RECT 1.28 20.3 1.48 20.5 ;
      RECT 10.02 10.78 10.22 10.98 ;
      RECT 83.62 -0.1 83.82 0.1 ;
      RECT 54.18 -0.1 54.38 0.1 ;
    LAYER via3 ;
      RECT 83.62 97.82 83.82 98.02 ;
      RECT 54.18 97.82 54.38 98.02 ;
      RECT 10.02 97.82 10.22 98.02 ;
      RECT 121.34 81.5 121.54 81.7 ;
      RECT 10.02 10.78 10.22 10.98 ;
      RECT 83.62 -0.1 83.82 0.1 ;
      RECT 54.18 -0.1 54.38 0.1 ;
    LAYER OVERLAP ;
      POLYGON 27.6 0 27.6 10.88 0 10.88 0 97.92 123.28 97.92 123.28 10.88 95.68 10.88 95.68 0 ;
  END
END sb_1__2_

END LIBRARY
