//
//
//
//
//
//
module mux_tree_tapbuf_size3_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__39 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size3_0 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size3 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__37 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__36 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size5 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size5_0 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__35 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__34 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size6 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size6_0 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__33 ( .A ( mem_out[1] ) , 
    .X ( net_aps_33 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_65 ( .A ( net_aps_33 ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__32 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__31 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__30 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__29 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__28 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__27 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__26 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_9 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__25 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__24 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_10 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__23 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__22 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_7 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_6 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_5 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_4 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_3 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_2 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_1 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_0 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_9 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_43 ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_10 ( in , sram , sram_inv , out , VDD , VSS , 
    p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_41 ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_8 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module sb_0__0_ ( prog_clk , chany_top_in , top_left_grid_pin_1_ , 
    chanx_right_in , right_top_grid_pin_42_ , right_top_grid_pin_43_ , 
    right_top_grid_pin_44_ , right_top_grid_pin_45_ , right_top_grid_pin_46_ , 
    right_top_grid_pin_47_ , right_top_grid_pin_48_ , right_top_grid_pin_49_ , 
    right_bottom_grid_pin_1_ , ccff_head , chany_top_out , chanx_right_out , 
    ccff_tail , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_top_in ;
input  [0:0] top_left_grid_pin_1_ ;
input  [0:19] chanx_right_in ;
input  [0:0] right_top_grid_pin_42_ ;
input  [0:0] right_top_grid_pin_43_ ;
input  [0:0] right_top_grid_pin_44_ ;
input  [0:0] right_top_grid_pin_45_ ;
input  [0:0] right_top_grid_pin_46_ ;
input  [0:0] right_top_grid_pin_47_ ;
input  [0:0] right_top_grid_pin_48_ ;
input  [0:0] right_top_grid_pin_49_ ;
input  [0:0] right_bottom_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chany_top_out ;
output [0:19] chanx_right_out ;
output [0:0] ccff_tail ;
input  VDD ;
input  VSS ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_10_sram ;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_11_sram ;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_5_sram ;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_6_sram ;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_7_sram ;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_8_sram ;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_9_sram ;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size5_0_sram ;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_1_sram ;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;
supply1 VDD ;
supply0 VSS ;
//

mux_tree_tapbuf_size2_8 mux_top_track_0 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[1] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chany_top_out[0] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_10 mux_top_track_4 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[3] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) ,
    .out ( { ropt_net_116 } ) ,
    .VDD ( VDD ) , .VSS ( VSS ) , .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2 mux_top_track_8 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[5] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) , 
    .out ( chany_top_out[4] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_9 mux_top_track_24 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) ,
    .out ( { ropt_net_119 } ) ,
    .VDD ( VDD ) , .VSS ( VSS ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_0 mux_right_track_10 (
    .in ( { chany_top_in[4] , right_top_grid_pin_43_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chanx_right_out[5] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size2_1 mux_right_track_12 (
    .in ( { chany_top_in[5] , right_top_grid_pin_44_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_5_sram_inv ) , 
    .out ( chanx_right_out[6] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_2 mux_right_track_14 (
    .in ( { chany_top_in[6] , right_top_grid_pin_45_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_6_sram_inv ) , 
    .out ( chanx_right_out[7] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_3 mux_right_track_16 (
    .in ( { chany_top_in[7] , right_top_grid_pin_46_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_7_sram_inv ) , 
    .out ( chanx_right_out[8] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_4 mux_right_track_18 (
    .in ( { chany_top_in[8] , right_top_grid_pin_47_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_8_sram_inv ) , 
    .out ( chanx_right_out[9] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_5 mux_right_track_20 (
    .in ( { chany_top_in[9] , right_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_9_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_9_sram_inv ) , 
    .out ( chanx_right_out[10] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_6 mux_right_track_22 (
    .in ( { chany_top_in[10] , right_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_10_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_10_sram_inv ) , 
    .out ( chanx_right_out[11] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_7 mux_right_track_26 (
    .in ( { chany_top_in[12] , right_top_grid_pin_43_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_11_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_11_sram_inv ) , 
    .out ( chanx_right_out[13] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_mem_8 mem_top_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_10 mem_top_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem mem_top_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_9 mem_top_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_0 mem_right_track_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_1 mem_right_track_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_5_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_2 mem_right_track_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_6_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_3 mem_right_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_7_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_4 mem_right_track_18 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_8_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_5 mem_right_track_20 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_9_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_9_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_6 mem_right_track_22 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_10_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_10_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_7 mem_right_track_26 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) ,
    .ccff_tail ( { ropt_net_117 } ) ,
    .mem_out ( mux_tree_tapbuf_size2_11_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_11_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size6_0 mux_right_track_0 (
    .in ( { chany_top_in[19] , right_top_grid_pin_42_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_46_[0] , 
        right_top_grid_pin_48_[0] , right_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chanx_right_out[0] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size6 mux_right_track_4 (
    .in ( { chany_top_in[1] , right_top_grid_pin_42_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_46_[0] , 
        right_top_grid_pin_48_[0] , right_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chanx_right_out[2] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size6_mem_0 mem_right_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size6_mem mem_right_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size5_0 mux_right_track_2 (
    .in ( { chany_top_in[0] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_45_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size5_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_0_sram_inv ) , 
    .out ( chanx_right_out[1] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size5 mux_right_track_6 (
    .in ( { chany_top_in[2] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_45_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size5_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_1_sram_inv ) , 
    .out ( chanx_right_out[3] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size5_mem_0 mem_right_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_0_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size5_mem mem_right_track_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_1_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size3 mux_right_track_8 (
    .in ( { chany_top_in[3] , right_top_grid_pin_42_[0] , 
        right_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chanx_right_out[4] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size3_0 mux_right_track_24 (
    .in ( { chany_top_in[11] , right_top_grid_pin_42_[0] , 
        right_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) , 
    .out ( chanx_right_out[12] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size3_mem mem_right_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size3_mem_0 mem_right_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
sky130_fd_sc_hd__conb_1 optlc_105 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_112 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__conb_1 optlc_107 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_113 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__conb_1 optlc_109 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_114 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__conb_1 optlc_111 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_115 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_728 ( .A ( ropt_net_116 ) , 
    .X ( ropt_net_141 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_6__5 ( .A ( chany_top_in[18] ) , 
    .X ( ropt_net_134 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_757 ( .A ( ropt_net_139 ) , 
    .X ( chany_top_out[5] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_758 ( .A ( ropt_net_140 ) , 
    .X ( chany_top_out[16] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_759 ( .A ( ropt_net_141 ) , 
    .X ( chany_top_out[2] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_761 ( .A ( ropt_net_142 ) , 
    .X ( chanx_right_out[15] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_729 ( .A ( ropt_net_117 ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_730 ( .A ( chanx_right_in[0] ) , 
    .X ( chany_top_out[19] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_731 ( .A ( ropt_net_119 ) , 
    .X ( chany_top_out[12] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_732 ( .A ( ropt_net_120 ) , 
    .X ( chany_top_out[15] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_765 ( .A ( ropt_net_143 ) , 
    .X ( chany_top_out[14] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_767 ( .A ( ropt_net_144 ) , 
    .X ( chany_top_out[1] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_768 ( .A ( ropt_net_145 ) , 
    .X ( chany_top_out[3] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_733 ( .A ( chanx_right_in[12] ) , 
    .X ( chany_top_out[11] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_771 ( .A ( ropt_net_146 ) , 
    .X ( chanx_right_out[16] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_772 ( .A ( ropt_net_147 ) , 
    .X ( chanx_right_out[17] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_734 ( .A ( chanx_right_in[2] ) , 
    .X ( ropt_net_144 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_735 ( .A ( chanx_right_in[14] ) , 
    .X ( chany_top_out[13] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_57 ( .A ( chanx_right_in[11] ) , 
    .X ( BUF_net_57 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_736 ( .A ( chanx_right_in[18] ) , 
    .X ( chany_top_out[17] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_62 ( .A ( chanx_right_in[17] ) , 
    .X ( BUF_net_62 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_64 ( .A ( chanx_right_in[19] ) , 
    .X ( BUF_net_64 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_737 ( .A ( ropt_net_125 ) , 
    .X ( ropt_net_139 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_73 ( .A ( chanx_right_in[6] ) , 
    .X ( ropt_net_125 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_739 ( .A ( chanx_right_in[4] ) , 
    .X ( ropt_net_145 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_742 ( .A ( chanx_right_in[8] ) , 
    .X ( chany_top_out[7] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_743 ( .A ( chany_top_in[15] ) , 
    .X ( ropt_net_146 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_744 ( .A ( chanx_right_in[10] ) , 
    .X ( chany_top_out[9] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_78 ( .A ( BUF_net_57 ) , 
    .X ( chany_top_out[10] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_745 ( .A ( chany_top_in[16] ) , 
    .X ( ropt_net_147 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_82 ( .A ( chanx_right_in[16] ) , 
    .X ( ropt_net_120 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_83 ( .A ( BUF_net_62 ) , 
    .X ( ropt_net_140 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_85 ( .A ( BUF_net_64 ) , 
    .X ( chany_top_out[18] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_97 ( .A ( chany_top_in[14] ) , 
    .X ( ropt_net_135 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_98 ( .A ( chanx_right_in[7] ) , 
    .X ( chany_top_out[6] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_746 ( .A ( chanx_right_in[9] ) , 
    .X ( chany_top_out[8] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_747 ( .A ( chany_top_in[17] ) , 
    .X ( chanx_right_out[18] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_101 ( .A ( chanx_right_in[15] ) , 
    .X ( ropt_net_143 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_748 ( .A ( chany_top_in[13] ) , 
    .X ( chanx_right_out[14] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_750 ( .A ( ropt_net_134 ) , 
    .X ( chanx_right_out[19] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_752 ( .A ( ropt_net_135 ) , 
    .X ( ropt_net_142 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x883200y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x920000y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x956800y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x993600y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1030400y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1067200y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x883200y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x920000y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x956800y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x993600y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1030400y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1067200y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x883200y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x920000y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x956800y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x993600y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1030400y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1067200y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x883200y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x920000y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x956800y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x993600y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1030400y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1067200y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x883200y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x920000y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x956800y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x993600y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1030400y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1067200y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x883200y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x920000y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x956800y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x993600y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1030400y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1067200y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x883200y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x920000y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x956800y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x993600y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1030400y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1067200y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x883200y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x920000y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x956800y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x993600y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1030400y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1048800y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x883200y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x920000y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x956800y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x993600y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1030400y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1048800y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x883200y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x920000y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x956800y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x993600y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1030400y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1067200y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x883200y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x920000y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x956800y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x993600y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1030400y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1067200y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x883200y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x920000y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x956800y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x993600y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1030400y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1067200y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x883200y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x920000y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x956800y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1002800y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1039600y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1076400y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1113200y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x662400y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x671600y353600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x713000y353600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x805000y353600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x897000y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x915400y353600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x947600y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x984400y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1021200y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x588800y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x598000y380800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x690000y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x726800y380800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x846400y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x883200y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x929200y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x966000y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1002800y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1021200y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x662400y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x754400y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x791200y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x841800y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x864800y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x901600y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x938400y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x975200y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1012000y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x1021200y408000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x478400y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x496800y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x506000y435200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x588800y435200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x680800y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x717600y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x754400y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x763600y435200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x805000y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x841800y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x860200y435200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x943000y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x979800y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x1016600y435200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1048800y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x368000y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x386400y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x395600y462400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x529000y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x538200y462400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x708400y462400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x887800y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x906200y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1002800y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1039600y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1076400y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1113200y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x331200y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x349600y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x358800y489600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x400200y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x437000y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x473800y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x510600y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x547400y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x584200y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x621000y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x657800y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x694600y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x818800y489600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x910800y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x947600y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x984400y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1021200y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1058000y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x331200y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x349600y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x358800y516800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x450800y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x529000y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x565800y516800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x782000y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x841800y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x878600y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x915400y516800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1048800y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x409400y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x446200y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x464600y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x473800y544000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x506000y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x542800y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x579600y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x846400y544000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x933800y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x970600y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1007400y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x1025800y544000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x478400y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x496800y571200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x860200y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x897000y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1085600y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x331200y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x427800y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x460000y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x496800y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x533600y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x630200y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x726800y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x763600y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x800400y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x809600y598400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x943000y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x979800y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1016600y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1053400y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1090200y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x1127000y598400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x331200y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x391000y625600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x432400y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x469200y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x487600y625600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x529000y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x565800y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x602600y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x676200y625600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x722200y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x731400y625600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x823400y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x883200y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x901600y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x910800y625600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x952200y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1012000y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x220800y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x262200y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x299000y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x335800y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x372600y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x409400y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x446200y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x483000y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x501400y652800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x593400y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x630200y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x667000y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x703800y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x740600y652800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x846400y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x368000y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x464600y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x501400y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x552000y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x561200y680000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x607200y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x625600y680000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x754400y680000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x795800y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x855600y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x874000y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x883200y680000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x924600y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x961400y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x970600y680000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1002800y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1039600y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1104000y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1122400y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x368000y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x386400y707200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x556600y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x593400y707200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x639400y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x657800y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x708400y707200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x754400y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x763600y707200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x846400y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x897000y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x915400y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x924600y707200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x970600y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1007400y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1044200y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1081000y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x1117800y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x1127000y707200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x331200y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x386400y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x423200y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x460000y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x478400y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x575000y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x611800y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x630200y734400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x676200y734400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x713000y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x818800y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x855600y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x892400y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x929200y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x966000y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1002800y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1039600y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x1076400y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x1113200y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x294400y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x312800y761600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x478400y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x510600y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x625600y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x731400y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x368000y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x386400y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x437000y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x473800y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x598000y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x634800y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x671600y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x708400y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x745200y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x782000y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x818800y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x837200y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x368000y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x386400y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x395600y816000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x441600y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x450800y816000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x487600y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x506000y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x547400y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x584200y816000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x630200y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x667000y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x703800y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x740600y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x759000y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x768200y816000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x814200y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x832600y816000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y816000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x331200y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x427800y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x464600y843200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x510600y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x547400y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x584200y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x621000y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x717600y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x754400y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x805000y843200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y843200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x331200y870400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x363400y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x400200y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x418600y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x460000y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x496800y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x547400y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x584200y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x602600y870400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x644000y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x680800y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x759000y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x768200y870400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x814200y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x832600y870400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y870400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x184000y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x234600y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x271400y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x308200y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x345000y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x381800y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x437000y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x446200y897600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x492200y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x529000y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x565800y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x602600y897600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x694600y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x754400y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x805000y897600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y897600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x73600y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x92000y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x331200y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x349600y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x358800y924800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x584200y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x621000y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x657800y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x736000y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x754400y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x763600y924800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y924800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y952000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x36800y952000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x133400y952000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x170200y952000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x207000y952000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x308200y952000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x317400y952000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x354200y952000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x372600y952000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x607200y952000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x800400y952000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x837200y952000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y979200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x36800y979200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x55200y979200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x151800y979200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x188600y979200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x621000y979200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x639400y979200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x818800y979200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x837200y979200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x552000y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x662400y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y1006400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
endmodule


