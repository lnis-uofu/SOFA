VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_2__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 84.64 BY 97.92 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 2.23 80.24 2.37 81.6 ;
    END
  END prog_clk[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.51 96.56 56.65 97.92 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.05 96.56 33.19 97.92 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.89 96.56 57.19 97.92 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.13 96.56 32.27 97.92 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.93 96.56 23.07 97.92 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.15 96.56 49.29 97.92 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.87 96.56 64.01 97.92 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 96.56 57.57 97.92 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.03 96.56 62.17 97.92 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.85 96.56 46.15 97.92 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.61 96.56 48.91 97.92 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 96.56 48.37 97.92 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 96.56 52.97 97.92 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.79 96.56 64.93 97.92 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.11 96.56 61.25 97.92 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.27 96.56 59.41 97.92 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 96.56 50.21 97.92 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.95 96.56 63.09 97.92 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.35 96.56 58.49 97.92 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.19 96.56 60.33 97.92 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.69 96.56 24.99 97.92 ;
    END
  END top_left_grid_pin_42_[0]
  PIN top_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.65 96.56 36.95 97.92 ;
    END
  END top_left_grid_pin_43_[0]
  PIN top_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.85 96.56 23.15 97.92 ;
    END
  END top_left_grid_pin_44_[0]
  PIN top_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.55 96.56 21.69 97.92 ;
    END
  END top_left_grid_pin_45_[0]
  PIN top_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 34.81 96.56 35.11 97.92 ;
    END
  END top_left_grid_pin_46_[0]
  PIN top_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.67 80.24 8.81 81.6 ;
    END
  END top_left_grid_pin_47_[0]
  PIN top_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.63 96.56 20.77 97.92 ;
    END
  END top_left_grid_pin_48_[0]
  PIN top_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.27 80.24 13.41 81.6 ;
    END
  END top_left_grid_pin_49_[0]
  PIN top_right_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.85 96.56 23.99 97.92 ;
    END
  END top_right_grid_pin_1_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.33 0 41.47 1.36 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.15 0 49.29 1.36 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 0 51.13 1.36 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.25 0 42.39 1.36 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.01 0 22.15 1.36 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.57 0 38.71 1.36 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.49 0 39.63 1.36 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.95 0 63.09 1.36 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.57 0 61.71 1.36 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.79 0 64.93 1.36 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.73 0 36.87 1.36 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 0 57.57 1.36 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.41 0 40.55 1.36 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.21 0 31.35 1.36 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 0 52.05 1.36 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.73 0 59.87 1.36 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.35 0 58.49 1.36 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.65 0 60.79 1.36 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.87 0 64.01 1.36 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.51 0 56.65 1.36 ;
    END
  END chany_bottom_in[19]
  PIN bottom_right_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.69 0 25.83 1.36 ;
    END
  END bottom_right_grid_pin_1_[0]
  PIN bottom_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.61 16.32 3.75 17.68 ;
    END
  END bottom_left_grid_pin_42_[0]
  PIN bottom_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.85 0 23.15 1.36 ;
    END
  END bottom_left_grid_pin_43_[0]
  PIN bottom_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.29 1.38 22.59 ;
    END
  END bottom_left_grid_pin_44_[0]
  PIN bottom_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.53 16.32 4.67 17.68 ;
    END
  END bottom_left_grid_pin_45_[0]
  PIN bottom_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.69 16.32 2.83 17.68 ;
    END
  END bottom_left_grid_pin_46_[0]
  PIN bottom_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 20.93 1.38 21.23 ;
    END
  END bottom_left_grid_pin_47_[0]
  PIN bottom_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.83 16.32 6.97 17.68 ;
    END
  END bottom_left_grid_pin_48_[0]
  PIN bottom_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 19.57 1.38 19.87 ;
    END
  END bottom_left_grid_pin_49_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 51.53 1.38 51.83 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 23.65 1.38 23.95 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.69 1.38 42.99 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 34.53 1.38 34.83 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 35.89 1.38 36.19 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 30.45 1.38 30.75 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 4.45 16.32 4.75 17.68 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 65.81 1.38 66.11 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.89 1.38 70.19 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 61.05 1.38 61.35 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 41.33 1.38 41.63 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 58.33 1.38 58.63 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 64.45 1.38 64.75 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 55.61 1.38 55.91 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 77.37 1.38 77.67 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.89 1.38 53.19 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 73.29 1.38 73.59 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 74.65 1.38 74.95 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 76.01 1.38 76.31 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.09 1.38 29.39 ;
    END
  END chanx_left_in[19]
  PIN left_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 18.4 6.65 19.78 6.95 ;
    END
  END left_bottom_grid_pin_34_[0]
  PIN left_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 18.4 5.29 19.78 5.59 ;
    END
  END left_bottom_grid_pin_35_[0]
  PIN left_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.67 16.32 8.81 17.68 ;
    END
  END left_bottom_grid_pin_36_[0]
  PIN left_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.45 16.32 5.59 17.68 ;
    END
  END left_bottom_grid_pin_37_[0]
  PIN left_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.63 0 20.77 1.36 ;
    END
  END left_bottom_grid_pin_38_[0]
  PIN left_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.59 16.32 9.73 17.68 ;
    END
  END left_bottom_grid_pin_39_[0]
  PIN left_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.69 0 24.99 1.36 ;
    END
  END left_bottom_grid_pin_40_[0]
  PIN left_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.75 16.32 7.89 17.68 ;
    END
  END left_bottom_grid_pin_41_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.03 96.56 39.17 97.92 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.87 96.56 41.01 97.92 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.97 96.56 34.11 97.92 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 96.56 46.53 97.92 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 96.56 52.05 97.92 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.17 96.56 43.31 97.92 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.69 96.56 25.83 97.92 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.35 96.56 35.49 97.92 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 96.56 47.45 97.92 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.65 96.56 37.79 97.92 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 96.56 51.13 97.92 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.73 96.56 36.87 97.92 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.75 96.56 53.89 97.92 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.37 96.56 29.51 97.92 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.95 96.56 40.09 97.92 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.61 96.56 26.75 97.92 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 96.56 45.61 97.92 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.77 96.56 24.91 97.92 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.45 96.56 28.59 97.92 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.25 96.56 42.39 97.92 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.53 96.56 27.67 97.92 ;
    END
  END chany_top_out[19]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.13 0 32.27 1.36 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.05 0 79.19 1.36 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.13 0 78.27 1.36 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.65 0 37.79 1.36 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.37 0 29.51 1.36 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.93 0 23.07 1.36 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.85 0 23.99 1.36 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 0 46.53 1.36 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.17 0 43.31 1.36 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 0 50.21 1.36 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.43 0 34.57 1.36 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.45 0 28.59 1.36 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.61 0 26.75 1.36 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.77 0 24.91 1.36 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.29 0 30.43 1.36 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 0 47.45 1.36 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.53 0 27.67 1.36 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.05 0 33.19 1.36 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 0 48.37 1.36 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 0 45.61 1.36 ;
    END
  END chany_bottom_out[19]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 45.41 1.38 45.71 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.97 1.38 57.27 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 71.25 1.38 71.55 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 27.73 1.38 28.03 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.81 1.38 49.11 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 46.77 1.38 47.07 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 38.61 1.38 38.91 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 54.25 1.38 54.55 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.05 1.38 44.35 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.17 1.38 33.47 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 67.17 1.38 67.47 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.17 1.38 50.47 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 26.37 1.38 26.67 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 6.29 16.32 6.59 17.68 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.01 1.38 25.31 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.97 1.38 40.27 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.69 1.38 59.99 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.25 1.38 37.55 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.81 1.38 32.11 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 68.53 1.38 68.83 ;
    END
  END chanx_left_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 63.09 1.38 63.39 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 18.4 2.48 18.88 2.96 ;
        RECT 84.16 2.48 84.64 2.96 ;
        RECT 18.4 7.92 18.88 8.4 ;
        RECT 84.16 7.92 84.64 8.4 ;
        RECT 18.4 13.36 18.88 13.84 ;
        RECT 84.16 13.36 84.64 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 84.16 18.8 84.64 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 84.16 24.24 84.64 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 84.16 29.68 84.64 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 84.16 35.12 84.64 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 84.16 40.56 84.64 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 84.16 46 84.64 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 84.16 51.44 84.64 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 84.16 56.88 84.64 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 84.16 62.32 84.64 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 84.16 67.76 84.64 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 84.16 73.2 84.64 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 84.16 78.64 84.64 79.12 ;
        RECT 18.4 84.08 18.88 84.56 ;
        RECT 84.16 84.08 84.64 84.56 ;
        RECT 18.4 89.52 18.88 90 ;
        RECT 84.16 89.52 84.64 90 ;
        RECT 18.4 94.96 18.88 95.44 ;
        RECT 84.16 94.96 84.64 95.44 ;
      LAYER met4 ;
        RECT 29.14 0 29.74 0.6 ;
        RECT 58.58 0 59.18 0.6 ;
        RECT 29.14 97.32 29.74 97.92 ;
        RECT 58.58 97.32 59.18 97.92 ;
      LAYER met5 ;
        RECT 0 26.96 3.2 30.16 ;
        RECT 81.44 26.96 84.64 30.16 ;
        RECT 0 67.76 3.2 70.96 ;
        RECT 81.44 67.76 84.64 70.96 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 18.4 0 84.64 0.24 ;
        RECT 18.4 5.2 18.88 5.68 ;
        RECT 84.16 5.2 84.64 5.68 ;
        RECT 18.4 10.64 18.88 11.12 ;
        RECT 84.16 10.64 84.64 11.12 ;
        RECT 0 16.08 84.64 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 84.16 21.52 84.64 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 84.16 26.96 84.64 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 84.16 32.4 84.64 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 84.16 37.84 84.64 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 84.16 43.28 84.64 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 84.16 48.72 84.64 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 84.16 54.16 84.64 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 84.16 59.6 84.64 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 84.16 65.04 84.64 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 84.16 70.48 84.64 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 84.16 75.92 84.64 76.4 ;
        RECT 0 81.36 84.64 81.84 ;
        RECT 18.4 86.8 18.88 87.28 ;
        RECT 84.16 86.8 84.64 87.28 ;
        RECT 18.4 92.24 18.88 92.72 ;
        RECT 84.16 92.24 84.64 92.72 ;
        RECT 18.4 97.68 84.64 97.92 ;
      LAYER met4 ;
        RECT 43.86 0 44.46 0.6 ;
        RECT 73.3 0 73.9 0.6 ;
        RECT 43.86 97.32 44.46 97.92 ;
        RECT 73.3 97.32 73.9 97.92 ;
      LAYER met5 ;
        RECT 0 47.36 3.2 50.56 ;
        RECT 81.44 47.36 84.64 50.56 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 18.4 97.835 84.64 98.005 ;
      RECT 84.18 95.115 84.64 95.285 ;
      RECT 18.4 95.115 22.08 95.285 ;
      RECT 84.18 92.395 84.64 92.565 ;
      RECT 18.4 92.395 20.24 92.565 ;
      RECT 83.72 89.675 84.64 89.845 ;
      RECT 18.4 89.675 22.08 89.845 ;
      RECT 83.72 86.955 84.64 87.125 ;
      RECT 18.4 86.955 22.08 87.125 ;
      RECT 80.96 84.235 84.64 84.405 ;
      RECT 18.4 84.235 20.24 84.405 ;
      RECT 80.96 81.515 84.64 81.685 ;
      RECT 0 81.515 20.24 81.685 ;
      RECT 80.96 78.795 84.64 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 80.96 76.075 84.64 76.245 ;
      RECT 0 76.075 1.84 76.245 ;
      RECT 83.72 73.355 84.64 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 80.96 70.635 84.64 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 80.96 67.915 84.64 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 83.72 65.195 84.64 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 83.72 62.475 84.64 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 83.72 59.755 84.64 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 83.72 57.035 84.64 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 83.72 54.315 84.64 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 83.72 51.595 84.64 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 83.72 48.875 84.64 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 83.72 46.155 84.64 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 83.72 43.435 84.64 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 83.72 40.715 84.64 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 83.72 37.995 84.64 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 83.72 35.275 84.64 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 83.72 32.555 84.64 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 83.72 29.835 84.64 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 83.72 27.115 84.64 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 83.72 24.395 84.64 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 83.72 21.675 84.64 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 83.72 18.955 84.64 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 83.72 16.235 84.64 16.405 ;
      RECT 0 16.235 22.08 16.405 ;
      RECT 83.72 13.515 84.64 13.685 ;
      RECT 18.4 13.515 20.24 13.685 ;
      RECT 83.72 10.795 84.64 10.965 ;
      RECT 18.4 10.795 22.08 10.965 ;
      RECT 83.72 8.075 84.64 8.245 ;
      RECT 18.4 8.075 22.08 8.245 ;
      RECT 84.18 5.355 84.64 5.525 ;
      RECT 18.4 5.355 20.24 5.525 ;
      RECT 84.18 2.635 84.64 2.805 ;
      RECT 18.4 2.635 22.08 2.805 ;
      RECT 18.4 -0.085 84.64 0.085 ;
    LAYER met2 ;
      RECT 73.46 97.735 73.74 98.105 ;
      RECT 44.02 97.735 44.3 98.105 ;
      RECT 33.45 96.06 33.71 96.38 ;
      RECT 41.73 1.54 41.99 1.86 ;
      RECT 28.85 1.54 29.11 1.86 ;
      RECT 73.46 -0.185 73.74 0.185 ;
      RECT 44.02 -0.185 44.3 0.185 ;
      POLYGON 84.36 97.64 84.36 0.28 79.47 0.28 79.47 1.64 78.77 1.64 78.77 0.28 78.55 0.28 78.55 1.64 77.85 1.64 77.85 0.28 65.21 0.28 65.21 1.64 64.51 1.64 64.51 0.28 64.29 0.28 64.29 1.64 63.59 1.64 63.59 0.28 63.37 0.28 63.37 1.64 62.67 1.64 62.67 0.28 61.99 0.28 61.99 1.64 61.29 1.64 61.29 0.28 61.07 0.28 61.07 1.64 60.37 1.64 60.37 0.28 60.15 0.28 60.15 1.64 59.45 1.64 59.45 0.28 58.77 0.28 58.77 1.64 58.07 1.64 58.07 0.28 57.85 0.28 57.85 1.64 57.15 1.64 57.15 0.28 56.93 0.28 56.93 1.64 56.23 1.64 56.23 0.28 52.33 0.28 52.33 1.64 51.63 1.64 51.63 0.28 51.41 0.28 51.41 1.64 50.71 1.64 50.71 0.28 50.49 0.28 50.49 1.64 49.79 1.64 49.79 0.28 49.57 0.28 49.57 1.64 48.87 1.64 48.87 0.28 48.65 0.28 48.65 1.64 47.95 1.64 47.95 0.28 47.73 0.28 47.73 1.64 47.03 1.64 47.03 0.28 46.81 0.28 46.81 1.64 46.11 1.64 46.11 0.28 45.89 0.28 45.89 1.64 45.19 1.64 45.19 0.28 43.59 0.28 43.59 1.64 42.89 1.64 42.89 0.28 42.67 0.28 42.67 1.64 41.97 1.64 41.97 0.28 41.75 0.28 41.75 1.64 41.05 1.64 41.05 0.28 40.83 0.28 40.83 1.64 40.13 1.64 40.13 0.28 39.91 0.28 39.91 1.64 39.21 1.64 39.21 0.28 38.99 0.28 38.99 1.64 38.29 1.64 38.29 0.28 38.07 0.28 38.07 1.64 37.37 1.64 37.37 0.28 37.15 0.28 37.15 1.64 36.45 1.64 36.45 0.28 34.85 0.28 34.85 1.64 34.15 1.64 34.15 0.28 33.47 0.28 33.47 1.64 32.77 1.64 32.77 0.28 32.55 0.28 32.55 1.64 31.85 1.64 31.85 0.28 31.63 0.28 31.63 1.64 30.93 1.64 30.93 0.28 30.71 0.28 30.71 1.64 30.01 1.64 30.01 0.28 29.79 0.28 29.79 1.64 29.09 1.64 29.09 0.28 28.87 0.28 28.87 1.64 28.17 1.64 28.17 0.28 27.95 0.28 27.95 1.64 27.25 1.64 27.25 0.28 27.03 0.28 27.03 1.64 26.33 1.64 26.33 0.28 26.11 0.28 26.11 1.64 25.41 1.64 25.41 0.28 25.19 0.28 25.19 1.64 24.49 1.64 24.49 0.28 24.27 0.28 24.27 1.64 23.57 1.64 23.57 0.28 23.35 0.28 23.35 1.64 22.65 1.64 22.65 0.28 22.43 0.28 22.43 1.64 21.73 1.64 21.73 0.28 21.05 0.28 21.05 1.64 20.35 1.64 20.35 0.28 18.68 0.28 18.68 16.6 10.01 16.6 10.01 17.96 9.31 17.96 9.31 16.6 9.09 16.6 9.09 17.96 8.39 17.96 8.39 16.6 8.17 16.6 8.17 17.96 7.47 17.96 7.47 16.6 7.25 16.6 7.25 17.96 6.55 17.96 6.55 16.6 5.87 16.6 5.87 17.96 5.17 17.96 5.17 16.6 4.95 16.6 4.95 17.96 4.25 17.96 4.25 16.6 4.03 16.6 4.03 17.96 3.33 17.96 3.33 16.6 3.11 16.6 3.11 17.96 2.41 17.96 2.41 16.6 0.28 16.6 0.28 81.32 1.95 81.32 1.95 79.96 2.65 79.96 2.65 81.32 8.39 81.32 8.39 79.96 9.09 79.96 9.09 81.32 12.99 81.32 12.99 79.96 13.69 79.96 13.69 81.32 18.68 81.32 18.68 97.64 20.35 97.64 20.35 96.28 21.05 96.28 21.05 97.64 21.27 97.64 21.27 96.28 21.97 96.28 21.97 97.64 22.65 97.64 22.65 96.28 23.35 96.28 23.35 97.64 23.57 97.64 23.57 96.28 24.27 96.28 24.27 97.64 24.49 97.64 24.49 96.28 25.19 96.28 25.19 97.64 25.41 97.64 25.41 96.28 26.11 96.28 26.11 97.64 26.33 97.64 26.33 96.28 27.03 96.28 27.03 97.64 27.25 97.64 27.25 96.28 27.95 96.28 27.95 97.64 28.17 97.64 28.17 96.28 28.87 96.28 28.87 97.64 29.09 97.64 29.09 96.28 29.79 96.28 29.79 97.64 31.85 97.64 31.85 96.28 32.55 96.28 32.55 97.64 32.77 97.64 32.77 96.28 33.47 96.28 33.47 97.64 33.69 97.64 33.69 96.28 34.39 96.28 34.39 97.64 35.07 97.64 35.07 96.28 35.77 96.28 35.77 97.64 36.45 97.64 36.45 96.28 37.15 96.28 37.15 97.64 37.37 97.64 37.37 96.28 38.07 96.28 38.07 97.64 38.75 97.64 38.75 96.28 39.45 96.28 39.45 97.64 39.67 97.64 39.67 96.28 40.37 96.28 40.37 97.64 40.59 97.64 40.59 96.28 41.29 96.28 41.29 97.64 41.97 97.64 41.97 96.28 42.67 96.28 42.67 97.64 42.89 97.64 42.89 96.28 43.59 96.28 43.59 97.64 45.19 97.64 45.19 96.28 45.89 96.28 45.89 97.64 46.11 97.64 46.11 96.28 46.81 96.28 46.81 97.64 47.03 97.64 47.03 96.28 47.73 96.28 47.73 97.64 47.95 97.64 47.95 96.28 48.65 96.28 48.65 97.64 48.87 97.64 48.87 96.28 49.57 96.28 49.57 97.64 49.79 97.64 49.79 96.28 50.49 96.28 50.49 97.64 50.71 97.64 50.71 96.28 51.41 96.28 51.41 97.64 51.63 97.64 51.63 96.28 52.33 96.28 52.33 97.64 52.55 97.64 52.55 96.28 53.25 96.28 53.25 97.64 53.47 97.64 53.47 96.28 54.17 96.28 54.17 97.64 56.23 97.64 56.23 96.28 56.93 96.28 56.93 97.64 57.15 97.64 57.15 96.28 57.85 96.28 57.85 97.64 58.07 97.64 58.07 96.28 58.77 96.28 58.77 97.64 58.99 97.64 58.99 96.28 59.69 96.28 59.69 97.64 59.91 97.64 59.91 96.28 60.61 96.28 60.61 97.64 60.83 97.64 60.83 96.28 61.53 96.28 61.53 97.64 61.75 97.64 61.75 96.28 62.45 96.28 62.45 97.64 62.67 97.64 62.67 96.28 63.37 96.28 63.37 97.64 63.59 97.64 63.59 96.28 64.29 96.28 64.29 97.64 64.51 97.64 64.51 96.28 65.21 96.28 65.21 97.64 ;
    LAYER met4 ;
      POLYGON 84.24 97.52 84.24 0.4 74.3 0.4 74.3 1 72.9 1 72.9 0.4 59.58 0.4 59.58 1 58.18 1 58.18 0.4 44.86 0.4 44.86 1 43.46 1 43.46 0.4 30.14 0.4 30.14 1 28.74 1 28.74 0.4 25.39 0.4 25.39 1.76 24.29 1.76 24.29 0.4 23.55 0.4 23.55 1.76 22.45 1.76 22.45 0.4 18.8 0.4 18.8 16.72 6.99 16.72 6.99 18.08 5.89 18.08 5.89 16.72 5.15 16.72 5.15 18.08 4.05 18.08 4.05 16.72 0.4 16.72 0.4 81.2 18.8 81.2 18.8 97.52 22.45 97.52 22.45 96.16 23.55 96.16 23.55 97.52 24.29 97.52 24.29 96.16 25.39 96.16 25.39 97.52 28.74 97.52 28.74 96.92 30.14 96.92 30.14 97.52 34.41 97.52 34.41 96.16 35.51 96.16 35.51 97.52 36.25 97.52 36.25 96.16 37.35 96.16 37.35 97.52 43.46 97.52 43.46 96.92 44.86 96.92 44.86 97.52 45.45 97.52 45.45 96.16 46.55 96.16 46.55 97.52 48.21 97.52 48.21 96.16 49.31 96.16 49.31 97.52 56.49 97.52 56.49 96.16 57.59 96.16 57.59 97.52 58.18 97.52 58.18 96.92 59.58 96.92 59.58 97.52 72.9 97.52 72.9 96.92 74.3 96.92 74.3 97.52 ;
    LAYER met3 ;
      POLYGON 73.765 98.085 73.765 98.08 73.98 98.08 73.98 97.76 73.765 97.76 73.765 97.755 73.435 97.755 73.435 97.76 73.22 97.76 73.22 98.08 73.435 98.08 73.435 98.085 ;
      POLYGON 44.325 98.085 44.325 98.08 44.54 98.08 44.54 97.76 44.325 97.76 44.325 97.755 43.995 97.755 43.995 97.76 43.78 97.76 43.78 98.08 43.995 98.08 43.995 98.085 ;
      POLYGON 2.03 68.16 2.03 68.15 4.75 68.15 4.75 67.85 2.03 67.85 2.03 67.84 1.65 67.84 1.65 68.16 ;
      POLYGON 44.77 57.95 44.77 57.65 1.23 57.65 1.23 57.93 1.78 57.93 1.78 57.95 ;
      POLYGON 39.71 55.23 39.71 54.93 1.23 54.93 1.23 55.21 1.78 55.21 1.78 55.23 ;
      POLYGON 2.03 24.64 2.03 24.63 6.13 24.63 6.13 24.33 2.03 24.33 2.03 24.32 1.65 24.32 1.65 24.64 ;
      POLYGON 73.765 0.165 73.765 0.16 73.98 0.16 73.98 -0.16 73.765 -0.16 73.765 -0.165 73.435 -0.165 73.435 -0.16 73.22 -0.16 73.22 0.16 73.435 0.16 73.435 0.165 ;
      POLYGON 44.325 0.165 44.325 0.16 44.54 0.16 44.54 -0.16 44.325 -0.16 44.325 -0.165 43.995 -0.165 43.995 -0.16 43.78 -0.16 43.78 0.16 43.995 0.16 43.995 0.165 ;
      POLYGON 84.24 97.52 84.24 0.4 18.8 0.4 18.8 4.89 20.18 4.89 20.18 5.99 18.8 5.99 18.8 6.25 20.18 6.25 20.18 7.35 18.8 7.35 18.8 16.72 0.4 16.72 0.4 19.17 1.78 19.17 1.78 20.27 0.4 20.27 0.4 20.53 1.78 20.53 1.78 21.63 0.4 21.63 0.4 21.89 1.78 21.89 1.78 22.99 0.4 22.99 0.4 23.25 1.78 23.25 1.78 24.35 0.4 24.35 0.4 24.61 1.78 24.61 1.78 25.71 0.4 25.71 0.4 25.97 1.78 25.97 1.78 27.07 0.4 27.07 0.4 27.33 1.78 27.33 1.78 28.43 0.4 28.43 0.4 28.69 1.78 28.69 1.78 29.79 0.4 29.79 0.4 30.05 1.78 30.05 1.78 31.15 0.4 31.15 0.4 31.41 1.78 31.41 1.78 32.51 0.4 32.51 0.4 32.77 1.78 32.77 1.78 33.87 0.4 33.87 0.4 34.13 1.78 34.13 1.78 35.23 0.4 35.23 0.4 35.49 1.78 35.49 1.78 36.59 0.4 36.59 0.4 36.85 1.78 36.85 1.78 37.95 0.4 37.95 0.4 38.21 1.78 38.21 1.78 39.31 0.4 39.31 0.4 39.57 1.78 39.57 1.78 40.67 0.4 40.67 0.4 40.93 1.78 40.93 1.78 42.03 0.4 42.03 0.4 42.29 1.78 42.29 1.78 43.39 0.4 43.39 0.4 43.65 1.78 43.65 1.78 44.75 0.4 44.75 0.4 45.01 1.78 45.01 1.78 46.11 0.4 46.11 0.4 46.37 1.78 46.37 1.78 47.47 0.4 47.47 0.4 48.41 1.78 48.41 1.78 49.51 0.4 49.51 0.4 49.77 1.78 49.77 1.78 50.87 0.4 50.87 0.4 51.13 1.78 51.13 1.78 52.23 0.4 52.23 0.4 52.49 1.78 52.49 1.78 53.59 0.4 53.59 0.4 53.85 1.78 53.85 1.78 54.95 0.4 54.95 0.4 55.21 1.78 55.21 1.78 56.31 0.4 56.31 0.4 56.57 1.78 56.57 1.78 57.67 0.4 57.67 0.4 57.93 1.78 57.93 1.78 59.03 0.4 59.03 0.4 59.29 1.78 59.29 1.78 60.39 0.4 60.39 0.4 60.65 1.78 60.65 1.78 61.75 0.4 61.75 0.4 62.69 1.78 62.69 1.78 63.79 0.4 63.79 0.4 64.05 1.78 64.05 1.78 65.15 0.4 65.15 0.4 65.41 1.78 65.41 1.78 66.51 0.4 66.51 0.4 66.77 1.78 66.77 1.78 67.87 0.4 67.87 0.4 68.13 1.78 68.13 1.78 69.23 0.4 69.23 0.4 69.49 1.78 69.49 1.78 70.59 0.4 70.59 0.4 70.85 1.78 70.85 1.78 71.95 0.4 71.95 0.4 72.89 1.78 72.89 1.78 73.99 0.4 73.99 0.4 74.25 1.78 74.25 1.78 75.35 0.4 75.35 0.4 75.61 1.78 75.61 1.78 76.71 0.4 76.71 0.4 76.97 1.78 76.97 1.78 78.07 0.4 78.07 0.4 81.2 18.8 81.2 18.8 97.52 ;
    LAYER met5 ;
      POLYGON 83.04 96.32 83.04 72.56 79.84 72.56 79.84 66.16 83.04 66.16 83.04 52.16 79.84 52.16 79.84 45.76 83.04 45.76 83.04 31.76 79.84 31.76 79.84 25.36 83.04 25.36 83.04 1.6 20 1.6 20 17.92 1.6 17.92 1.6 25.36 4.8 25.36 4.8 31.76 1.6 31.76 1.6 45.76 4.8 45.76 4.8 52.16 1.6 52.16 1.6 66.16 4.8 66.16 4.8 72.56 1.6 72.56 1.6 80 20 80 20 96.32 ;
    LAYER met1 ;
      POLYGON 84.36 97.4 84.36 95.72 83.88 95.72 83.88 94.68 84.36 94.68 84.36 93 83.88 93 83.88 91.96 84.36 91.96 84.36 90.28 83.88 90.28 83.88 89.24 84.36 89.24 84.36 87.56 83.88 87.56 83.88 86.52 84.36 86.52 84.36 84.84 83.88 84.84 83.88 83.8 84.36 83.8 84.36 82.12 18.68 82.12 18.68 83.8 19.16 83.8 19.16 84.84 18.68 84.84 18.68 86.52 19.16 86.52 19.16 87.56 18.68 87.56 18.68 89.24 19.16 89.24 19.16 90.28 18.68 90.28 18.68 91.96 19.16 91.96 19.16 93 18.68 93 18.68 94.68 19.16 94.68 19.16 95.72 18.68 95.72 18.68 97.4 ;
      POLYGON 84.36 81.08 84.36 79.4 83.88 79.4 83.88 78.36 84.36 78.36 84.36 76.68 83.88 76.68 83.88 75.64 84.36 75.64 84.36 73.96 83.88 73.96 83.88 72.92 84.36 72.92 84.36 71.24 83.88 71.24 83.88 70.2 84.36 70.2 84.36 68.52 83.88 68.52 83.88 67.48 84.36 67.48 84.36 65.8 83.88 65.8 83.88 64.76 84.36 64.76 84.36 63.08 83.88 63.08 83.88 62.04 84.36 62.04 84.36 60.36 83.88 60.36 83.88 59.32 84.36 59.32 84.36 57.64 83.88 57.64 83.88 56.6 84.36 56.6 84.36 54.92 83.88 54.92 83.88 53.88 84.36 53.88 84.36 52.2 83.88 52.2 83.88 51.16 84.36 51.16 84.36 49.48 83.88 49.48 83.88 48.44 84.36 48.44 84.36 46.76 83.88 46.76 83.88 45.72 84.36 45.72 84.36 44.04 83.88 44.04 83.88 43 84.36 43 84.36 41.32 83.88 41.32 83.88 40.28 84.36 40.28 84.36 38.6 83.88 38.6 83.88 37.56 84.36 37.56 84.36 35.88 83.88 35.88 83.88 34.84 84.36 34.84 84.36 33.16 83.88 33.16 83.88 32.12 84.36 32.12 84.36 30.44 83.88 30.44 83.88 29.4 84.36 29.4 84.36 27.72 83.88 27.72 83.88 26.68 84.36 26.68 84.36 25 83.88 25 83.88 23.96 84.36 23.96 84.36 22.28 83.88 22.28 83.88 21.24 84.36 21.24 84.36 19.56 83.88 19.56 83.88 18.52 84.36 18.52 84.36 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 ;
      POLYGON 84.36 15.8 84.36 14.12 83.88 14.12 83.88 13.08 84.36 13.08 84.36 11.4 83.88 11.4 83.88 10.36 84.36 10.36 84.36 8.68 83.88 8.68 83.88 7.64 84.36 7.64 84.36 5.96 83.88 5.96 83.88 4.92 84.36 4.92 84.36 3.24 83.88 3.24 83.88 2.2 84.36 2.2 84.36 0.52 18.68 0.52 18.68 2.2 19.16 2.2 19.16 3.24 18.68 3.24 18.68 4.92 19.16 4.92 19.16 5.96 18.68 5.96 18.68 7.64 19.16 7.64 19.16 8.68 18.68 8.68 18.68 10.36 19.16 10.36 19.16 11.4 18.68 11.4 18.68 13.08 19.16 13.08 19.16 14.12 18.68 14.12 18.68 15.8 ;
    LAYER li1 ;
      POLYGON 84.47 97.75 84.47 0.17 18.57 0.17 18.57 16.49 0.17 16.49 0.17 81.43 18.57 81.43 18.57 97.75 ;
    LAYER mcon ;
      RECT 84.325 97.835 84.495 98.005 ;
      RECT 83.865 97.835 84.035 98.005 ;
      RECT 83.405 97.835 83.575 98.005 ;
      RECT 82.945 97.835 83.115 98.005 ;
      RECT 82.485 97.835 82.655 98.005 ;
      RECT 82.025 97.835 82.195 98.005 ;
      RECT 81.565 97.835 81.735 98.005 ;
      RECT 81.105 97.835 81.275 98.005 ;
      RECT 80.645 97.835 80.815 98.005 ;
      RECT 80.185 97.835 80.355 98.005 ;
      RECT 79.725 97.835 79.895 98.005 ;
      RECT 79.265 97.835 79.435 98.005 ;
      RECT 78.805 97.835 78.975 98.005 ;
      RECT 78.345 97.835 78.515 98.005 ;
      RECT 77.885 97.835 78.055 98.005 ;
      RECT 77.425 97.835 77.595 98.005 ;
      RECT 76.965 97.835 77.135 98.005 ;
      RECT 76.505 97.835 76.675 98.005 ;
      RECT 76.045 97.835 76.215 98.005 ;
      RECT 75.585 97.835 75.755 98.005 ;
      RECT 75.125 97.835 75.295 98.005 ;
      RECT 74.665 97.835 74.835 98.005 ;
      RECT 74.205 97.835 74.375 98.005 ;
      RECT 73.745 97.835 73.915 98.005 ;
      RECT 73.285 97.835 73.455 98.005 ;
      RECT 72.825 97.835 72.995 98.005 ;
      RECT 72.365 97.835 72.535 98.005 ;
      RECT 71.905 97.835 72.075 98.005 ;
      RECT 71.445 97.835 71.615 98.005 ;
      RECT 70.985 97.835 71.155 98.005 ;
      RECT 70.525 97.835 70.695 98.005 ;
      RECT 70.065 97.835 70.235 98.005 ;
      RECT 69.605 97.835 69.775 98.005 ;
      RECT 69.145 97.835 69.315 98.005 ;
      RECT 68.685 97.835 68.855 98.005 ;
      RECT 68.225 97.835 68.395 98.005 ;
      RECT 67.765 97.835 67.935 98.005 ;
      RECT 67.305 97.835 67.475 98.005 ;
      RECT 66.845 97.835 67.015 98.005 ;
      RECT 66.385 97.835 66.555 98.005 ;
      RECT 65.925 97.835 66.095 98.005 ;
      RECT 65.465 97.835 65.635 98.005 ;
      RECT 65.005 97.835 65.175 98.005 ;
      RECT 64.545 97.835 64.715 98.005 ;
      RECT 64.085 97.835 64.255 98.005 ;
      RECT 63.625 97.835 63.795 98.005 ;
      RECT 63.165 97.835 63.335 98.005 ;
      RECT 62.705 97.835 62.875 98.005 ;
      RECT 62.245 97.835 62.415 98.005 ;
      RECT 61.785 97.835 61.955 98.005 ;
      RECT 61.325 97.835 61.495 98.005 ;
      RECT 60.865 97.835 61.035 98.005 ;
      RECT 60.405 97.835 60.575 98.005 ;
      RECT 59.945 97.835 60.115 98.005 ;
      RECT 59.485 97.835 59.655 98.005 ;
      RECT 59.025 97.835 59.195 98.005 ;
      RECT 58.565 97.835 58.735 98.005 ;
      RECT 58.105 97.835 58.275 98.005 ;
      RECT 57.645 97.835 57.815 98.005 ;
      RECT 57.185 97.835 57.355 98.005 ;
      RECT 56.725 97.835 56.895 98.005 ;
      RECT 56.265 97.835 56.435 98.005 ;
      RECT 55.805 97.835 55.975 98.005 ;
      RECT 55.345 97.835 55.515 98.005 ;
      RECT 54.885 97.835 55.055 98.005 ;
      RECT 54.425 97.835 54.595 98.005 ;
      RECT 53.965 97.835 54.135 98.005 ;
      RECT 53.505 97.835 53.675 98.005 ;
      RECT 53.045 97.835 53.215 98.005 ;
      RECT 52.585 97.835 52.755 98.005 ;
      RECT 52.125 97.835 52.295 98.005 ;
      RECT 51.665 97.835 51.835 98.005 ;
      RECT 51.205 97.835 51.375 98.005 ;
      RECT 50.745 97.835 50.915 98.005 ;
      RECT 50.285 97.835 50.455 98.005 ;
      RECT 49.825 97.835 49.995 98.005 ;
      RECT 49.365 97.835 49.535 98.005 ;
      RECT 48.905 97.835 49.075 98.005 ;
      RECT 48.445 97.835 48.615 98.005 ;
      RECT 47.985 97.835 48.155 98.005 ;
      RECT 47.525 97.835 47.695 98.005 ;
      RECT 47.065 97.835 47.235 98.005 ;
      RECT 46.605 97.835 46.775 98.005 ;
      RECT 46.145 97.835 46.315 98.005 ;
      RECT 45.685 97.835 45.855 98.005 ;
      RECT 45.225 97.835 45.395 98.005 ;
      RECT 44.765 97.835 44.935 98.005 ;
      RECT 44.305 97.835 44.475 98.005 ;
      RECT 43.845 97.835 44.015 98.005 ;
      RECT 43.385 97.835 43.555 98.005 ;
      RECT 42.925 97.835 43.095 98.005 ;
      RECT 42.465 97.835 42.635 98.005 ;
      RECT 42.005 97.835 42.175 98.005 ;
      RECT 41.545 97.835 41.715 98.005 ;
      RECT 41.085 97.835 41.255 98.005 ;
      RECT 40.625 97.835 40.795 98.005 ;
      RECT 40.165 97.835 40.335 98.005 ;
      RECT 39.705 97.835 39.875 98.005 ;
      RECT 39.245 97.835 39.415 98.005 ;
      RECT 38.785 97.835 38.955 98.005 ;
      RECT 38.325 97.835 38.495 98.005 ;
      RECT 37.865 97.835 38.035 98.005 ;
      RECT 37.405 97.835 37.575 98.005 ;
      RECT 36.945 97.835 37.115 98.005 ;
      RECT 36.485 97.835 36.655 98.005 ;
      RECT 36.025 97.835 36.195 98.005 ;
      RECT 35.565 97.835 35.735 98.005 ;
      RECT 35.105 97.835 35.275 98.005 ;
      RECT 34.645 97.835 34.815 98.005 ;
      RECT 34.185 97.835 34.355 98.005 ;
      RECT 33.725 97.835 33.895 98.005 ;
      RECT 33.265 97.835 33.435 98.005 ;
      RECT 32.805 97.835 32.975 98.005 ;
      RECT 32.345 97.835 32.515 98.005 ;
      RECT 31.885 97.835 32.055 98.005 ;
      RECT 31.425 97.835 31.595 98.005 ;
      RECT 30.965 97.835 31.135 98.005 ;
      RECT 30.505 97.835 30.675 98.005 ;
      RECT 30.045 97.835 30.215 98.005 ;
      RECT 29.585 97.835 29.755 98.005 ;
      RECT 29.125 97.835 29.295 98.005 ;
      RECT 28.665 97.835 28.835 98.005 ;
      RECT 28.205 97.835 28.375 98.005 ;
      RECT 27.745 97.835 27.915 98.005 ;
      RECT 27.285 97.835 27.455 98.005 ;
      RECT 26.825 97.835 26.995 98.005 ;
      RECT 26.365 97.835 26.535 98.005 ;
      RECT 25.905 97.835 26.075 98.005 ;
      RECT 25.445 97.835 25.615 98.005 ;
      RECT 24.985 97.835 25.155 98.005 ;
      RECT 24.525 97.835 24.695 98.005 ;
      RECT 24.065 97.835 24.235 98.005 ;
      RECT 23.605 97.835 23.775 98.005 ;
      RECT 23.145 97.835 23.315 98.005 ;
      RECT 22.685 97.835 22.855 98.005 ;
      RECT 22.225 97.835 22.395 98.005 ;
      RECT 21.765 97.835 21.935 98.005 ;
      RECT 21.305 97.835 21.475 98.005 ;
      RECT 20.845 97.835 21.015 98.005 ;
      RECT 20.385 97.835 20.555 98.005 ;
      RECT 19.925 97.835 20.095 98.005 ;
      RECT 19.465 97.835 19.635 98.005 ;
      RECT 19.005 97.835 19.175 98.005 ;
      RECT 18.545 97.835 18.715 98.005 ;
      RECT 84.325 95.115 84.495 95.285 ;
      RECT 83.865 95.115 84.035 95.285 ;
      RECT 19.005 95.115 19.175 95.285 ;
      RECT 18.545 95.115 18.715 95.285 ;
      RECT 84.325 92.395 84.495 92.565 ;
      RECT 83.865 92.395 84.035 92.565 ;
      RECT 19.005 92.395 19.175 92.565 ;
      RECT 18.545 92.395 18.715 92.565 ;
      RECT 84.325 89.675 84.495 89.845 ;
      RECT 83.865 89.675 84.035 89.845 ;
      RECT 19.005 89.675 19.175 89.845 ;
      RECT 18.545 89.675 18.715 89.845 ;
      RECT 84.325 86.955 84.495 87.125 ;
      RECT 83.865 86.955 84.035 87.125 ;
      RECT 19.005 86.955 19.175 87.125 ;
      RECT 18.545 86.955 18.715 87.125 ;
      RECT 84.325 84.235 84.495 84.405 ;
      RECT 83.865 84.235 84.035 84.405 ;
      RECT 19.005 84.235 19.175 84.405 ;
      RECT 18.545 84.235 18.715 84.405 ;
      RECT 84.325 81.515 84.495 81.685 ;
      RECT 83.865 81.515 84.035 81.685 ;
      RECT 83.405 81.515 83.575 81.685 ;
      RECT 82.945 81.515 83.115 81.685 ;
      RECT 82.485 81.515 82.655 81.685 ;
      RECT 82.025 81.515 82.195 81.685 ;
      RECT 81.565 81.515 81.735 81.685 ;
      RECT 81.105 81.515 81.275 81.685 ;
      RECT 80.645 81.515 80.815 81.685 ;
      RECT 80.185 81.515 80.355 81.685 ;
      RECT 79.725 81.515 79.895 81.685 ;
      RECT 79.265 81.515 79.435 81.685 ;
      RECT 78.805 81.515 78.975 81.685 ;
      RECT 78.345 81.515 78.515 81.685 ;
      RECT 77.885 81.515 78.055 81.685 ;
      RECT 77.425 81.515 77.595 81.685 ;
      RECT 76.965 81.515 77.135 81.685 ;
      RECT 76.505 81.515 76.675 81.685 ;
      RECT 76.045 81.515 76.215 81.685 ;
      RECT 75.585 81.515 75.755 81.685 ;
      RECT 75.125 81.515 75.295 81.685 ;
      RECT 74.665 81.515 74.835 81.685 ;
      RECT 74.205 81.515 74.375 81.685 ;
      RECT 73.745 81.515 73.915 81.685 ;
      RECT 73.285 81.515 73.455 81.685 ;
      RECT 72.825 81.515 72.995 81.685 ;
      RECT 72.365 81.515 72.535 81.685 ;
      RECT 71.905 81.515 72.075 81.685 ;
      RECT 71.445 81.515 71.615 81.685 ;
      RECT 70.985 81.515 71.155 81.685 ;
      RECT 70.525 81.515 70.695 81.685 ;
      RECT 70.065 81.515 70.235 81.685 ;
      RECT 69.605 81.515 69.775 81.685 ;
      RECT 69.145 81.515 69.315 81.685 ;
      RECT 68.685 81.515 68.855 81.685 ;
      RECT 68.225 81.515 68.395 81.685 ;
      RECT 67.765 81.515 67.935 81.685 ;
      RECT 67.305 81.515 67.475 81.685 ;
      RECT 66.845 81.515 67.015 81.685 ;
      RECT 66.385 81.515 66.555 81.685 ;
      RECT 65.925 81.515 66.095 81.685 ;
      RECT 65.465 81.515 65.635 81.685 ;
      RECT 65.005 81.515 65.175 81.685 ;
      RECT 64.545 81.515 64.715 81.685 ;
      RECT 64.085 81.515 64.255 81.685 ;
      RECT 63.625 81.515 63.795 81.685 ;
      RECT 63.165 81.515 63.335 81.685 ;
      RECT 62.705 81.515 62.875 81.685 ;
      RECT 62.245 81.515 62.415 81.685 ;
      RECT 61.785 81.515 61.955 81.685 ;
      RECT 61.325 81.515 61.495 81.685 ;
      RECT 60.865 81.515 61.035 81.685 ;
      RECT 60.405 81.515 60.575 81.685 ;
      RECT 59.945 81.515 60.115 81.685 ;
      RECT 59.485 81.515 59.655 81.685 ;
      RECT 59.025 81.515 59.195 81.685 ;
      RECT 58.565 81.515 58.735 81.685 ;
      RECT 58.105 81.515 58.275 81.685 ;
      RECT 57.645 81.515 57.815 81.685 ;
      RECT 57.185 81.515 57.355 81.685 ;
      RECT 56.725 81.515 56.895 81.685 ;
      RECT 56.265 81.515 56.435 81.685 ;
      RECT 55.805 81.515 55.975 81.685 ;
      RECT 55.345 81.515 55.515 81.685 ;
      RECT 54.885 81.515 55.055 81.685 ;
      RECT 54.425 81.515 54.595 81.685 ;
      RECT 53.965 81.515 54.135 81.685 ;
      RECT 53.505 81.515 53.675 81.685 ;
      RECT 53.045 81.515 53.215 81.685 ;
      RECT 52.585 81.515 52.755 81.685 ;
      RECT 52.125 81.515 52.295 81.685 ;
      RECT 51.665 81.515 51.835 81.685 ;
      RECT 51.205 81.515 51.375 81.685 ;
      RECT 50.745 81.515 50.915 81.685 ;
      RECT 50.285 81.515 50.455 81.685 ;
      RECT 49.825 81.515 49.995 81.685 ;
      RECT 49.365 81.515 49.535 81.685 ;
      RECT 48.905 81.515 49.075 81.685 ;
      RECT 48.445 81.515 48.615 81.685 ;
      RECT 47.985 81.515 48.155 81.685 ;
      RECT 47.525 81.515 47.695 81.685 ;
      RECT 47.065 81.515 47.235 81.685 ;
      RECT 46.605 81.515 46.775 81.685 ;
      RECT 46.145 81.515 46.315 81.685 ;
      RECT 45.685 81.515 45.855 81.685 ;
      RECT 45.225 81.515 45.395 81.685 ;
      RECT 44.765 81.515 44.935 81.685 ;
      RECT 44.305 81.515 44.475 81.685 ;
      RECT 43.845 81.515 44.015 81.685 ;
      RECT 43.385 81.515 43.555 81.685 ;
      RECT 42.925 81.515 43.095 81.685 ;
      RECT 42.465 81.515 42.635 81.685 ;
      RECT 42.005 81.515 42.175 81.685 ;
      RECT 41.545 81.515 41.715 81.685 ;
      RECT 41.085 81.515 41.255 81.685 ;
      RECT 40.625 81.515 40.795 81.685 ;
      RECT 40.165 81.515 40.335 81.685 ;
      RECT 39.705 81.515 39.875 81.685 ;
      RECT 39.245 81.515 39.415 81.685 ;
      RECT 38.785 81.515 38.955 81.685 ;
      RECT 38.325 81.515 38.495 81.685 ;
      RECT 37.865 81.515 38.035 81.685 ;
      RECT 37.405 81.515 37.575 81.685 ;
      RECT 36.945 81.515 37.115 81.685 ;
      RECT 36.485 81.515 36.655 81.685 ;
      RECT 36.025 81.515 36.195 81.685 ;
      RECT 35.565 81.515 35.735 81.685 ;
      RECT 35.105 81.515 35.275 81.685 ;
      RECT 34.645 81.515 34.815 81.685 ;
      RECT 34.185 81.515 34.355 81.685 ;
      RECT 33.725 81.515 33.895 81.685 ;
      RECT 33.265 81.515 33.435 81.685 ;
      RECT 32.805 81.515 32.975 81.685 ;
      RECT 32.345 81.515 32.515 81.685 ;
      RECT 31.885 81.515 32.055 81.685 ;
      RECT 31.425 81.515 31.595 81.685 ;
      RECT 30.965 81.515 31.135 81.685 ;
      RECT 30.505 81.515 30.675 81.685 ;
      RECT 30.045 81.515 30.215 81.685 ;
      RECT 29.585 81.515 29.755 81.685 ;
      RECT 29.125 81.515 29.295 81.685 ;
      RECT 28.665 81.515 28.835 81.685 ;
      RECT 28.205 81.515 28.375 81.685 ;
      RECT 27.745 81.515 27.915 81.685 ;
      RECT 27.285 81.515 27.455 81.685 ;
      RECT 26.825 81.515 26.995 81.685 ;
      RECT 26.365 81.515 26.535 81.685 ;
      RECT 25.905 81.515 26.075 81.685 ;
      RECT 25.445 81.515 25.615 81.685 ;
      RECT 24.985 81.515 25.155 81.685 ;
      RECT 24.525 81.515 24.695 81.685 ;
      RECT 24.065 81.515 24.235 81.685 ;
      RECT 23.605 81.515 23.775 81.685 ;
      RECT 23.145 81.515 23.315 81.685 ;
      RECT 22.685 81.515 22.855 81.685 ;
      RECT 22.225 81.515 22.395 81.685 ;
      RECT 21.765 81.515 21.935 81.685 ;
      RECT 21.305 81.515 21.475 81.685 ;
      RECT 20.845 81.515 21.015 81.685 ;
      RECT 20.385 81.515 20.555 81.685 ;
      RECT 19.925 81.515 20.095 81.685 ;
      RECT 19.465 81.515 19.635 81.685 ;
      RECT 19.005 81.515 19.175 81.685 ;
      RECT 18.545 81.515 18.715 81.685 ;
      RECT 18.085 81.515 18.255 81.685 ;
      RECT 17.625 81.515 17.795 81.685 ;
      RECT 17.165 81.515 17.335 81.685 ;
      RECT 16.705 81.515 16.875 81.685 ;
      RECT 16.245 81.515 16.415 81.685 ;
      RECT 15.785 81.515 15.955 81.685 ;
      RECT 15.325 81.515 15.495 81.685 ;
      RECT 14.865 81.515 15.035 81.685 ;
      RECT 14.405 81.515 14.575 81.685 ;
      RECT 13.945 81.515 14.115 81.685 ;
      RECT 13.485 81.515 13.655 81.685 ;
      RECT 13.025 81.515 13.195 81.685 ;
      RECT 12.565 81.515 12.735 81.685 ;
      RECT 12.105 81.515 12.275 81.685 ;
      RECT 11.645 81.515 11.815 81.685 ;
      RECT 11.185 81.515 11.355 81.685 ;
      RECT 10.725 81.515 10.895 81.685 ;
      RECT 10.265 81.515 10.435 81.685 ;
      RECT 9.805 81.515 9.975 81.685 ;
      RECT 9.345 81.515 9.515 81.685 ;
      RECT 8.885 81.515 9.055 81.685 ;
      RECT 8.425 81.515 8.595 81.685 ;
      RECT 7.965 81.515 8.135 81.685 ;
      RECT 7.505 81.515 7.675 81.685 ;
      RECT 7.045 81.515 7.215 81.685 ;
      RECT 6.585 81.515 6.755 81.685 ;
      RECT 6.125 81.515 6.295 81.685 ;
      RECT 5.665 81.515 5.835 81.685 ;
      RECT 5.205 81.515 5.375 81.685 ;
      RECT 4.745 81.515 4.915 81.685 ;
      RECT 4.285 81.515 4.455 81.685 ;
      RECT 3.825 81.515 3.995 81.685 ;
      RECT 3.365 81.515 3.535 81.685 ;
      RECT 2.905 81.515 3.075 81.685 ;
      RECT 2.445 81.515 2.615 81.685 ;
      RECT 1.985 81.515 2.155 81.685 ;
      RECT 1.525 81.515 1.695 81.685 ;
      RECT 1.065 81.515 1.235 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 84.325 78.795 84.495 78.965 ;
      RECT 83.865 78.795 84.035 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 84.325 76.075 84.495 76.245 ;
      RECT 83.865 76.075 84.035 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 84.325 73.355 84.495 73.525 ;
      RECT 83.865 73.355 84.035 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 84.325 70.635 84.495 70.805 ;
      RECT 83.865 70.635 84.035 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 84.325 67.915 84.495 68.085 ;
      RECT 83.865 67.915 84.035 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 84.325 65.195 84.495 65.365 ;
      RECT 83.865 65.195 84.035 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 84.325 62.475 84.495 62.645 ;
      RECT 83.865 62.475 84.035 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 84.325 59.755 84.495 59.925 ;
      RECT 83.865 59.755 84.035 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 84.325 57.035 84.495 57.205 ;
      RECT 83.865 57.035 84.035 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 84.325 54.315 84.495 54.485 ;
      RECT 83.865 54.315 84.035 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 84.325 51.595 84.495 51.765 ;
      RECT 83.865 51.595 84.035 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 84.325 48.875 84.495 49.045 ;
      RECT 83.865 48.875 84.035 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 84.325 46.155 84.495 46.325 ;
      RECT 83.865 46.155 84.035 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 84.325 43.435 84.495 43.605 ;
      RECT 83.865 43.435 84.035 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 84.325 40.715 84.495 40.885 ;
      RECT 83.865 40.715 84.035 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 84.325 37.995 84.495 38.165 ;
      RECT 83.865 37.995 84.035 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 84.325 35.275 84.495 35.445 ;
      RECT 83.865 35.275 84.035 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 84.325 32.555 84.495 32.725 ;
      RECT 83.865 32.555 84.035 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 84.325 29.835 84.495 30.005 ;
      RECT 83.865 29.835 84.035 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 84.325 27.115 84.495 27.285 ;
      RECT 83.865 27.115 84.035 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 84.325 24.395 84.495 24.565 ;
      RECT 83.865 24.395 84.035 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 84.325 21.675 84.495 21.845 ;
      RECT 83.865 21.675 84.035 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 84.325 18.955 84.495 19.125 ;
      RECT 83.865 18.955 84.035 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 84.325 16.235 84.495 16.405 ;
      RECT 83.865 16.235 84.035 16.405 ;
      RECT 83.405 16.235 83.575 16.405 ;
      RECT 82.945 16.235 83.115 16.405 ;
      RECT 82.485 16.235 82.655 16.405 ;
      RECT 82.025 16.235 82.195 16.405 ;
      RECT 81.565 16.235 81.735 16.405 ;
      RECT 81.105 16.235 81.275 16.405 ;
      RECT 80.645 16.235 80.815 16.405 ;
      RECT 80.185 16.235 80.355 16.405 ;
      RECT 79.725 16.235 79.895 16.405 ;
      RECT 79.265 16.235 79.435 16.405 ;
      RECT 78.805 16.235 78.975 16.405 ;
      RECT 78.345 16.235 78.515 16.405 ;
      RECT 77.885 16.235 78.055 16.405 ;
      RECT 77.425 16.235 77.595 16.405 ;
      RECT 76.965 16.235 77.135 16.405 ;
      RECT 76.505 16.235 76.675 16.405 ;
      RECT 76.045 16.235 76.215 16.405 ;
      RECT 75.585 16.235 75.755 16.405 ;
      RECT 75.125 16.235 75.295 16.405 ;
      RECT 74.665 16.235 74.835 16.405 ;
      RECT 74.205 16.235 74.375 16.405 ;
      RECT 73.745 16.235 73.915 16.405 ;
      RECT 73.285 16.235 73.455 16.405 ;
      RECT 72.825 16.235 72.995 16.405 ;
      RECT 72.365 16.235 72.535 16.405 ;
      RECT 71.905 16.235 72.075 16.405 ;
      RECT 71.445 16.235 71.615 16.405 ;
      RECT 70.985 16.235 71.155 16.405 ;
      RECT 70.525 16.235 70.695 16.405 ;
      RECT 70.065 16.235 70.235 16.405 ;
      RECT 69.605 16.235 69.775 16.405 ;
      RECT 69.145 16.235 69.315 16.405 ;
      RECT 68.685 16.235 68.855 16.405 ;
      RECT 68.225 16.235 68.395 16.405 ;
      RECT 67.765 16.235 67.935 16.405 ;
      RECT 67.305 16.235 67.475 16.405 ;
      RECT 66.845 16.235 67.015 16.405 ;
      RECT 66.385 16.235 66.555 16.405 ;
      RECT 65.925 16.235 66.095 16.405 ;
      RECT 65.465 16.235 65.635 16.405 ;
      RECT 65.005 16.235 65.175 16.405 ;
      RECT 64.545 16.235 64.715 16.405 ;
      RECT 64.085 16.235 64.255 16.405 ;
      RECT 63.625 16.235 63.795 16.405 ;
      RECT 63.165 16.235 63.335 16.405 ;
      RECT 62.705 16.235 62.875 16.405 ;
      RECT 62.245 16.235 62.415 16.405 ;
      RECT 61.785 16.235 61.955 16.405 ;
      RECT 61.325 16.235 61.495 16.405 ;
      RECT 60.865 16.235 61.035 16.405 ;
      RECT 60.405 16.235 60.575 16.405 ;
      RECT 59.945 16.235 60.115 16.405 ;
      RECT 59.485 16.235 59.655 16.405 ;
      RECT 59.025 16.235 59.195 16.405 ;
      RECT 58.565 16.235 58.735 16.405 ;
      RECT 58.105 16.235 58.275 16.405 ;
      RECT 57.645 16.235 57.815 16.405 ;
      RECT 57.185 16.235 57.355 16.405 ;
      RECT 56.725 16.235 56.895 16.405 ;
      RECT 56.265 16.235 56.435 16.405 ;
      RECT 55.805 16.235 55.975 16.405 ;
      RECT 55.345 16.235 55.515 16.405 ;
      RECT 54.885 16.235 55.055 16.405 ;
      RECT 54.425 16.235 54.595 16.405 ;
      RECT 53.965 16.235 54.135 16.405 ;
      RECT 53.505 16.235 53.675 16.405 ;
      RECT 53.045 16.235 53.215 16.405 ;
      RECT 52.585 16.235 52.755 16.405 ;
      RECT 52.125 16.235 52.295 16.405 ;
      RECT 51.665 16.235 51.835 16.405 ;
      RECT 51.205 16.235 51.375 16.405 ;
      RECT 50.745 16.235 50.915 16.405 ;
      RECT 50.285 16.235 50.455 16.405 ;
      RECT 49.825 16.235 49.995 16.405 ;
      RECT 49.365 16.235 49.535 16.405 ;
      RECT 48.905 16.235 49.075 16.405 ;
      RECT 48.445 16.235 48.615 16.405 ;
      RECT 47.985 16.235 48.155 16.405 ;
      RECT 47.525 16.235 47.695 16.405 ;
      RECT 47.065 16.235 47.235 16.405 ;
      RECT 46.605 16.235 46.775 16.405 ;
      RECT 46.145 16.235 46.315 16.405 ;
      RECT 45.685 16.235 45.855 16.405 ;
      RECT 45.225 16.235 45.395 16.405 ;
      RECT 44.765 16.235 44.935 16.405 ;
      RECT 44.305 16.235 44.475 16.405 ;
      RECT 43.845 16.235 44.015 16.405 ;
      RECT 43.385 16.235 43.555 16.405 ;
      RECT 42.925 16.235 43.095 16.405 ;
      RECT 42.465 16.235 42.635 16.405 ;
      RECT 42.005 16.235 42.175 16.405 ;
      RECT 41.545 16.235 41.715 16.405 ;
      RECT 41.085 16.235 41.255 16.405 ;
      RECT 40.625 16.235 40.795 16.405 ;
      RECT 40.165 16.235 40.335 16.405 ;
      RECT 39.705 16.235 39.875 16.405 ;
      RECT 39.245 16.235 39.415 16.405 ;
      RECT 38.785 16.235 38.955 16.405 ;
      RECT 38.325 16.235 38.495 16.405 ;
      RECT 37.865 16.235 38.035 16.405 ;
      RECT 37.405 16.235 37.575 16.405 ;
      RECT 36.945 16.235 37.115 16.405 ;
      RECT 36.485 16.235 36.655 16.405 ;
      RECT 36.025 16.235 36.195 16.405 ;
      RECT 35.565 16.235 35.735 16.405 ;
      RECT 35.105 16.235 35.275 16.405 ;
      RECT 34.645 16.235 34.815 16.405 ;
      RECT 34.185 16.235 34.355 16.405 ;
      RECT 33.725 16.235 33.895 16.405 ;
      RECT 33.265 16.235 33.435 16.405 ;
      RECT 32.805 16.235 32.975 16.405 ;
      RECT 32.345 16.235 32.515 16.405 ;
      RECT 31.885 16.235 32.055 16.405 ;
      RECT 31.425 16.235 31.595 16.405 ;
      RECT 30.965 16.235 31.135 16.405 ;
      RECT 30.505 16.235 30.675 16.405 ;
      RECT 30.045 16.235 30.215 16.405 ;
      RECT 29.585 16.235 29.755 16.405 ;
      RECT 29.125 16.235 29.295 16.405 ;
      RECT 28.665 16.235 28.835 16.405 ;
      RECT 28.205 16.235 28.375 16.405 ;
      RECT 27.745 16.235 27.915 16.405 ;
      RECT 27.285 16.235 27.455 16.405 ;
      RECT 26.825 16.235 26.995 16.405 ;
      RECT 26.365 16.235 26.535 16.405 ;
      RECT 25.905 16.235 26.075 16.405 ;
      RECT 25.445 16.235 25.615 16.405 ;
      RECT 24.985 16.235 25.155 16.405 ;
      RECT 24.525 16.235 24.695 16.405 ;
      RECT 24.065 16.235 24.235 16.405 ;
      RECT 23.605 16.235 23.775 16.405 ;
      RECT 23.145 16.235 23.315 16.405 ;
      RECT 22.685 16.235 22.855 16.405 ;
      RECT 22.225 16.235 22.395 16.405 ;
      RECT 21.765 16.235 21.935 16.405 ;
      RECT 21.305 16.235 21.475 16.405 ;
      RECT 20.845 16.235 21.015 16.405 ;
      RECT 20.385 16.235 20.555 16.405 ;
      RECT 19.925 16.235 20.095 16.405 ;
      RECT 19.465 16.235 19.635 16.405 ;
      RECT 19.005 16.235 19.175 16.405 ;
      RECT 18.545 16.235 18.715 16.405 ;
      RECT 18.085 16.235 18.255 16.405 ;
      RECT 17.625 16.235 17.795 16.405 ;
      RECT 17.165 16.235 17.335 16.405 ;
      RECT 16.705 16.235 16.875 16.405 ;
      RECT 16.245 16.235 16.415 16.405 ;
      RECT 15.785 16.235 15.955 16.405 ;
      RECT 15.325 16.235 15.495 16.405 ;
      RECT 14.865 16.235 15.035 16.405 ;
      RECT 14.405 16.235 14.575 16.405 ;
      RECT 13.945 16.235 14.115 16.405 ;
      RECT 13.485 16.235 13.655 16.405 ;
      RECT 13.025 16.235 13.195 16.405 ;
      RECT 12.565 16.235 12.735 16.405 ;
      RECT 12.105 16.235 12.275 16.405 ;
      RECT 11.645 16.235 11.815 16.405 ;
      RECT 11.185 16.235 11.355 16.405 ;
      RECT 10.725 16.235 10.895 16.405 ;
      RECT 10.265 16.235 10.435 16.405 ;
      RECT 9.805 16.235 9.975 16.405 ;
      RECT 9.345 16.235 9.515 16.405 ;
      RECT 8.885 16.235 9.055 16.405 ;
      RECT 8.425 16.235 8.595 16.405 ;
      RECT 7.965 16.235 8.135 16.405 ;
      RECT 7.505 16.235 7.675 16.405 ;
      RECT 7.045 16.235 7.215 16.405 ;
      RECT 6.585 16.235 6.755 16.405 ;
      RECT 6.125 16.235 6.295 16.405 ;
      RECT 5.665 16.235 5.835 16.405 ;
      RECT 5.205 16.235 5.375 16.405 ;
      RECT 4.745 16.235 4.915 16.405 ;
      RECT 4.285 16.235 4.455 16.405 ;
      RECT 3.825 16.235 3.995 16.405 ;
      RECT 3.365 16.235 3.535 16.405 ;
      RECT 2.905 16.235 3.075 16.405 ;
      RECT 2.445 16.235 2.615 16.405 ;
      RECT 1.985 16.235 2.155 16.405 ;
      RECT 1.525 16.235 1.695 16.405 ;
      RECT 1.065 16.235 1.235 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 84.325 13.515 84.495 13.685 ;
      RECT 83.865 13.515 84.035 13.685 ;
      RECT 19.005 13.515 19.175 13.685 ;
      RECT 18.545 13.515 18.715 13.685 ;
      RECT 84.325 10.795 84.495 10.965 ;
      RECT 83.865 10.795 84.035 10.965 ;
      RECT 19.005 10.795 19.175 10.965 ;
      RECT 18.545 10.795 18.715 10.965 ;
      RECT 84.325 8.075 84.495 8.245 ;
      RECT 83.865 8.075 84.035 8.245 ;
      RECT 19.005 8.075 19.175 8.245 ;
      RECT 18.545 8.075 18.715 8.245 ;
      RECT 84.325 5.355 84.495 5.525 ;
      RECT 83.865 5.355 84.035 5.525 ;
      RECT 19.005 5.355 19.175 5.525 ;
      RECT 18.545 5.355 18.715 5.525 ;
      RECT 84.325 2.635 84.495 2.805 ;
      RECT 83.865 2.635 84.035 2.805 ;
      RECT 19.005 2.635 19.175 2.805 ;
      RECT 18.545 2.635 18.715 2.805 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
    LAYER via ;
      RECT 73.525 97.845 73.675 97.995 ;
      RECT 44.085 97.845 44.235 97.995 ;
      RECT 59.265 96.145 59.415 96.295 ;
      RECT 40.865 96.145 41.015 96.295 ;
      RECT 73.525 81.525 73.675 81.675 ;
      RECT 44.085 81.525 44.235 81.675 ;
      RECT 13.265 79.825 13.415 79.975 ;
      RECT 5.445 17.945 5.595 18.095 ;
      RECT 73.525 16.245 73.675 16.395 ;
      RECT 44.085 16.245 44.235 16.395 ;
      RECT 37.645 1.625 37.795 1.775 ;
      RECT 24.765 1.625 24.915 1.775 ;
      RECT 73.525 -0.075 73.675 0.075 ;
      RECT 44.085 -0.075 44.235 0.075 ;
    LAYER via2 ;
      RECT 73.5 97.82 73.7 98.02 ;
      RECT 44.06 97.82 44.26 98.02 ;
      RECT 1.28 73.34 1.48 73.54 ;
      RECT 1.74 61.1 1.94 61.3 ;
      RECT 1.74 46.82 1.94 47.02 ;
      RECT 1.28 25.06 1.48 25.26 ;
      RECT 19.68 5.34 19.88 5.54 ;
      RECT 73.5 -0.1 73.7 0.1 ;
      RECT 44.06 -0.1 44.26 0.1 ;
    LAYER via3 ;
      RECT 73.5 97.82 73.7 98.02 ;
      RECT 44.06 97.82 44.26 98.02 ;
      RECT 1.74 30.5 1.94 30.7 ;
      RECT 1.74 26.42 1.94 26.62 ;
      RECT 73.5 -0.1 73.7 0.1 ;
      RECT 44.06 -0.1 44.26 0.1 ;
    LAYER OVERLAP ;
      POLYGON 18.4 0 18.4 16.32 0 16.32 0 81.6 18.4 81.6 18.4 97.92 84.64 97.92 84.64 0 ;
  END
END sb_2__1_

END LIBRARY
