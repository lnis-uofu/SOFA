//
//
//
//
//
//
module fpga_top ( vdda1 , vdda2 , vssa1 , vssa2 , vccd1 , vccd2 , vssd1 , 
    vssd2 , wb_clk_i , wb_rst_i , wbs_stb_i , wbs_cyc_i , wbs_we_i , 
    wbs_sel_i , wbs_dat_i , wbs_adr_i , wbs_ack_o , wbs_dat_o , la_data_in , 
    la_data_out , la_oen , io_in , io_out , io_oeb , analog_io_0_ , 
    analog_io_10_ , analog_io_11_ , analog_io_12_ , analog_io_13_ , 
    analog_io_14_ , analog_io_15_ , analog_io_16_ , analog_io_17_ , 
    analog_io_18_ , analog_io_19_ , analog_io_1_ , analog_io_20_ , 
    analog_io_21_ , analog_io_22_ , analog_io_23_ , analog_io_24_ , 
    analog_io_25_ , analog_io_26_ , analog_io_27_ , analog_io_28_ , 
    analog_io_29_ , analog_io_2_ , analog_io_30_ , analog_io_3_ , 
    analog_io_4_ , analog_io_5_ , analog_io_6_ , analog_io_7_ , analog_io_8_ , 
    analog_io_9_ , user_clock2 ) ;
inout  vdda1 ;
inout  vdda2 ;
inout  vssa1 ;
inout  vssa2 ;
inout  vccd1 ;
inout  vccd2 ;
inout  vssd1 ;
inout  vssd2 ;
input  wb_clk_i ;
input  wb_rst_i ;
input  wbs_stb_i ;
input  wbs_cyc_i ;
input  wbs_we_i ;
input  [3:0] wbs_sel_i ;
input  [31:0] wbs_dat_i ;
input  [31:0] wbs_adr_i ;
output wbs_ack_o ;
output [31:0] wbs_dat_o ;
input  [127:0] la_data_in ;
output [127:0] la_data_out ;
input  [127:0] la_oen ;
input  [37:0] io_in ;
output [37:0] io_out ;
output [37:0] io_oeb ;
inout  analog_io_0_ ;
inout  analog_io_10_ ;
inout  analog_io_11_ ;
inout  analog_io_12_ ;
inout  analog_io_13_ ;
inout  analog_io_14_ ;
inout  analog_io_15_ ;
inout  analog_io_16_ ;
inout  analog_io_17_ ;
inout  analog_io_18_ ;
inout  analog_io_19_ ;
inout  analog_io_1_ ;
inout  analog_io_20_ ;
inout  analog_io_21_ ;
inout  analog_io_22_ ;
inout  analog_io_23_ ;
inout  analog_io_24_ ;
inout  analog_io_25_ ;
inout  analog_io_26_ ;
inout  analog_io_27_ ;
inout  analog_io_28_ ;
inout  analog_io_29_ ;
inout  analog_io_2_ ;
inout  analog_io_30_ ;
inout  analog_io_3_ ;
inout  analog_io_4_ ;
inout  analog_io_5_ ;
inout  analog_io_6_ ;
inout  analog_io_7_ ;
inout  analog_io_8_ ;
inout  analog_io_9_ ;
input  user_clock2 ;

wire [0:143] gfpga_pad_EMBEDDED_IO_HD_SOC_IN ;
wire [0:143] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT ;
wire [0:143] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR ;
wire ccff_head ;
wire sc_tail ;
wire pReset ;
wire Reset ;
wire IO_ISOL_N ;
wire Test_en ;
wire prog_clk ;
wire clk ;
wire ccff_tail ;
wire sc_head ;
wire wb_la_switch ;

assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0] = io_in[24] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0] = io_out[24] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0] = io_oeb[24] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1] = io_in[23] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1] = io_out[23] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1] = io_oeb[23] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2] = io_in[22] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2] = io_out[22] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2] = io_oeb[22] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3] = io_in[21] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3] = io_out[21] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3] = io_oeb[21] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4] = io_in[20] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4] = io_out[20] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4] = io_oeb[20] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5] = io_in[19] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5] = io_out[19] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5] = io_oeb[19] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6] = io_in[18] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6] = io_out[18] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6] = io_oeb[18] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7] = io_in[17] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7] = io_out[17] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7] = io_oeb[17] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8] = io_in[16] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8] = io_out[16] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8] = io_oeb[16] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9] = io_in[15] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9] = io_out[15] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9] = io_oeb[15] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10] = io_in[14] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10] = io_out[14] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10] = io_oeb[14] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11] = io_in[13] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11] = io_out[13] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11] = io_oeb[13] ;
assign ccff_head = io_in[12] ;
assign sc_tail = io_out[11] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12] = io_in[10] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12] = io_out[10] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12] = io_oeb[10] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13] = io_in[9] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13] = io_out[9] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13] = io_oeb[9] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14] = io_in[8] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14] = io_out[8] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14] = io_oeb[8] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15] = io_in[7] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15] = io_out[7] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15] = io_oeb[7] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16] = io_in[6] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16] = io_out[6] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16] = io_oeb[6] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17] = io_in[5] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17] = io_out[5] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17] = io_oeb[5] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18] = io_in[4] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18] = io_out[4] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18] = io_oeb[4] ;
assign pReset = io_in[3] ;
assign Reset = io_in[2] ;
assign IO_ISOL_N = io_in[1] ;
assign Test_en = io_in[0] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19] = la_data_in[127] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19] = la_data_out[127] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20] = la_data_in[126] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20] = la_data_out[126] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21] = la_data_in[125] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21] = la_data_out[125] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22] = la_data_in[124] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22] = la_data_out[124] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23] = la_data_in[123] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23] = la_data_out[123] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24] = la_data_in[122] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24] = la_data_out[122] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25] = la_data_in[121] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25] = la_data_out[121] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26] = la_data_in[120] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26] = la_data_out[120] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27] = la_data_in[119] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27] = la_data_out[119] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28] = la_data_in[118] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28] = la_data_out[118] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29] = la_data_in[117] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29] = la_data_out[117] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30] = la_data_in[116] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31] = la_data_in[115] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32] = la_data_in[114] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33] = la_data_in[113] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34] = la_data_in[112] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35] = la_data_in[111] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36] = la_data_in[110] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37] = la_data_in[109] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38] = la_data_in[108] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39] = la_data_in[107] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40] = la_data_in[106] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41] = la_data_in[105] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42] = la_data_in[104] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43] = la_data_in[103] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44] = la_data_in[102] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45] = la_data_in[101] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46] = la_data_in[100] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47] = la_data_in[99] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48] = la_data_in[98] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49] = la_data_in[97] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50] = la_data_in[96] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51] = la_data_in[95] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52] = la_data_in[94] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53] = la_data_in[93] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54] = la_data_in[92] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55] = la_data_in[91] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56] = la_data_in[90] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57] = la_data_in[89] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58] = la_data_in[88] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59] = la_data_in[87] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60] = la_data_in[86] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61] = la_data_in[85] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62] = la_data_out[84] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63] = la_data_out[83] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64] = la_data_out[82] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65] = la_data_out[81] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66] = la_data_out[80] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67] = la_data_out[79] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68] = la_data_out[78] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69] = la_data_out[77] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70] = la_data_out[76] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71] = la_data_out[75] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72] = la_data_out[74] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73] = la_data_out[73] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74] = la_data_out[72] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75] = la_data_out[71] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76] = la_data_out[70] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77] = la_data_out[69] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78] = la_data_out[68] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79] = la_data_out[67] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80] = la_data_out[66] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81] = la_data_out[65] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82] = la_data_out[64] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83] = la_data_out[63] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84] = la_data_out[62] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85] = la_data_out[61] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86] = la_data_out[60] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87] = la_data_out[59] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88] = la_data_out[58] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89] = la_data_out[57] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90] = la_data_out[56] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91] = la_data_out[55] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92] = la_data_out[54] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93] = la_data_out[53] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94] = la_data_out[52] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95] = la_data_out[51] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[96] = la_data_out[50] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[97] = la_data_out[49] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[98] = la_data_out[48] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[99] = la_data_out[47] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[100] = la_data_out[46] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[101] = la_data_out[45] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[102] = la_data_out[44] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[103] = la_data_out[43] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[104] = la_data_out[42] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[105] = la_data_out[41] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[106] = la_data_out[40] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[107] = la_data_out[39] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[108] = la_data_out[38] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[109] = la_data_out[37] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[110] = la_data_out[36] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[111] = la_data_out[35] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[112] = la_data_out[34] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[113] = la_data_out[33] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[114] = la_data_out[32] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[115] = la_data_out[31] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[116] = la_data_out[30] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[117] = la_data_out[29] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[118] = la_data_out[28] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[119] = la_data_out[27] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[120] = la_data_out[26] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[121] = la_data_out[25] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[122] = la_data_out[24] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[123] = la_data_out[23] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[124] = la_data_out[22] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[125] = la_data_out[21] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[126] = la_data_out[20] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[127] = la_data_out[19] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[128] = la_data_out[18] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[129] = la_data_out[17] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[130] = la_data_out[16] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[131] = la_data_out[15] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[132] = la_data_out[14] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[133] = la_data_in[13] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[134] = la_data_out[12] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[135] = la_data_out[11] ;
assign prog_clk = io_in[37] ;
assign clk = io_in[36] ;
assign ccff_tail = io_out[35] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[136] = io_in[34] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[136] = io_out[34] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[136] = io_oeb[34] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[137] = io_in[33] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[137] = io_out[33] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[137] = io_oeb[33] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[138] = io_in[32] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[138] = io_out[32] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[138] = io_oeb[32] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[139] = io_in[31] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[139] = io_out[31] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[139] = io_oeb[31] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[140] = io_in[30] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[140] = io_out[30] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[140] = io_oeb[30] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[141] = io_in[29] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[141] = io_out[29] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[141] = io_oeb[29] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[142] = io_in[28] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[142] = io_out[28] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[142] = io_oeb[28] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[143] = io_in[27] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[143] = io_out[27] ;
assign gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[143] = io_oeb[27] ;
assign sc_head = io_in[26] ;
assign wb_la_switch = io_in[25] ;

sky130_fd_sc_hd__inv_8 WB_LA_SWITCH_INV ( .A ( io_in[25] ) , 
    .Y ( wb_la_switch_b ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_30_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[0] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_30_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[116] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_31_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[1] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_31_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[115] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_32_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[2] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_32_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[114] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_33_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[3] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_33_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[113] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_34_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[4] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_34_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[112] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_35_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[5] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_35_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[111] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_36_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[6] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_36_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[110] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_37_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[7] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_37_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[109] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_38_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[8] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_38_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[108] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_39_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[9] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_39_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[107] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_40_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[10] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_40_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[106] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_41_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[11] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_41_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[105] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_42_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[12] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_42_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[104] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_43_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[13] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_43_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[103] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_44_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[14] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_44_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[102] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_45_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[15] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_45_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[101] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_46_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[16] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_46_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[100] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_47_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[17] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_47_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[99] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_48_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[18] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_48_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[98] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_49_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[19] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_49_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[97] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_50_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[20] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_50_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[96] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_51_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[21] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_51_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[95] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_52_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[22] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_52_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[94] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_53_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[23] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_53_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[93] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_54_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[24] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_54_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[92] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_55_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[25] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_55_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[91] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_56_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[26] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_56_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[90] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_57_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[27] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_57_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[89] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_58_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[28] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_58_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[88] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_59_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[29] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_59_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[87] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_60_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[30] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_60_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[86] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_61_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_dat_o[31] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_61_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[85] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_62_MUX ( .A0 ( la_data_in[84] ) , 
    .A1 ( wbs_dat_i[0] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_63_MUX ( .A0 ( la_data_in[83] ) , 
    .A1 ( wbs_dat_i[1] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_64_MUX ( .A0 ( la_data_in[82] ) , 
    .A1 ( wbs_dat_i[2] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_65_MUX ( .A0 ( la_data_in[81] ) , 
    .A1 ( wbs_dat_i[3] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_66_MUX ( .A0 ( la_data_in[80] ) , 
    .A1 ( wbs_dat_i[4] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_67_MUX ( .A0 ( la_data_in[79] ) , 
    .A1 ( wbs_dat_i[5] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_68_MUX ( .A0 ( la_data_in[78] ) , 
    .A1 ( wbs_dat_i[6] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_69_MUX ( .A0 ( la_data_in[77] ) , 
    .A1 ( wbs_dat_i[7] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_70_MUX ( .A0 ( la_data_in[76] ) , 
    .A1 ( wbs_dat_i[8] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_71_MUX ( .A0 ( la_data_in[75] ) , 
    .A1 ( wbs_dat_i[9] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_72_MUX ( .A0 ( la_data_in[74] ) , 
    .A1 ( wbs_dat_i[10] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_73_MUX ( .A0 ( la_data_in[73] ) , 
    .A1 ( wbs_dat_i[11] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_74_MUX ( .A0 ( la_data_in[72] ) , 
    .A1 ( wbs_dat_i[12] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_75_MUX ( .A0 ( la_data_in[71] ) , 
    .A1 ( wbs_dat_i[13] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_76_MUX ( .A0 ( la_data_in[70] ) , 
    .A1 ( wbs_dat_i[14] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_77_MUX ( .A0 ( la_data_in[69] ) , 
    .A1 ( wbs_dat_i[15] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_78_MUX ( .A0 ( la_data_in[68] ) , 
    .A1 ( wbs_dat_i[16] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_79_MUX ( .A0 ( la_data_in[67] ) , 
    .A1 ( wbs_dat_i[17] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_80_MUX ( .A0 ( la_data_in[66] ) , 
    .A1 ( wbs_dat_i[18] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_81_MUX ( .A0 ( la_data_in[65] ) , 
    .A1 ( wbs_dat_i[19] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_82_MUX ( .A0 ( la_data_in[64] ) , 
    .A1 ( wbs_dat_i[20] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_83_MUX ( .A0 ( la_data_in[63] ) , 
    .A1 ( wbs_dat_i[21] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_84_MUX ( .A0 ( la_data_in[62] ) , 
    .A1 ( wbs_dat_i[22] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_85_MUX ( .A0 ( la_data_in[61] ) , 
    .A1 ( wbs_dat_i[23] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_86_MUX ( .A0 ( la_data_in[60] ) , 
    .A1 ( wbs_dat_i[24] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_87_MUX ( .A0 ( la_data_in[59] ) , 
    .A1 ( wbs_dat_i[25] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_88_MUX ( .A0 ( la_data_in[58] ) , 
    .A1 ( wbs_dat_i[26] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_89_MUX ( .A0 ( la_data_in[57] ) , 
    .A1 ( wbs_dat_i[27] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_90_MUX ( .A0 ( la_data_in[56] ) , 
    .A1 ( wbs_dat_i[28] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_91_MUX ( .A0 ( la_data_in[55] ) , 
    .A1 ( wbs_dat_i[29] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_92_MUX ( .A0 ( la_data_in[54] ) , 
    .A1 ( wbs_dat_i[30] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_93_MUX ( .A0 ( la_data_in[53] ) , 
    .A1 ( wbs_dat_i[31] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_94_MUX ( .A0 ( la_data_in[52] ) , 
    .A1 ( wbs_adr_i[0] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_95_MUX ( .A0 ( la_data_in[51] ) , 
    .A1 ( wbs_adr_i[1] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_96_MUX ( .A0 ( la_data_in[50] ) , 
    .A1 ( wbs_adr_i[2] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[96] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_97_MUX ( .A0 ( la_data_in[49] ) , 
    .A1 ( wbs_adr_i[3] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[97] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_98_MUX ( .A0 ( la_data_in[48] ) , 
    .A1 ( wbs_adr_i[4] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[98] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_99_MUX ( .A0 ( la_data_in[47] ) , 
    .A1 ( wbs_adr_i[5] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[99] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_100_MUX ( .A0 ( la_data_in[46] ) , 
    .A1 ( wbs_adr_i[6] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[100] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_101_MUX ( .A0 ( la_data_in[45] ) , 
    .A1 ( wbs_adr_i[7] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[101] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_102_MUX ( .A0 ( la_data_in[44] ) , 
    .A1 ( wbs_adr_i[8] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[102] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_103_MUX ( .A0 ( la_data_in[43] ) , 
    .A1 ( wbs_adr_i[9] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[103] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_104_MUX ( .A0 ( la_data_in[42] ) , 
    .A1 ( wbs_adr_i[10] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[104] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_105_MUX ( .A0 ( la_data_in[41] ) , 
    .A1 ( wbs_adr_i[11] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[105] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_106_MUX ( .A0 ( la_data_in[40] ) , 
    .A1 ( wbs_adr_i[12] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[106] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_107_MUX ( .A0 ( la_data_in[39] ) , 
    .A1 ( wbs_adr_i[13] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[107] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_108_MUX ( .A0 ( la_data_in[38] ) , 
    .A1 ( wbs_adr_i[14] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[108] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_109_MUX ( .A0 ( la_data_in[37] ) , 
    .A1 ( wbs_adr_i[15] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[109] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_110_MUX ( .A0 ( la_data_in[36] ) , 
    .A1 ( wbs_adr_i[16] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[110] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_111_MUX ( .A0 ( la_data_in[35] ) , 
    .A1 ( wbs_adr_i[17] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[111] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_112_MUX ( .A0 ( la_data_in[34] ) , 
    .A1 ( wbs_adr_i[18] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[112] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_113_MUX ( .A0 ( la_data_in[33] ) , 
    .A1 ( wbs_adr_i[19] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[113] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_114_MUX ( .A0 ( la_data_in[32] ) , 
    .A1 ( wbs_adr_i[20] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[114] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_115_MUX ( .A0 ( la_data_in[31] ) , 
    .A1 ( wbs_adr_i[21] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[115] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_116_MUX ( .A0 ( la_data_in[30] ) , 
    .A1 ( wbs_adr_i[22] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[116] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_117_MUX ( .A0 ( la_data_in[29] ) , 
    .A1 ( wbs_adr_i[23] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[117] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_118_MUX ( .A0 ( la_data_in[28] ) , 
    .A1 ( wbs_adr_i[24] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[118] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_119_MUX ( .A0 ( la_data_in[27] ) , 
    .A1 ( wbs_adr_i[25] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[119] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_120_MUX ( .A0 ( la_data_in[26] ) , 
    .A1 ( wbs_adr_i[26] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[120] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_121_MUX ( .A0 ( la_data_in[25] ) , 
    .A1 ( wbs_adr_i[27] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[121] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_122_MUX ( .A0 ( la_data_in[24] ) , 
    .A1 ( wbs_adr_i[28] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[122] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_123_MUX ( .A0 ( la_data_in[23] ) , 
    .A1 ( wbs_adr_i[29] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[123] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_124_MUX ( .A0 ( la_data_in[22] ) , 
    .A1 ( wbs_adr_i[30] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[124] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_125_MUX ( .A0 ( la_data_in[21] ) , 
    .A1 ( wbs_adr_i[31] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[125] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_126_MUX ( .A0 ( la_data_in[20] ) , 
    .A1 ( wbs_sel_i[0] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[126] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_127_MUX ( .A0 ( la_data_in[19] ) , 
    .A1 ( wbs_sel_i[1] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[127] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_128_MUX ( .A0 ( la_data_in[18] ) , 
    .A1 ( wbs_sel_i[2] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[128] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_129_MUX ( .A0 ( la_data_in[17] ) , 
    .A1 ( wbs_sel_i[3] ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[129] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_130_MUX ( .A0 ( la_data_in[16] ) , 
    .A1 ( wbs_we_i ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[130] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_131_MUX ( .A0 ( la_data_in[15] ) , 
    .A1 ( wbs_stb_i ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[131] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_132_MUX ( .A0 ( la_data_in[14] ) , 
    .A1 ( wbs_cyc_i ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[132] ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_133_DEMUX_WB ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[133] ) , .TE_B ( wb_la_switch_b ) , 
    .Z ( wbs_ack_o ) ) ;
sky130_fd_sc_hd__ebufn_4 FPGA2SOC_OUT_133_DEMUX_LA ( 
    .A ( gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[133] ) , .TE_B ( io_in[25] ) , 
    .Z ( la_data_out[13] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_134_MUX ( .A0 ( la_data_in[12] ) , 
    .A1 ( wb_rst_i ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[134] ) ) ;
sky130_fd_sc_hd__mux2_1 FPGA2SOC_IN_135_MUX ( .A0 ( la_data_in[11] ) , 
    .A1 ( wb_clk_i ) , .S ( io_in[25] ) , 
    .X ( gfpga_pad_EMBEDDED_IO_HD_SOC_IN[135] ) ) ;
fpga_core fpga_core_uut ( .pReset ( io_in[3] ) , .prog_clk ( io_in[37] ) , 
    .Test_en ( io_in[0] ) , .IO_ISOL_N ( io_in[1] ) , .clk ( io_in[36] ) , 
    .Reset ( io_in[2] ) ,
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN ( { io_in[24] , io_in[23] , io_in[22] , 
        io_in[21] , io_in[20] , io_in[19] , io_in[18] , io_in[17] , 
        io_in[16] , io_in[15] , io_in[14] , io_in[13] , io_in[10] , io_in[9] , 
        io_in[8] , io_in[7] , io_in[6] , io_in[5] , io_in[4] , 
        la_data_in[127] , la_data_in[126] , la_data_in[125] , 
        la_data_in[124] , la_data_in[123] , la_data_in[122] , 
        la_data_in[121] , la_data_in[120] , la_data_in[119] , 
        la_data_in[118] , la_data_in[117] , la_data_in[116] , 
        la_data_in[115] , la_data_in[114] , la_data_in[113] , 
        la_data_in[112] , la_data_in[111] , la_data_in[110] , 
        la_data_in[109] , la_data_in[108] , la_data_in[107] , 
        la_data_in[106] , la_data_in[105] , la_data_in[104] , 
        la_data_in[103] , la_data_in[102] , la_data_in[101] , 
        la_data_in[100] , la_data_in[99] , la_data_in[98] , la_data_in[97] , 
        la_data_in[96] , la_data_in[95] , la_data_in[94] , la_data_in[93] , 
        la_data_in[92] , la_data_in[91] , la_data_in[90] , la_data_in[89] , 
        la_data_in[88] , la_data_in[87] , la_data_in[86] , la_data_in[85] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[96] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[97] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[98] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[99] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[100] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[101] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[102] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[103] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[104] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[105] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[106] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[107] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[108] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[109] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[110] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[111] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[112] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[113] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[114] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[115] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[116] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[117] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[118] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[119] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[120] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[121] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[122] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[123] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[124] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[125] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[126] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[127] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[128] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[129] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[130] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[131] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[132] , la_data_in[13] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[134] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_IN[135] , io_in[34] , io_in[33] , 
        io_in[32] , io_in[31] , io_in[30] , io_in[29] , io_in[28] , 
        io_in[27] } ) ,
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT ( { io_out[24] , io_out[23] , 
        io_out[22] , io_out[21] , io_out[20] , io_out[19] , io_out[18] , 
        io_out[17] , io_out[16] , io_out[15] , io_out[14] , io_out[13] , 
        io_out[10] , io_out[9] , io_out[8] , io_out[7] , io_out[6] , 
        io_out[5] , io_out[4] , la_data_out[127] , la_data_out[126] , 
        la_data_out[125] , la_data_out[124] , la_data_out[123] , 
        la_data_out[122] , la_data_out[121] , la_data_out[120] , 
        la_data_out[119] , la_data_out[118] , la_data_out[117] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61] , la_data_out[84] , 
        la_data_out[83] , la_data_out[82] , la_data_out[81] , 
        la_data_out[80] , la_data_out[79] , la_data_out[78] , 
        la_data_out[77] , la_data_out[76] , la_data_out[75] , 
        la_data_out[74] , la_data_out[73] , la_data_out[72] , 
        la_data_out[71] , la_data_out[70] , la_data_out[69] , 
        la_data_out[68] , la_data_out[67] , la_data_out[66] , 
        la_data_out[65] , la_data_out[64] , la_data_out[63] , 
        la_data_out[62] , la_data_out[61] , la_data_out[60] , 
        la_data_out[59] , la_data_out[58] , la_data_out[57] , 
        la_data_out[56] , la_data_out[55] , la_data_out[54] , 
        la_data_out[53] , la_data_out[52] , la_data_out[51] , 
        la_data_out[50] , la_data_out[49] , la_data_out[48] , 
        la_data_out[47] , la_data_out[46] , la_data_out[45] , 
        la_data_out[44] , la_data_out[43] , la_data_out[42] , 
        la_data_out[41] , la_data_out[40] , la_data_out[39] , 
        la_data_out[38] , la_data_out[37] , la_data_out[36] , 
        la_data_out[35] , la_data_out[34] , la_data_out[33] , 
        la_data_out[32] , la_data_out[31] , la_data_out[30] , 
        la_data_out[29] , la_data_out[28] , la_data_out[27] , 
        la_data_out[26] , la_data_out[25] , la_data_out[24] , 
        la_data_out[23] , la_data_out[22] , la_data_out[21] , 
        la_data_out[20] , la_data_out[19] , la_data_out[18] , 
        la_data_out[17] , la_data_out[16] , la_data_out[15] , 
        la_data_out[14] , gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[133] , 
        la_data_out[12] , la_data_out[11] , io_out[34] , io_out[33] , 
        io_out[32] , io_out[31] , io_out[30] , io_out[29] , io_out[28] , 
        io_out[27] } ) ,
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR ( { io_oeb[24] , io_oeb[23] , 
        io_oeb[22] , io_oeb[21] , io_oeb[20] , io_oeb[19] , io_oeb[18] , 
        io_oeb[17] , io_oeb[16] , io_oeb[15] , io_oeb[14] , io_oeb[13] , 
        io_oeb[10] , io_oeb[9] , io_oeb[8] , io_oeb[7] , io_oeb[6] , 
        io_oeb[5] , io_oeb[4] , gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[96] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[97] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[98] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[99] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[100] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[101] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[102] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[103] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[104] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[105] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[106] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[107] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[108] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[109] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[110] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[111] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[112] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[113] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[114] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[115] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[116] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[117] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[118] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[119] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[120] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[121] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[122] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[123] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[124] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[125] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[126] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[127] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[128] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[129] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[130] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[131] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[132] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[133] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[134] , 
        gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[135] , io_oeb[34] , io_oeb[33] , 
        io_oeb[32] , io_oeb[31] , io_oeb[30] , io_oeb[29] , io_oeb[28] , 
        io_oeb[27] } ) ,
    .ccff_head ( io_in[12] ) , .ccff_tail ( io_out[35] ) , 
    .sc_head ( io_in[26] ) , .sc_tail ( io_out[11] ) , 
    .h_incr0 ( SYNOPSYS_UNCONNECTED_1 ) , .p0 ( optlc_net_20 ) , 
    .p1 ( optlc_net_21 ) , .p2 ( optlc_net_22 ) , .p3 ( optlc_net_23 ) , 
    .p4 ( optlc_net_24 ) , .p5 ( optlc_net_25 ) , .p6 ( optlc_net_26 ) , 
    .p7 ( optlc_net_27 ) , .p8 ( optlc_net_28 ) , .p9 ( optlc_net_29 ) , 
    .p10 ( optlc_net_30 ) , .p11 ( optlc_net_31 ) , .p12 ( optlc_net_32 ) , 
    .p13 ( optlc_net_33 ) , .p14 ( optlc_net_34 ) , .p15 ( optlc_net_35 ) , 
    .p16 ( optlc_net_36 ) , .p17 ( optlc_net_37 ) , .p18 ( optlc_net_38 ) , 
    .p19 ( optlc_net_39 ) , .p20 ( optlc_net_40 ) , .p21 ( optlc_net_41 ) , 
    .p22 ( optlc_net_42 ) , .p23 ( optlc_net_43 ) , .p24 ( optlc_net_44 ) , 
    .p25 ( optlc_net_45 ) , .p26 ( optlc_net_46 ) , .p27 ( optlc_net_47 ) , 
    .p28 ( optlc_net_48 ) , .p29 ( optlc_net_49 ) , .p30 ( optlc_net_50 ) , 
    .p31 ( optlc_net_51 ) , .p32 ( optlc_net_52 ) , .p33 ( optlc_net_53 ) , 
    .p34 ( optlc_net_54 ) , .p35 ( optlc_net_55 ) , .p36 ( optlc_net_56 ) , 
    .p37 ( optlc_net_57 ) , .p38 ( optlc_net_58 ) , .p39 ( optlc_net_59 ) , 
    .p40 ( optlc_net_60 ) , .p41 ( optlc_net_61 ) , .p42 ( optlc_net_62 ) , 
    .p43 ( optlc_net_63 ) , .p44 ( optlc_net_64 ) , .p45 ( optlc_net_65 ) , 
    .p46 ( optlc_net_66 ) , .p47 ( optlc_net_67 ) , .p48 ( optlc_net_68 ) , 
    .p49 ( optlc_net_69 ) , .p50 ( optlc_net_70 ) , .p51 ( optlc_net_71 ) , 
    .p52 ( optlc_net_72 ) , .p53 ( optlc_net_73 ) , .p54 ( optlc_net_74 ) , 
    .p55 ( optlc_net_75 ) , .p56 ( optlc_net_76 ) , .p57 ( optlc_net_77 ) , 
    .p58 ( optlc_net_78 ) , .p59 ( optlc_net_79 ) , .p60 ( optlc_net_80 ) , 
    .p61 ( optlc_net_81 ) , .p62 ( optlc_net_82 ) , .p63 ( optlc_net_83 ) , 
    .p64 ( optlc_net_84 ) , .p65 ( optlc_net_85 ) , .p66 ( optlc_net_86 ) , 
    .p67 ( optlc_net_87 ) , .p68 ( optlc_net_88 ) , .p69 ( optlc_net_89 ) , 
    .p70 ( optlc_net_90 ) , .p71 ( optlc_net_91 ) , .p72 ( optlc_net_92 ) , 
    .p73 ( optlc_net_93 ) , .p74 ( optlc_net_94 ) , .p75 ( optlc_net_95 ) , 
    .p76 ( optlc_net_96 ) , .p77 ( optlc_net_97 ) , .p78 ( optlc_net_98 ) , 
    .p79 ( optlc_net_99 ) , .p80 ( optlc_net_100 ) , .p81 ( optlc_net_101 ) , 
    .p82 ( optlc_net_102 ) , .p83 ( optlc_net_103 ) , .p84 ( optlc_net_104 ) , 
    .p85 ( optlc_net_105 ) , .p86 ( optlc_net_106 ) , .p87 ( optlc_net_107 ) , 
    .p88 ( optlc_net_108 ) , .p89 ( optlc_net_109 ) , .p90 ( optlc_net_110 ) , 
    .p91 ( optlc_net_111 ) , .p92 ( optlc_net_112 ) , .p93 ( optlc_net_113 ) , 
    .p94 ( optlc_net_114 ) , .p95 ( optlc_net_115 ) , .p96 ( optlc_net_116 ) , 
    .p97 ( optlc_net_117 ) , .p98 ( optlc_net_118 ) , .p99 ( optlc_net_119 ) , 
    .p100 ( optlc_net_120 ) , .p101 ( optlc_net_121 ) , 
    .p102 ( optlc_net_122 ) , .p103 ( optlc_net_123 ) , 
    .p104 ( optlc_net_124 ) , .p105 ( optlc_net_125 ) , 
    .p106 ( optlc_net_126 ) , .p107 ( optlc_net_127 ) , 
    .p108 ( optlc_net_128 ) , .p109 ( optlc_net_129 ) , 
    .p110 ( optlc_net_130 ) , .p111 ( optlc_net_131 ) , 
    .p112 ( optlc_net_132 ) , .p113 ( optlc_net_133 ) , 
    .p114 ( optlc_net_134 ) , .p115 ( optlc_net_135 ) , 
    .p116 ( optlc_net_136 ) , .p117 ( optlc_net_137 ) , 
    .p118 ( optlc_net_138 ) , .p119 ( optlc_net_139 ) , 
    .p120 ( optlc_net_140 ) , .p121 ( optlc_net_141 ) , 
    .p122 ( optlc_net_142 ) , .p123 ( optlc_net_143 ) , 
    .p124 ( optlc_net_144 ) , .p125 ( optlc_net_145 ) , 
    .p126 ( optlc_net_146 ) , .p127 ( optlc_net_147 ) , 
    .p128 ( optlc_net_148 ) , .p129 ( optlc_net_149 ) , 
    .p130 ( optlc_net_150 ) , .p131 ( optlc_net_151 ) , 
    .p132 ( optlc_net_152 ) , .p133 ( optlc_net_153 ) , 
    .p134 ( optlc_net_154 ) , .p135 ( optlc_net_155 ) , 
    .p136 ( optlc_net_156 ) , .p137 ( optlc_net_157 ) , 
    .p138 ( optlc_net_158 ) , .p139 ( optlc_net_159 ) , 
    .p140 ( optlc_net_160 ) , .p141 ( optlc_net_161 ) , 
    .p142 ( optlc_net_162 ) , .p143 ( optlc_net_163 ) , 
    .p144 ( optlc_net_164 ) , .p145 ( optlc_net_165 ) , 
    .p146 ( optlc_net_166 ) , .p147 ( optlc_net_167 ) , 
    .p148 ( optlc_net_168 ) , .p149 ( optlc_net_169 ) , 
    .p150 ( optlc_net_170 ) , .p151 ( optlc_net_171 ) , 
    .p152 ( optlc_net_172 ) , .p153 ( optlc_net_173 ) , 
    .p154 ( optlc_net_174 ) , .p155 ( optlc_net_175 ) , 
    .p156 ( optlc_net_176 ) , .p157 ( optlc_net_177 ) , 
    .p158 ( optlc_net_178 ) , .p159 ( optlc_net_179 ) , 
    .p160 ( optlc_net_180 ) , .p161 ( optlc_net_181 ) , 
    .p162 ( optlc_net_182 ) , .p163 ( optlc_net_183 ) , 
    .p164 ( optlc_net_184 ) , .p165 ( optlc_net_185 ) , 
    .p166 ( optlc_net_186 ) , .p167 ( optlc_net_187 ) , 
    .p168 ( optlc_net_188 ) , .p169 ( optlc_net_189 ) , 
    .p170 ( optlc_net_190 ) , .p171 ( optlc_net_191 ) , 
    .p172 ( optlc_net_192 ) , .p173 ( optlc_net_193 ) , 
    .p174 ( optlc_net_194 ) , .p175 ( optlc_net_195 ) , 
    .p176 ( optlc_net_196 ) , .p177 ( optlc_net_197 ) , 
    .p178 ( optlc_net_198 ) , .p179 ( optlc_net_199 ) , 
    .p180 ( optlc_net_200 ) , .p181 ( optlc_net_201 ) , 
    .p182 ( optlc_net_202 ) , .p183 ( optlc_net_203 ) , 
    .p184 ( optlc_net_204 ) , .p185 ( optlc_net_205 ) , 
    .p186 ( optlc_net_206 ) , .p187 ( optlc_net_207 ) , 
    .p188 ( optlc_net_208 ) , .p189 ( optlc_net_209 ) , 
    .p190 ( optlc_net_210 ) , .p191 ( optlc_net_211 ) , 
    .p192 ( optlc_net_212 ) , .p193 ( optlc_net_213 ) , 
    .p194 ( optlc_net_214 ) , .p195 ( optlc_net_215 ) , 
    .p196 ( optlc_net_216 ) , .p197 ( optlc_net_217 ) , 
    .p198 ( optlc_net_218 ) , .p199 ( optlc_net_219 ) , 
    .p200 ( optlc_net_220 ) , .p201 ( optlc_net_221 ) , 
    .p202 ( optlc_net_222 ) , .p203 ( optlc_net_223 ) , 
    .p204 ( optlc_net_224 ) , .p205 ( optlc_net_225 ) , 
    .p206 ( optlc_net_226 ) , .p207 ( optlc_net_227 ) , 
    .p208 ( optlc_net_228 ) , .p209 ( optlc_net_229 ) , 
    .p210 ( optlc_net_230 ) , .p211 ( optlc_net_231 ) , 
    .p212 ( optlc_net_232 ) , .p213 ( optlc_net_233 ) , 
    .p214 ( optlc_net_234 ) , .p215 ( optlc_net_235 ) , 
    .p216 ( optlc_net_236 ) , .p217 ( optlc_net_237 ) , 
    .p218 ( optlc_net_238 ) , .p219 ( optlc_net_239 ) , 
    .p220 ( optlc_net_240 ) , .p221 ( optlc_net_241 ) , 
    .p222 ( optlc_net_242 ) , .p223 ( optlc_net_243 ) , 
    .p224 ( optlc_net_244 ) , .p225 ( optlc_net_245 ) , 
    .p226 ( optlc_net_246 ) , .p227 ( optlc_net_247 ) , 
    .p228 ( optlc_net_248 ) , .p229 ( optlc_net_249 ) , 
    .p230 ( optlc_net_250 ) , .p231 ( optlc_net_251 ) , 
    .p232 ( optlc_net_252 ) , .p233 ( optlc_net_253 ) , 
    .p234 ( optlc_net_254 ) , .p235 ( optlc_net_255 ) , 
    .p236 ( optlc_net_256 ) , .p237 ( optlc_net_257 ) , 
    .p238 ( optlc_net_258 ) , .p239 ( optlc_net_259 ) , 
    .p240 ( optlc_net_260 ) , .p241 ( optlc_net_261 ) , 
    .p242 ( optlc_net_262 ) , .p243 ( optlc_net_263 ) , 
    .p244 ( optlc_net_264 ) , .p245 ( optlc_net_265 ) , 
    .p246 ( optlc_net_266 ) , .p247 ( optlc_net_267 ) , 
    .p248 ( optlc_net_268 ) , .p249 ( optlc_net_269 ) , 
    .p250 ( optlc_net_270 ) , .p251 ( optlc_net_271 ) , 
    .p252 ( optlc_net_272 ) , .p253 ( optlc_net_273 ) , 
    .p254 ( optlc_net_274 ) , .p255 ( optlc_net_275 ) , 
    .p256 ( optlc_net_276 ) , .p257 ( optlc_net_277 ) , 
    .p258 ( optlc_net_278 ) , .p259 ( optlc_net_279 ) , 
    .p260 ( optlc_net_280 ) , .p261 ( optlc_net_281 ) , 
    .p262 ( optlc_net_282 ) , .p263 ( optlc_net_283 ) , 
    .p264 ( optlc_net_284 ) , .p265 ( optlc_net_285 ) , 
    .p266 ( optlc_net_286 ) , .p267 ( optlc_net_287 ) , 
    .p268 ( optlc_net_288 ) , .p269 ( optlc_net_289 ) , 
    .p270 ( optlc_net_290 ) , .p271 ( optlc_net_291 ) , 
    .p272 ( optlc_net_292 ) , .p273 ( optlc_net_293 ) , 
    .p274 ( optlc_net_294 ) , .p275 ( optlc_net_295 ) , 
    .p276 ( optlc_net_296 ) , .p277 ( optlc_net_297 ) , 
    .p278 ( optlc_net_298 ) , .p279 ( optlc_net_299 ) , 
    .p280 ( optlc_net_300 ) , .p281 ( optlc_net_301 ) , 
    .p282 ( optlc_net_302 ) , .p283 ( optlc_net_303 ) , 
    .p284 ( optlc_net_304 ) , .p285 ( optlc_net_305 ) , 
    .p286 ( optlc_net_306 ) , .p287 ( optlc_net_307 ) , 
    .p288 ( optlc_net_308 ) , .p289 ( optlc_net_309 ) , 
    .p290 ( optlc_net_310 ) , .p291 ( optlc_net_311 ) , 
    .p292 ( optlc_net_312 ) , .p293 ( optlc_net_313 ) , 
    .p294 ( optlc_net_314 ) , .p295 ( optlc_net_315 ) , 
    .p296 ( optlc_net_316 ) , .p297 ( optlc_net_317 ) , 
    .p298 ( optlc_net_318 ) , .p299 ( optlc_net_319 ) , 
    .p300 ( optlc_net_320 ) , .p301 ( optlc_net_321 ) , 
    .p302 ( optlc_net_322 ) , .p303 ( optlc_net_323 ) , 
    .p304 ( optlc_net_324 ) , .p305 ( optlc_net_325 ) , 
    .p306 ( optlc_net_326 ) , .p307 ( optlc_net_327 ) , 
    .p308 ( optlc_net_328 ) , .p309 ( optlc_net_329 ) , 
    .p310 ( optlc_net_330 ) , .p311 ( optlc_net_331 ) , 
    .p312 ( optlc_net_332 ) , .p313 ( optlc_net_333 ) , 
    .p314 ( optlc_net_334 ) , .p315 ( optlc_net_335 ) , 
    .p316 ( optlc_net_336 ) , .p317 ( optlc_net_337 ) , 
    .p318 ( optlc_net_338 ) , .p319 ( optlc_net_339 ) , 
    .p320 ( optlc_net_340 ) , .p321 ( optlc_net_341 ) , 
    .p322 ( optlc_net_342 ) , .p323 ( optlc_net_343 ) , 
    .p324 ( optlc_net_344 ) , .p325 ( optlc_net_345 ) , 
    .p326 ( optlc_net_346 ) , .p327 ( optlc_net_347 ) , 
    .p328 ( optlc_net_348 ) , .p329 ( optlc_net_349 ) , 
    .p330 ( optlc_net_350 ) , .p331 ( optlc_net_351 ) , 
    .p332 ( optlc_net_352 ) , .p333 ( optlc_net_353 ) , 
    .p334 ( optlc_net_354 ) , .p335 ( optlc_net_355 ) , 
    .p336 ( optlc_net_356 ) , .p337 ( optlc_net_357 ) , 
    .p338 ( optlc_net_358 ) , .p339 ( optlc_net_359 ) , 
    .p340 ( optlc_net_360 ) , .p341 ( optlc_net_361 ) , 
    .p342 ( optlc_net_362 ) , .p343 ( optlc_net_363 ) , 
    .p344 ( optlc_net_364 ) , .p345 ( optlc_net_365 ) , 
    .p346 ( optlc_net_366 ) , .p347 ( optlc_net_367 ) , 
    .p348 ( optlc_net_368 ) , .p349 ( optlc_net_369 ) , 
    .p350 ( optlc_net_370 ) , .p351 ( optlc_net_371 ) , 
    .p352 ( optlc_net_372 ) , .p353 ( optlc_net_373 ) , 
    .p354 ( optlc_net_374 ) , .p355 ( optlc_net_375 ) , 
    .p356 ( optlc_net_376 ) , .p357 ( optlc_net_377 ) , 
    .p358 ( optlc_net_378 ) , .p359 ( optlc_net_379 ) , 
    .p360 ( optlc_net_380 ) , .p361 ( optlc_net_381 ) , 
    .p362 ( optlc_net_382 ) , .p363 ( optlc_net_383 ) , 
    .p364 ( optlc_net_384 ) , .p365 ( optlc_net_385 ) , 
    .p366 ( optlc_net_386 ) , .p367 ( optlc_net_387 ) , 
    .p368 ( optlc_net_388 ) , .p369 ( optlc_net_389 ) , 
    .p370 ( optlc_net_390 ) , .p371 ( optlc_net_391 ) , 
    .p372 ( optlc_net_392 ) , .p373 ( optlc_net_393 ) , 
    .p374 ( optlc_net_394 ) , .p375 ( optlc_net_395 ) , 
    .p376 ( optlc_net_396 ) , .p377 ( optlc_net_397 ) , 
    .p378 ( optlc_net_398 ) , .p379 ( optlc_net_399 ) , 
    .p380 ( optlc_net_400 ) , .p381 ( optlc_net_401 ) , 
    .p382 ( optlc_net_402 ) , .p383 ( optlc_net_403 ) , 
    .p384 ( optlc_net_404 ) , .p385 ( optlc_net_405 ) , 
    .p386 ( optlc_net_406 ) , .p387 ( optlc_net_407 ) , 
    .p388 ( optlc_net_408 ) , .p389 ( optlc_net_409 ) , 
    .p390 ( optlc_net_410 ) , .p391 ( optlc_net_411 ) , 
    .p392 ( optlc_net_412 ) , .p393 ( optlc_net_413 ) , 
    .p394 ( optlc_net_414 ) , .p395 ( optlc_net_415 ) , 
    .p396 ( optlc_net_416 ) , .p397 ( optlc_net_417 ) , 
    .p398 ( optlc_net_418 ) , .p399 ( optlc_net_419 ) , 
    .p400 ( optlc_net_420 ) , .p401 ( optlc_net_421 ) , 
    .p402 ( optlc_net_422 ) , .p403 ( optlc_net_423 ) , 
    .p404 ( optlc_net_424 ) , .p405 ( optlc_net_425 ) , 
    .p406 ( optlc_net_426 ) , .p407 ( optlc_net_427 ) , 
    .p408 ( optlc_net_428 ) , .p409 ( optlc_net_429 ) , 
    .p410 ( optlc_net_430 ) , .p411 ( optlc_net_431 ) , 
    .p412 ( optlc_net_432 ) , .p413 ( optlc_net_433 ) , 
    .p414 ( optlc_net_434 ) , .p415 ( optlc_net_435 ) , 
    .p416 ( optlc_net_436 ) , .p417 ( optlc_net_437 ) , 
    .p418 ( optlc_net_438 ) , .p419 ( optlc_net_439 ) , 
    .p420 ( optlc_net_440 ) , .p421 ( optlc_net_441 ) , 
    .p422 ( optlc_net_442 ) , .p423 ( optlc_net_443 ) , 
    .p424 ( optlc_net_444 ) , .p425 ( optlc_net_445 ) , 
    .p426 ( optlc_net_446 ) , .p427 ( optlc_net_447 ) , 
    .p428 ( optlc_net_448 ) , .p429 ( optlc_net_449 ) , 
    .p430 ( optlc_net_450 ) , .p431 ( optlc_net_451 ) , 
    .p432 ( optlc_net_452 ) , .p433 ( optlc_net_453 ) , 
    .p434 ( optlc_net_454 ) , .p435 ( optlc_net_455 ) , 
    .p436 ( optlc_net_456 ) , .p437 ( optlc_net_457 ) , 
    .p438 ( optlc_net_458 ) , .p439 ( optlc_net_459 ) , 
    .p440 ( optlc_net_460 ) , .p441 ( optlc_net_461 ) , 
    .p442 ( optlc_net_462 ) , .p443 ( optlc_net_463 ) , 
    .p444 ( optlc_net_464 ) , .p445 ( optlc_net_465 ) , 
    .p446 ( optlc_net_466 ) , .p447 ( optlc_net_467 ) , 
    .p448 ( optlc_net_468 ) , .p449 ( optlc_net_469 ) , 
    .p450 ( optlc_net_470 ) , .p451 ( optlc_net_471 ) , 
    .p452 ( optlc_net_472 ) , .p453 ( optlc_net_473 ) , 
    .p454 ( optlc_net_474 ) , .p455 ( optlc_net_475 ) , 
    .p456 ( optlc_net_476 ) , .p457 ( optlc_net_477 ) , 
    .p458 ( optlc_net_478 ) , .p459 ( optlc_net_479 ) , 
    .p460 ( optlc_net_480 ) , .p461 ( optlc_net_481 ) , 
    .p462 ( optlc_net_482 ) , .p463 ( optlc_net_483 ) , 
    .p464 ( optlc_net_484 ) , .p465 ( optlc_net_485 ) , 
    .p466 ( optlc_net_486 ) , .p467 ( optlc_net_487 ) , 
    .p468 ( optlc_net_488 ) , .p469 ( optlc_net_489 ) , 
    .p470 ( optlc_net_490 ) , .p471 ( optlc_net_491 ) , 
    .p472 ( optlc_net_492 ) , .p473 ( optlc_net_493 ) , 
    .p474 ( optlc_net_494 ) , .p475 ( optlc_net_495 ) , 
    .p476 ( optlc_net_496 ) , .p477 ( optlc_net_497 ) , 
    .p478 ( optlc_net_498 ) , .p479 ( optlc_net_499 ) , 
    .p480 ( optlc_net_500 ) , .p481 ( optlc_net_501 ) , 
    .p482 ( optlc_net_502 ) , .p483 ( optlc_net_503 ) , 
    .p484 ( optlc_net_504 ) , .p485 ( optlc_net_505 ) , 
    .p486 ( optlc_net_506 ) , .p487 ( optlc_net_507 ) , 
    .p488 ( optlc_net_508 ) , .p489 ( optlc_net_509 ) , 
    .p490 ( optlc_net_510 ) , .p491 ( optlc_net_511 ) , 
    .p492 ( optlc_net_512 ) , .p493 ( optlc_net_513 ) , 
    .p494 ( optlc_net_514 ) , .p495 ( optlc_net_515 ) , 
    .p496 ( optlc_net_516 ) , .p497 ( optlc_net_517 ) , 
    .p498 ( optlc_net_518 ) , .p499 ( optlc_net_519 ) , 
    .p500 ( optlc_net_520 ) , .p501 ( optlc_net_521 ) , 
    .p502 ( optlc_net_522 ) , .p503 ( optlc_net_523 ) , 
    .p504 ( optlc_net_524 ) , .p505 ( optlc_net_525 ) , 
    .p506 ( optlc_net_526 ) , .p507 ( optlc_net_527 ) , 
    .p508 ( optlc_net_528 ) , .p509 ( optlc_net_529 ) , 
    .p510 ( optlc_net_530 ) , .p511 ( optlc_net_531 ) , 
    .p512 ( optlc_net_532 ) , .p513 ( optlc_net_533 ) , 
    .p514 ( optlc_net_534 ) , .p515 ( optlc_net_535 ) , 
    .p516 ( optlc_net_536 ) , .p517 ( optlc_net_537 ) , 
    .p518 ( optlc_net_538 ) , .p519 ( optlc_net_539 ) , 
    .p520 ( optlc_net_540 ) , .p521 ( optlc_net_541 ) , 
    .p522 ( optlc_net_542 ) , .p523 ( optlc_net_543 ) , 
    .p524 ( optlc_net_544 ) , .p525 ( optlc_net_545 ) , 
    .p526 ( optlc_net_546 ) , .p527 ( optlc_net_547 ) , 
    .p528 ( optlc_net_548 ) , .p529 ( optlc_net_549 ) , 
    .p530 ( optlc_net_550 ) , .p531 ( optlc_net_551 ) , 
    .p532 ( optlc_net_552 ) , .p533 ( optlc_net_553 ) , 
    .p534 ( optlc_net_554 ) , .p535 ( optlc_net_555 ) , 
    .p536 ( optlc_net_556 ) , .p537 ( optlc_net_557 ) , 
    .p538 ( optlc_net_558 ) , .p539 ( optlc_net_559 ) , 
    .p540 ( optlc_net_560 ) , .p541 ( optlc_net_561 ) , 
    .p542 ( optlc_net_562 ) , .p543 ( optlc_net_563 ) , 
    .p544 ( optlc_net_564 ) , .p545 ( optlc_net_565 ) , 
    .p546 ( optlc_net_566 ) , .p547 ( optlc_net_567 ) , 
    .p548 ( optlc_net_568 ) , .p549 ( optlc_net_569 ) , 
    .p550 ( optlc_net_570 ) , .p551 ( optlc_net_571 ) , 
    .p552 ( optlc_net_572 ) , .p553 ( optlc_net_573 ) , 
    .p554 ( optlc_net_574 ) , .p555 ( optlc_net_575 ) , 
    .p556 ( optlc_net_576 ) , .p557 ( optlc_net_577 ) , 
    .p558 ( optlc_net_578 ) , .p559 ( optlc_net_579 ) , 
    .p560 ( optlc_net_580 ) , .p561 ( optlc_net_581 ) , 
    .p562 ( optlc_net_582 ) , .p563 ( optlc_net_583 ) , 
    .p564 ( optlc_net_584 ) , .p565 ( optlc_net_585 ) , 
    .p566 ( optlc_net_586 ) , .p567 ( optlc_net_587 ) , 
    .p568 ( optlc_net_588 ) , .p569 ( optlc_net_589 ) , 
    .p570 ( optlc_net_590 ) , .p571 ( optlc_net_591 ) , 
    .p572 ( optlc_net_592 ) , .p573 ( optlc_net_593 ) , 
    .p574 ( optlc_net_594 ) , .p575 ( optlc_net_595 ) , 
    .p576 ( optlc_net_596 ) , .p577 ( optlc_net_597 ) , 
    .p578 ( optlc_net_598 ) , .p579 ( optlc_net_599 ) , 
    .p580 ( optlc_net_600 ) , .p581 ( optlc_net_601 ) , 
    .p582 ( optlc_net_602 ) , .p583 ( optlc_net_603 ) , 
    .p584 ( optlc_net_604 ) , .p585 ( optlc_net_605 ) , 
    .p586 ( optlc_net_606 ) , .p587 ( optlc_net_607 ) , 
    .p588 ( optlc_net_608 ) , .p589 ( optlc_net_609 ) , 
    .p590 ( optlc_net_610 ) , .p591 ( optlc_net_611 ) , 
    .p592 ( optlc_net_612 ) , .p593 ( optlc_net_613 ) , 
    .p594 ( optlc_net_614 ) , .p595 ( optlc_net_615 ) , 
    .p596 ( optlc_net_616 ) , .p597 ( optlc_net_617 ) , 
    .p598 ( optlc_net_618 ) , .p599 ( optlc_net_619 ) , 
    .p600 ( optlc_net_620 ) , .p601 ( optlc_net_621 ) , 
    .p602 ( optlc_net_622 ) , .p603 ( optlc_net_623 ) , 
    .p604 ( optlc_net_624 ) , .p605 ( optlc_net_625 ) , 
    .p606 ( optlc_net_626 ) , .p607 ( optlc_net_627 ) , 
    .p608 ( optlc_net_628 ) , .p609 ( optlc_net_629 ) , 
    .p610 ( optlc_net_630 ) , .p611 ( optlc_net_631 ) , 
    .p612 ( optlc_net_632 ) , .p613 ( optlc_net_633 ) , 
    .p614 ( optlc_net_634 ) , .p615 ( optlc_net_635 ) , 
    .p616 ( optlc_net_636 ) , .p617 ( optlc_net_637 ) , 
    .p618 ( optlc_net_638 ) , .p619 ( optlc_net_639 ) , 
    .p620 ( optlc_net_640 ) , .p621 ( optlc_net_641 ) , 
    .p622 ( optlc_net_642 ) , .p623 ( optlc_net_643 ) , 
    .p624 ( optlc_net_644 ) , .p625 ( optlc_net_645 ) , 
    .p626 ( optlc_net_646 ) , .p627 ( optlc_net_647 ) , 
    .p628 ( optlc_net_648 ) , .p629 ( optlc_net_649 ) , 
    .p630 ( optlc_net_650 ) , .p631 ( optlc_net_651 ) , 
    .p632 ( optlc_net_652 ) , .p633 ( optlc_net_653 ) , 
    .p634 ( optlc_net_654 ) , .p635 ( optlc_net_655 ) , 
    .p636 ( optlc_net_656 ) , .p637 ( optlc_net_657 ) , 
    .p638 ( optlc_net_658 ) , .p639 ( optlc_net_659 ) , 
    .p640 ( optlc_net_660 ) , .p641 ( optlc_net_661 ) , 
    .p642 ( optlc_net_662 ) , .p643 ( optlc_net_663 ) , 
    .p644 ( optlc_net_664 ) , .p645 ( optlc_net_665 ) , 
    .p646 ( optlc_net_666 ) , .p647 ( optlc_net_667 ) , 
    .p648 ( optlc_net_668 ) , .p649 ( optlc_net_669 ) , 
    .p650 ( optlc_net_670 ) , .p651 ( optlc_net_671 ) , 
    .p652 ( optlc_net_672 ) , .p653 ( optlc_net_673 ) , 
    .p654 ( optlc_net_674 ) , .p655 ( optlc_net_675 ) , 
    .p656 ( optlc_net_676 ) , .p657 ( optlc_net_677 ) , 
    .p658 ( optlc_net_678 ) , .p659 ( optlc_net_679 ) , 
    .p660 ( optlc_net_680 ) , .p661 ( optlc_net_681 ) , 
    .p662 ( optlc_net_682 ) , .p663 ( optlc_net_683 ) , 
    .p664 ( optlc_net_684 ) , .p665 ( optlc_net_685 ) , 
    .p666 ( optlc_net_686 ) , .p667 ( optlc_net_687 ) , 
    .p668 ( optlc_net_688 ) , .p669 ( optlc_net_689 ) , 
    .p670 ( optlc_net_690 ) , .p671 ( optlc_net_691 ) , 
    .p672 ( optlc_net_692 ) , .p673 ( optlc_net_693 ) , 
    .p674 ( optlc_net_694 ) , .p675 ( optlc_net_695 ) , 
    .p676 ( optlc_net_696 ) , .p677 ( optlc_net_697 ) , 
    .p678 ( optlc_net_698 ) , .p679 ( optlc_net_699 ) , 
    .p680 ( optlc_net_700 ) , .p681 ( optlc_net_701 ) , 
    .p682 ( optlc_net_702 ) , .p683 ( optlc_net_703 ) , 
    .p684 ( optlc_net_704 ) , .p685 ( optlc_net_705 ) , 
    .p686 ( optlc_net_706 ) , .p687 ( optlc_net_707 ) , 
    .p688 ( optlc_net_708 ) , .p689 ( optlc_net_709 ) , 
    .p690 ( optlc_net_710 ) , .p691 ( optlc_net_711 ) , 
    .p692 ( optlc_net_712 ) , .p693 ( optlc_net_713 ) , 
    .p694 ( optlc_net_714 ) , .p695 ( optlc_net_715 ) , 
    .p696 ( optlc_net_716 ) , .p697 ( optlc_net_717 ) , 
    .p698 ( optlc_net_718 ) , .p699 ( optlc_net_719 ) , 
    .p700 ( optlc_net_720 ) , .p701 ( optlc_net_721 ) , 
    .p702 ( optlc_net_722 ) , .p703 ( optlc_net_723 ) , 
    .p704 ( optlc_net_724 ) , .p705 ( optlc_net_725 ) , 
    .p706 ( optlc_net_726 ) , .p707 ( optlc_net_727 ) , 
    .p708 ( optlc_net_728 ) , .p709 ( optlc_net_729 ) , 
    .p710 ( optlc_net_730 ) , .p711 ( optlc_net_731 ) , 
    .p712 ( optlc_net_732 ) , .p713 ( optlc_net_733 ) , 
    .p714 ( optlc_net_734 ) , .p715 ( optlc_net_735 ) , 
    .p716 ( optlc_net_736 ) , .p717 ( optlc_net_737 ) , 
    .p718 ( optlc_net_738 ) , .p719 ( optlc_net_739 ) , 
    .p720 ( optlc_net_740 ) , .p721 ( optlc_net_741 ) , 
    .p722 ( optlc_net_742 ) , .p723 ( optlc_net_743 ) , 
    .p724 ( optlc_net_744 ) , .p725 ( optlc_net_745 ) , 
    .p726 ( optlc_net_746 ) , .p727 ( optlc_net_747 ) , 
    .p728 ( optlc_net_748 ) , .p729 ( optlc_net_749 ) , 
    .p730 ( optlc_net_750 ) , .p731 ( optlc_net_751 ) , 
    .p732 ( optlc_net_752 ) , .p733 ( optlc_net_753 ) , 
    .p734 ( optlc_net_754 ) , .p735 ( optlc_net_755 ) , 
    .p736 ( optlc_net_756 ) , .p737 ( optlc_net_757 ) , 
    .p738 ( optlc_net_758 ) , .p739 ( optlc_net_759 ) , 
    .p740 ( optlc_net_760 ) , .p741 ( optlc_net_761 ) , 
    .p742 ( optlc_net_762 ) , .p743 ( optlc_net_763 ) , 
    .p744 ( optlc_net_764 ) , .p745 ( optlc_net_765 ) , 
    .p746 ( optlc_net_766 ) , .p747 ( optlc_net_767 ) , 
    .p748 ( optlc_net_768 ) , .p749 ( optlc_net_769 ) , 
    .p750 ( optlc_net_770 ) , .p751 ( optlc_net_771 ) , 
    .p752 ( optlc_net_772 ) , .p753 ( optlc_net_773 ) , 
    .p754 ( optlc_net_774 ) , .p755 ( optlc_net_775 ) , 
    .p756 ( optlc_net_776 ) , .p757 ( optlc_net_777 ) , 
    .p758 ( optlc_net_778 ) , .p759 ( optlc_net_779 ) , 
    .p760 ( optlc_net_780 ) , .p761 ( optlc_net_781 ) , 
    .p762 ( optlc_net_782 ) , .p763 ( optlc_net_783 ) , 
    .p764 ( optlc_net_784 ) , .p765 ( optlc_net_785 ) , 
    .p766 ( optlc_net_786 ) , .p767 ( optlc_net_787 ) , 
    .p768 ( optlc_net_788 ) , .p769 ( optlc_net_789 ) , 
    .p770 ( optlc_net_790 ) , .p771 ( optlc_net_791 ) , 
    .p772 ( optlc_net_792 ) , .p773 ( optlc_net_793 ) , 
    .p774 ( optlc_net_794 ) , .p775 ( optlc_net_795 ) , 
    .p776 ( optlc_net_796 ) , .p777 ( optlc_net_797 ) , 
    .p778 ( optlc_net_798 ) , .p779 ( optlc_net_799 ) , 
    .p780 ( optlc_net_800 ) , .p781 ( optlc_net_801 ) , 
    .p782 ( optlc_net_802 ) , .p783 ( optlc_net_803 ) , 
    .p784 ( optlc_net_804 ) , .p785 ( optlc_net_805 ) , 
    .p786 ( optlc_net_806 ) , .p787 ( optlc_net_807 ) , 
    .p788 ( optlc_net_808 ) , .p789 ( optlc_net_809 ) , 
    .p790 ( optlc_net_810 ) , .p791 ( optlc_net_811 ) , 
    .p792 ( optlc_net_812 ) , .p793 ( optlc_net_813 ) , 
    .p794 ( optlc_net_814 ) , .p795 ( optlc_net_815 ) , 
    .p796 ( optlc_net_816 ) , .p797 ( optlc_net_817 ) , 
    .p798 ( optlc_net_818 ) , .p799 ( optlc_net_819 ) , 
    .p800 ( optlc_net_820 ) , .p801 ( optlc_net_821 ) , 
    .p802 ( optlc_net_822 ) , .p803 ( optlc_net_823 ) , 
    .p804 ( optlc_net_824 ) , .p805 ( optlc_net_825 ) , 
    .p806 ( optlc_net_826 ) , .p807 ( optlc_net_827 ) , 
    .p808 ( optlc_net_828 ) , .p809 ( optlc_net_829 ) , 
    .p810 ( optlc_net_830 ) , .p811 ( optlc_net_831 ) , 
    .p812 ( optlc_net_832 ) , .p813 ( optlc_net_833 ) , 
    .p814 ( optlc_net_834 ) , .p815 ( optlc_net_835 ) , 
    .p816 ( optlc_net_836 ) , .p817 ( optlc_net_837 ) , 
    .p818 ( optlc_net_838 ) , .p819 ( optlc_net_839 ) , 
    .p820 ( optlc_net_840 ) , .p821 ( optlc_net_841 ) , 
    .p822 ( optlc_net_842 ) , .p823 ( optlc_net_843 ) , 
    .p824 ( optlc_net_844 ) , .p825 ( optlc_net_845 ) , 
    .p826 ( optlc_net_846 ) , .p827 ( optlc_net_847 ) , 
    .p828 ( optlc_net_848 ) , .p829 ( optlc_net_849 ) , 
    .p830 ( optlc_net_850 ) , .p831 ( optlc_net_851 ) , 
    .p832 ( optlc_net_852 ) , .p833 ( optlc_net_853 ) , 
    .p834 ( optlc_net_854 ) , .p835 ( optlc_net_855 ) , 
    .p836 ( optlc_net_856 ) , .p837 ( optlc_net_857 ) , 
    .p838 ( optlc_net_858 ) , .p839 ( optlc_net_859 ) , 
    .p840 ( optlc_net_860 ) , .p841 ( optlc_net_861 ) , 
    .p842 ( optlc_net_862 ) , .p843 ( optlc_net_863 ) , 
    .p844 ( optlc_net_864 ) , .p845 ( optlc_net_865 ) , 
    .p846 ( optlc_net_866 ) , .p847 ( optlc_net_867 ) , 
    .p848 ( optlc_net_868 ) , .p849 ( optlc_net_869 ) , 
    .p850 ( optlc_net_870 ) , .p851 ( optlc_net_871 ) , 
    .p852 ( optlc_net_872 ) , .p853 ( optlc_net_873 ) , 
    .p854 ( optlc_net_874 ) , .p855 ( optlc_net_875 ) , 
    .p856 ( optlc_net_876 ) , .p857 ( optlc_net_877 ) , 
    .p858 ( optlc_net_878 ) , .p859 ( optlc_net_879 ) , 
    .p860 ( optlc_net_880 ) , .p861 ( optlc_net_881 ) , 
    .p862 ( optlc_net_882 ) , .p863 ( optlc_net_883 ) , 
    .p864 ( optlc_net_884 ) , .p865 ( optlc_net_885 ) , 
    .p866 ( optlc_net_886 ) , .p867 ( optlc_net_887 ) , 
    .p868 ( optlc_net_888 ) , .p869 ( optlc_net_889 ) , 
    .p870 ( optlc_net_890 ) , .p871 ( optlc_net_891 ) , 
    .p872 ( optlc_net_892 ) , .p873 ( optlc_net_893 ) , 
    .p874 ( optlc_net_894 ) , .p875 ( optlc_net_895 ) , 
    .p876 ( optlc_net_896 ) , .p877 ( optlc_net_897 ) , 
    .p878 ( optlc_net_898 ) , .p879 ( optlc_net_899 ) , 
    .p880 ( optlc_net_900 ) , .p881 ( optlc_net_901 ) , 
    .p882 ( optlc_net_902 ) , .p883 ( optlc_net_903 ) , 
    .p884 ( optlc_net_904 ) , .p885 ( optlc_net_905 ) , 
    .p886 ( optlc_net_906 ) , .p887 ( optlc_net_907 ) , 
    .p888 ( optlc_net_908 ) , .p889 ( optlc_net_909 ) , 
    .p890 ( optlc_net_910 ) , .p891 ( optlc_net_911 ) , 
    .p892 ( optlc_net_912 ) , .p893 ( optlc_net_913 ) , 
    .p894 ( optlc_net_914 ) , .p895 ( optlc_net_915 ) , 
    .p896 ( optlc_net_916 ) , .p897 ( optlc_net_917 ) , 
    .p898 ( optlc_net_918 ) , .p899 ( optlc_net_919 ) , 
    .p900 ( optlc_net_920 ) , .p901 ( optlc_net_921 ) , 
    .p902 ( optlc_net_922 ) , .p903 ( optlc_net_923 ) , 
    .p904 ( optlc_net_924 ) , .p905 ( optlc_net_925 ) , 
    .p906 ( optlc_net_926 ) , .p907 ( optlc_net_927 ) , 
    .p908 ( optlc_net_928 ) , .p909 ( optlc_net_929 ) , 
    .p910 ( optlc_net_930 ) , .p911 ( optlc_net_931 ) , 
    .p912 ( optlc_net_932 ) , .p913 ( optlc_net_933 ) , 
    .p914 ( optlc_net_934 ) , .p915 ( optlc_net_935 ) , 
    .p916 ( optlc_net_936 ) , .p917 ( optlc_net_937 ) , 
    .p918 ( optlc_net_938 ) , .p919 ( optlc_net_939 ) , 
    .p920 ( optlc_net_940 ) , .p921 ( optlc_net_941 ) , 
    .p922 ( optlc_net_942 ) , .p923 ( optlc_net_943 ) , 
    .p924 ( optlc_net_944 ) , .p925 ( optlc_net_945 ) , 
    .p926 ( optlc_net_946 ) , .p927 ( optlc_net_947 ) , 
    .p928 ( optlc_net_948 ) , .p929 ( optlc_net_949 ) , 
    .p930 ( optlc_net_950 ) , .p931 ( optlc_net_951 ) , 
    .p932 ( optlc_net_952 ) , .p933 ( optlc_net_953 ) , 
    .p934 ( optlc_net_954 ) , .p935 ( optlc_net_955 ) , 
    .p936 ( optlc_net_956 ) , .p937 ( optlc_net_957 ) , 
    .p938 ( optlc_net_958 ) , .p939 ( optlc_net_959 ) , 
    .p940 ( optlc_net_960 ) , .p941 ( optlc_net_961 ) , 
    .p942 ( optlc_net_962 ) , .p943 ( optlc_net_963 ) , 
    .p944 ( optlc_net_964 ) , .p945 ( optlc_net_965 ) , 
    .p946 ( optlc_net_966 ) , .p947 ( optlc_net_967 ) , 
    .p948 ( optlc_net_968 ) , .p949 ( optlc_net_969 ) , 
    .p950 ( optlc_net_970 ) , .p951 ( optlc_net_971 ) , 
    .p952 ( optlc_net_972 ) , .p953 ( optlc_net_973 ) , 
    .p954 ( optlc_net_974 ) , .p955 ( optlc_net_975 ) , 
    .p956 ( optlc_net_976 ) , .p957 ( optlc_net_977 ) , 
    .p958 ( optlc_net_978 ) , .p959 ( optlc_net_979 ) , 
    .p960 ( optlc_net_980 ) , .p961 ( optlc_net_981 ) , 
    .p962 ( optlc_net_982 ) , .p963 ( optlc_net_983 ) , 
    .p964 ( optlc_net_984 ) , .p965 ( optlc_net_985 ) , 
    .p966 ( optlc_net_986 ) , .p967 ( optlc_net_987 ) , 
    .p968 ( optlc_net_988 ) , .p969 ( optlc_net_989 ) , 
    .p970 ( optlc_net_990 ) , .p971 ( optlc_net_991 ) , 
    .p972 ( optlc_net_992 ) , .p973 ( optlc_net_993 ) , 
    .p974 ( optlc_net_994 ) , .p975 ( optlc_net_995 ) , 
    .p976 ( optlc_net_996 ) , .p977 ( optlc_net_997 ) , 
    .p978 ( optlc_net_998 ) , .p979 ( optlc_net_999 ) , 
    .p980 ( optlc_net_1000 ) , .p981 ( optlc_net_1001 ) , 
    .p982 ( optlc_net_1002 ) , .p983 ( optlc_net_1003 ) , 
    .p984 ( optlc_net_1004 ) , .p985 ( optlc_net_1005 ) , 
    .p986 ( optlc_net_1006 ) , .p987 ( optlc_net_1007 ) , 
    .p988 ( optlc_net_1008 ) , .p989 ( optlc_net_1009 ) , 
    .p990 ( optlc_net_1010 ) , .p991 ( optlc_net_1011 ) , 
    .p992 ( optlc_net_1012 ) , .p993 ( optlc_net_1013 ) , 
    .p994 ( optlc_net_1014 ) , .p995 ( optlc_net_1015 ) , 
    .p996 ( optlc_net_1016 ) , .p997 ( optlc_net_1017 ) , 
    .p998 ( optlc_net_1018 ) , .p999 ( optlc_net_1019 ) , 
    .p1000 ( optlc_net_1020 ) , .p1001 ( optlc_net_1021 ) , 
    .p1002 ( optlc_net_1022 ) , .p1003 ( optlc_net_1023 ) , 
    .p1004 ( optlc_net_1024 ) , .p1005 ( optlc_net_1025 ) , 
    .p1006 ( optlc_net_1026 ) , .p1007 ( optlc_net_1027 ) , 
    .p1008 ( optlc_net_1028 ) , .p1009 ( optlc_net_1029 ) , 
    .p1010 ( optlc_net_1030 ) , .p1011 ( optlc_net_1031 ) , 
    .p1012 ( optlc_net_1032 ) , .p1013 ( optlc_net_1033 ) , 
    .p1014 ( optlc_net_1034 ) , .p1015 ( optlc_net_1035 ) , 
    .p1016 ( optlc_net_1036 ) , .p1017 ( optlc_net_1037 ) , 
    .p1018 ( optlc_net_1038 ) , .p1019 ( optlc_net_1039 ) , 
    .p1020 ( optlc_net_1040 ) , .p1021 ( optlc_net_1041 ) , 
    .p1022 ( optlc_net_1042 ) , .p1023 ( optlc_net_1043 ) , 
    .p1024 ( optlc_net_1044 ) , .p1025 ( optlc_net_1045 ) , 
    .p1026 ( optlc_net_1046 ) , .p1027 ( optlc_net_1047 ) , 
    .p1028 ( optlc_net_1048 ) , .p1029 ( optlc_net_1049 ) , 
    .p1030 ( optlc_net_1050 ) , .p1031 ( optlc_net_1051 ) , 
    .p1032 ( optlc_net_1052 ) , .p1033 ( optlc_net_1053 ) , 
    .p1034 ( optlc_net_1054 ) , .p1035 ( optlc_net_1055 ) , 
    .p1036 ( optlc_net_1056 ) , .p1037 ( optlc_net_1057 ) , 
    .p1038 ( optlc_net_1058 ) , .p1039 ( optlc_net_1059 ) , 
    .p1040 ( optlc_net_1060 ) , .p1041 ( optlc_net_1061 ) , 
    .p1042 ( optlc_net_1062 ) , .p1043 ( optlc_net_1063 ) , 
    .p1044 ( optlc_net_1064 ) , .p1045 ( optlc_net_1065 ) , 
    .p1046 ( optlc_net_1066 ) , .p1047 ( optlc_net_1067 ) , 
    .p1048 ( optlc_net_1068 ) , .p1049 ( optlc_net_1069 ) , 
    .p1050 ( optlc_net_1070 ) , .p1051 ( optlc_net_1071 ) , 
    .p1052 ( optlc_net_1072 ) , .p1053 ( optlc_net_1073 ) , 
    .p1054 ( optlc_net_1074 ) , .p1055 ( optlc_net_1075 ) , 
    .p1056 ( optlc_net_1076 ) , .p1057 ( optlc_net_1077 ) , 
    .p1058 ( optlc_net_1078 ) , .p1059 ( optlc_net_1079 ) , 
    .p1060 ( optlc_net_1080 ) , .p1061 ( optlc_net_1081 ) , 
    .p1062 ( optlc_net_1082 ) , .p1063 ( optlc_net_1083 ) , 
    .p1064 ( optlc_net_1084 ) , .p1065 ( optlc_net_1085 ) , 
    .p1066 ( optlc_net_1086 ) , .p1067 ( optlc_net_1087 ) , 
    .p1068 ( optlc_net_1088 ) , .p1069 ( optlc_net_1089 ) , 
    .p1070 ( optlc_net_1090 ) , .p1071 ( optlc_net_1091 ) , 
    .p1072 ( optlc_net_1092 ) , .p1073 ( optlc_net_1093 ) , 
    .p1074 ( optlc_net_1094 ) , .p1075 ( optlc_net_1095 ) , 
    .p1076 ( optlc_net_1096 ) , .p1077 ( optlc_net_1097 ) , 
    .p1078 ( optlc_net_1098 ) , .p1079 ( optlc_net_1099 ) , 
    .p1080 ( optlc_net_1100 ) , .p1081 ( optlc_net_1101 ) , 
    .p1082 ( optlc_net_1102 ) , .p1083 ( optlc_net_1103 ) , 
    .p1084 ( optlc_net_1104 ) , .p1085 ( optlc_net_1105 ) , 
    .p1086 ( optlc_net_1106 ) , .p1087 ( optlc_net_1107 ) , 
    .p1088 ( optlc_net_1108 ) , .p1089 ( optlc_net_1109 ) , 
    .p1090 ( optlc_net_1110 ) , .p1091 ( optlc_net_1111 ) , 
    .p1092 ( optlc_net_1112 ) , .p1093 ( optlc_net_1113 ) , 
    .p1094 ( optlc_net_1114 ) , .p1095 ( optlc_net_1115 ) , 
    .p1096 ( optlc_net_1116 ) , .p1097 ( optlc_net_1117 ) , 
    .p1098 ( optlc_net_1118 ) , .p1099 ( optlc_net_1119 ) , 
    .p1100 ( optlc_net_1120 ) , .p1101 ( optlc_net_1121 ) , 
    .p1102 ( optlc_net_1122 ) , .p1103 ( optlc_net_1123 ) , 
    .p1104 ( optlc_net_1124 ) , .p1105 ( optlc_net_1125 ) , 
    .p1106 ( optlc_net_1126 ) , .p1107 ( optlc_net_1127 ) , 
    .p1108 ( optlc_net_1128 ) , .p1109 ( optlc_net_1129 ) , 
    .p1110 ( optlc_net_1130 ) , .p1111 ( optlc_net_1131 ) , 
    .p1112 ( optlc_net_1132 ) , .p1113 ( optlc_net_1133 ) , 
    .p1114 ( optlc_net_1134 ) , .p1115 ( optlc_net_1135 ) , 
    .p1116 ( optlc_net_1136 ) , .p1117 ( optlc_net_1137 ) , 
    .p1118 ( optlc_net_1138 ) , .p1119 ( optlc_net_1139 ) , 
    .p1120 ( optlc_net_1140 ) , .p1121 ( optlc_net_1141 ) , 
    .p1122 ( optlc_net_1142 ) , .p1123 ( optlc_net_1143 ) , 
    .p1124 ( optlc_net_1144 ) , .p1125 ( optlc_net_1145 ) , 
    .p1126 ( optlc_net_1146 ) , .p1127 ( optlc_net_1147 ) , 
    .p1128 ( optlc_net_1148 ) , .p1129 ( optlc_net_1149 ) , 
    .p1130 ( optlc_net_1150 ) , .p1131 ( optlc_net_1151 ) , 
    .p1132 ( optlc_net_1152 ) , .p1133 ( optlc_net_1153 ) , 
    .p1134 ( optlc_net_1154 ) , .p1135 ( optlc_net_1155 ) , 
    .p1136 ( optlc_net_1156 ) , .p1137 ( optlc_net_1157 ) , 
    .p1138 ( optlc_net_1158 ) , .p1139 ( optlc_net_1159 ) , 
    .p1140 ( optlc_net_1160 ) , .p1141 ( optlc_net_1161 ) , 
    .p1142 ( optlc_net_1162 ) , .p1143 ( optlc_net_1163 ) , 
    .p1144 ( optlc_net_1164 ) , .p1145 ( optlc_net_1165 ) , 
    .p1146 ( optlc_net_1166 ) , .p1147 ( optlc_net_1167 ) , 
    .p1148 ( optlc_net_1168 ) , .p1149 ( optlc_net_1169 ) , 
    .p1150 ( optlc_net_1170 ) , .p1151 ( optlc_net_1171 ) , 
    .p1152 ( optlc_net_1172 ) , .p1153 ( optlc_net_1173 ) , 
    .p1154 ( optlc_net_1174 ) , .p1155 ( optlc_net_1175 ) , 
    .p1156 ( optlc_net_1176 ) , .p1157 ( optlc_net_1177 ) , 
    .p1158 ( optlc_net_1178 ) , .p1159 ( optlc_net_1179 ) , 
    .p1160 ( optlc_net_1180 ) , .p1161 ( optlc_net_1181 ) , 
    .p1162 ( optlc_net_1182 ) , .p1163 ( optlc_net_1183 ) , 
    .p1164 ( optlc_net_1184 ) , .p1165 ( optlc_net_1185 ) , 
    .p1166 ( optlc_net_1186 ) , .p1167 ( optlc_net_1187 ) , 
    .p1168 ( optlc_net_1188 ) , .p1169 ( optlc_net_1189 ) , 
    .p1170 ( optlc_net_1190 ) , .p1171 ( optlc_net_1191 ) , 
    .p1172 ( optlc_net_1192 ) , .p1173 ( optlc_net_1193 ) , 
    .p1174 ( optlc_net_1194 ) , .p1175 ( optlc_net_1195 ) , 
    .p1176 ( optlc_net_1196 ) , .p1177 ( optlc_net_1197 ) , 
    .p1178 ( optlc_net_1198 ) , .p1179 ( optlc_net_1199 ) , 
    .p1180 ( optlc_net_1200 ) , .p1181 ( optlc_net_1201 ) , 
    .p1182 ( optlc_net_1202 ) , .p1183 ( optlc_net_1203 ) , 
    .p1184 ( optlc_net_1204 ) , .p1185 ( optlc_net_1205 ) , 
    .p1186 ( optlc_net_1206 ) , .p1187 ( optlc_net_1207 ) , 
    .p1188 ( optlc_net_1208 ) , .p1189 ( optlc_net_1209 ) , 
    .p1190 ( optlc_net_1210 ) , .p1191 ( optlc_net_1211 ) , 
    .p1192 ( optlc_net_1212 ) , .p1193 ( optlc_net_1213 ) , 
    .p1194 ( optlc_net_1214 ) , .p1195 ( optlc_net_1215 ) , 
    .p1196 ( optlc_net_1216 ) , .p1197 ( optlc_net_1217 ) , 
    .p1198 ( optlc_net_1218 ) , .p1199 ( optlc_net_1219 ) , 
    .p1200 ( optlc_net_1220 ) , .p1201 ( optlc_net_1221 ) , 
    .p1202 ( optlc_net_1222 ) , .p1203 ( optlc_net_1223 ) , 
    .p1204 ( optlc_net_1224 ) , .p1205 ( optlc_net_1225 ) , 
    .p1206 ( optlc_net_1226 ) , .p1207 ( optlc_net_1227 ) , 
    .p1208 ( optlc_net_1228 ) , .p1209 ( optlc_net_1229 ) , 
    .p1210 ( optlc_net_1230 ) , .p1211 ( optlc_net_1231 ) , 
    .p1212 ( optlc_net_1232 ) , .p1213 ( optlc_net_1233 ) , 
    .p1214 ( optlc_net_1234 ) , .p1215 ( optlc_net_1235 ) , 
    .p1216 ( optlc_net_1236 ) , .p1217 ( optlc_net_1237 ) , 
    .p1218 ( optlc_net_1238 ) , .p1219 ( optlc_net_1239 ) , 
    .p1220 ( optlc_net_1240 ) , .p1221 ( optlc_net_1241 ) , 
    .p1222 ( optlc_net_1242 ) , .p1223 ( optlc_net_1243 ) , 
    .p1224 ( optlc_net_1244 ) , .p1225 ( optlc_net_1245 ) , 
    .p1226 ( optlc_net_1246 ) , .p1227 ( optlc_net_1247 ) , 
    .p1228 ( optlc_net_1248 ) , .p1229 ( optlc_net_1249 ) , 
    .p1230 ( optlc_net_1250 ) , .p1231 ( optlc_net_1251 ) , 
    .p1232 ( optlc_net_1252 ) , .p1233 ( optlc_net_1253 ) , 
    .p1234 ( optlc_net_1254 ) , .p1235 ( optlc_net_1255 ) , 
    .p1236 ( optlc_net_1256 ) , .p1237 ( optlc_net_1257 ) , 
    .p1238 ( optlc_net_1258 ) , .p1239 ( optlc_net_1259 ) , 
    .p1240 ( optlc_net_1260 ) , .p1241 ( optlc_net_1261 ) , 
    .p1242 ( optlc_net_1262 ) , .p1243 ( optlc_net_1263 ) , 
    .p1244 ( optlc_net_1264 ) , .p1245 ( optlc_net_1265 ) , 
    .p1246 ( optlc_net_1266 ) , .p1247 ( optlc_net_1267 ) , 
    .p1248 ( optlc_net_1268 ) , .p1249 ( optlc_net_1269 ) , 
    .p1250 ( optlc_net_1270 ) , .p1251 ( optlc_net_1271 ) , 
    .p1252 ( optlc_net_1272 ) , .p1253 ( optlc_net_1273 ) , 
    .p1254 ( optlc_net_1274 ) , .p1255 ( optlc_net_1275 ) , 
    .p1256 ( optlc_net_1276 ) , .p1257 ( optlc_net_1277 ) , 
    .p1258 ( optlc_net_1278 ) , .p1259 ( optlc_net_1279 ) , 
    .p1260 ( optlc_net_1280 ) , .p1261 ( optlc_net_1281 ) , 
    .p1262 ( optlc_net_1282 ) , .p1263 ( optlc_net_1283 ) , 
    .p1264 ( optlc_net_1284 ) , .p1265 ( optlc_net_1285 ) , 
    .p1266 ( optlc_net_1286 ) , .p1267 ( optlc_net_1287 ) , 
    .p1268 ( optlc_net_1288 ) , .p1269 ( optlc_net_1289 ) , 
    .p1270 ( optlc_net_1290 ) , .p1271 ( optlc_net_1291 ) , 
    .p1272 ( optlc_net_1292 ) , .p1273 ( optlc_net_1293 ) , 
    .p1274 ( optlc_net_1294 ) , .p1275 ( optlc_net_1295 ) , 
    .p1276 ( optlc_net_1296 ) , .p1277 ( optlc_net_1297 ) , 
    .p1278 ( optlc_net_1298 ) , .p1279 ( optlc_net_1299 ) , 
    .p1280 ( optlc_net_1300 ) , .p1281 ( optlc_net_1301 ) , 
    .p1282 ( optlc_net_1302 ) , .p1283 ( optlc_net_1303 ) , 
    .p1284 ( optlc_net_1304 ) , .p1285 ( optlc_net_1305 ) , 
    .p1286 ( optlc_net_1306 ) , .p1287 ( optlc_net_1307 ) , 
    .p1288 ( optlc_net_1308 ) , .p1289 ( optlc_net_1309 ) , 
    .p1290 ( optlc_net_1310 ) , .p1291 ( optlc_net_1311 ) , 
    .p1292 ( optlc_net_1312 ) , .p1293 ( optlc_net_1313 ) , 
    .p1294 ( optlc_net_1314 ) , .p1295 ( optlc_net_1315 ) , 
    .p1296 ( optlc_net_1316 ) , .p1297 ( optlc_net_1317 ) , 
    .p1298 ( optlc_net_1318 ) , .p1299 ( optlc_net_1319 ) , 
    .p1300 ( optlc_net_1320 ) , .p1301 ( optlc_net_1321 ) , 
    .p1302 ( optlc_net_1322 ) , .p1303 ( optlc_net_1323 ) , 
    .p1304 ( optlc_net_1324 ) , .p1305 ( optlc_net_1325 ) , 
    .p1306 ( optlc_net_1326 ) , .p1307 ( optlc_net_1327 ) , 
    .p1308 ( optlc_net_1328 ) , .p1309 ( optlc_net_1329 ) , 
    .p1310 ( optlc_net_1330 ) , .p1311 ( optlc_net_1331 ) , 
    .p1312 ( optlc_net_1332 ) , .p1313 ( optlc_net_1333 ) , 
    .p1314 ( optlc_net_1334 ) , .p1315 ( optlc_net_1335 ) , 
    .p1316 ( optlc_net_1336 ) , .p1317 ( optlc_net_1337 ) , 
    .p1318 ( optlc_net_1338 ) , .p1319 ( optlc_net_1339 ) , 
    .p1320 ( optlc_net_1340 ) , .p1321 ( optlc_net_1341 ) , 
    .p1322 ( optlc_net_1342 ) , .p1323 ( optlc_net_1343 ) , 
    .p1324 ( optlc_net_1344 ) , .p1325 ( optlc_net_1345 ) , 
    .p1326 ( optlc_net_1346 ) , .p1327 ( optlc_net_1347 ) , 
    .p1328 ( optlc_net_1348 ) , .p1329 ( optlc_net_1349 ) , 
    .p1330 ( optlc_net_1350 ) , .p1331 ( optlc_net_1351 ) , 
    .p1332 ( optlc_net_1352 ) , .p1333 ( optlc_net_1353 ) , 
    .p1334 ( optlc_net_1354 ) , .p1335 ( optlc_net_1355 ) , 
    .p1336 ( optlc_net_1356 ) , .p1337 ( optlc_net_1357 ) , 
    .p1338 ( optlc_net_1358 ) , .p1339 ( optlc_net_1359 ) , 
    .p1340 ( optlc_net_1360 ) , .p1341 ( optlc_net_1361 ) , 
    .p1342 ( optlc_net_1362 ) , .p1343 ( optlc_net_1363 ) , 
    .p1344 ( optlc_net_1364 ) , .p1345 ( optlc_net_1365 ) , 
    .p1346 ( optlc_net_1366 ) , .p1347 ( optlc_net_1367 ) , 
    .p1348 ( optlc_net_1368 ) , .p1349 ( optlc_net_1369 ) , 
    .p1350 ( optlc_net_1370 ) , .p1351 ( optlc_net_1371 ) , 
    .p1352 ( optlc_net_1372 ) , .p1353 ( optlc_net_1373 ) , 
    .p1354 ( optlc_net_1374 ) , .p1355 ( optlc_net_1375 ) , 
    .p1356 ( optlc_net_1376 ) , .p1357 ( optlc_net_1377 ) , 
    .p1358 ( optlc_net_1378 ) , .p1359 ( optlc_net_1379 ) , 
    .p1360 ( optlc_net_1380 ) , .p1361 ( optlc_net_1381 ) , 
    .p1362 ( optlc_net_1382 ) , .p1363 ( optlc_net_1383 ) , 
    .p1364 ( optlc_net_1384 ) , .p1365 ( optlc_net_1385 ) , 
    .p1366 ( optlc_net_1386 ) , .p1367 ( optlc_net_1387 ) , 
    .p1368 ( optlc_net_1388 ) , .p1369 ( optlc_net_1389 ) , 
    .p1370 ( optlc_net_1390 ) , .p1371 ( optlc_net_1391 ) , 
    .p1372 ( optlc_net_1392 ) , .p1373 ( optlc_net_1393 ) , 
    .p1374 ( optlc_net_1394 ) , .p1375 ( optlc_net_1395 ) , 
    .p1376 ( optlc_net_1396 ) , .p1377 ( optlc_net_1397 ) , 
    .p1378 ( optlc_net_1398 ) , .p1379 ( optlc_net_1399 ) , 
    .p1380 ( optlc_net_1400 ) , .p1381 ( optlc_net_1401 ) , 
    .p1382 ( optlc_net_1402 ) , .p1383 ( optlc_net_1403 ) , 
    .p1384 ( optlc_net_1404 ) , .p1385 ( optlc_net_1405 ) , 
    .p1386 ( optlc_net_1406 ) , .p1387 ( optlc_net_1407 ) , 
    .p1388 ( optlc_net_1408 ) , .p1389 ( optlc_net_1409 ) , 
    .p1390 ( optlc_net_1410 ) , .p1391 ( optlc_net_1411 ) , 
    .p1392 ( optlc_net_1412 ) , .p1393 ( optlc_net_1413 ) , 
    .p1394 ( optlc_net_1414 ) , .p1395 ( optlc_net_1415 ) , 
    .p1396 ( optlc_net_1416 ) , .p1397 ( optlc_net_1417 ) , 
    .p1398 ( optlc_net_1418 ) , .p1399 ( optlc_net_1419 ) , 
    .p1400 ( optlc_net_1420 ) , .p1401 ( optlc_net_1421 ) , 
    .p1402 ( optlc_net_1422 ) , .p1403 ( optlc_net_1423 ) , 
    .p1404 ( optlc_net_1424 ) , .p1405 ( optlc_net_1425 ) , 
    .p1406 ( optlc_net_1426 ) , .p1407 ( optlc_net_1427 ) , 
    .p1408 ( optlc_net_1428 ) , .p1409 ( optlc_net_1429 ) , 
    .p1410 ( optlc_net_1430 ) , .p1411 ( optlc_net_1431 ) , 
    .p1412 ( optlc_net_1432 ) , .p1413 ( optlc_net_1433 ) , 
    .p1414 ( optlc_net_1434 ) , .p1415 ( optlc_net_1435 ) , 
    .p1416 ( optlc_net_1436 ) , .p1417 ( optlc_net_1437 ) , 
    .p1418 ( optlc_net_1438 ) , .p1419 ( optlc_net_1439 ) , 
    .p1420 ( optlc_net_1440 ) , .p1421 ( optlc_net_1441 ) , 
    .p1422 ( optlc_net_1442 ) , .p1423 ( optlc_net_1443 ) , 
    .p1424 ( optlc_net_1444 ) , .p1425 ( optlc_net_1445 ) , 
    .p1426 ( optlc_net_1446 ) , .p1427 ( optlc_net_1447 ) , 
    .p1428 ( optlc_net_1448 ) , .p1429 ( optlc_net_1449 ) , 
    .p1430 ( optlc_net_1450 ) , .p1431 ( optlc_net_1451 ) , 
    .p1432 ( optlc_net_1452 ) , .p1433 ( optlc_net_1453 ) , 
    .p1434 ( optlc_net_1454 ) , .p1435 ( optlc_net_1455 ) , 
    .p1436 ( optlc_net_1456 ) , .p1437 ( optlc_net_1457 ) , 
    .p1438 ( optlc_net_1458 ) , .p1439 ( optlc_net_1459 ) , 
    .p1440 ( optlc_net_1460 ) , .p1441 ( optlc_net_1461 ) , 
    .p1442 ( optlc_net_1462 ) , .p1443 ( optlc_net_1463 ) , 
    .p1444 ( optlc_net_1464 ) , .p1445 ( optlc_net_1465 ) , 
    .p1446 ( optlc_net_1466 ) , .p1447 ( optlc_net_1467 ) , 
    .p1448 ( optlc_net_1468 ) , .p1449 ( optlc_net_1469 ) , 
    .p1450 ( optlc_net_1470 ) , .p1451 ( optlc_net_1471 ) , 
    .p1452 ( optlc_net_1472 ) , .p1453 ( optlc_net_1473 ) , 
    .p1454 ( optlc_net_1474 ) , .p1455 ( optlc_net_1475 ) , 
    .p1456 ( optlc_net_1476 ) , .p1457 ( optlc_net_1477 ) , 
    .p1458 ( optlc_net_1478 ) , .p1459 ( optlc_net_1479 ) , 
    .p1460 ( optlc_net_1480 ) , .p1461 ( optlc_net_1481 ) , 
    .p1462 ( optlc_net_1482 ) , .p1463 ( optlc_net_1483 ) , 
    .p1464 ( optlc_net_1484 ) , .p1465 ( optlc_net_1485 ) , 
    .p1466 ( optlc_net_1486 ) , .p1467 ( optlc_net_1487 ) , 
    .p1468 ( optlc_net_1488 ) , .p1469 ( optlc_net_1489 ) , 
    .p1470 ( optlc_net_1490 ) , .p1471 ( optlc_net_1491 ) , 
    .p1472 ( optlc_net_1492 ) , .p1473 ( optlc_net_1493 ) , 
    .p1474 ( optlc_net_1494 ) , .p1475 ( optlc_net_1495 ) , 
    .p1476 ( optlc_net_1496 ) , .p1477 ( optlc_net_1497 ) , 
    .p1478 ( optlc_net_1498 ) , .p1479 ( optlc_net_1499 ) , 
    .p1480 ( optlc_net_1500 ) , .p1481 ( optlc_net_1501 ) , 
    .p1482 ( optlc_net_1502 ) , .p1483 ( optlc_net_1503 ) , 
    .p1484 ( optlc_net_1504 ) , .p1485 ( optlc_net_1505 ) , 
    .p1486 ( optlc_net_1506 ) , .p1487 ( optlc_net_1507 ) , 
    .p1488 ( optlc_net_1508 ) , .p1489 ( optlc_net_1509 ) , 
    .p1490 ( optlc_net_1510 ) , .p1491 ( optlc_net_1511 ) , 
    .p1492 ( optlc_net_1512 ) , .p1493 ( optlc_net_1513 ) , 
    .p1494 ( optlc_net_1514 ) , .p1495 ( optlc_net_1515 ) , 
    .p1496 ( optlc_net_1516 ) , .p1497 ( optlc_net_1517 ) , 
    .p1498 ( optlc_net_1518 ) , .p1499 ( optlc_net_1519 ) , 
    .p1500 ( optlc_net_1520 ) , .p1501 ( optlc_net_1521 ) , 
    .p1502 ( optlc_net_1522 ) , .p1503 ( optlc_net_1523 ) , 
    .p1504 ( optlc_net_1524 ) , .p1505 ( optlc_net_1525 ) , 
    .p1506 ( optlc_net_1526 ) , .p1507 ( optlc_net_1527 ) , 
    .p1508 ( optlc_net_1528 ) , .p1509 ( optlc_net_1529 ) , 
    .p1510 ( optlc_net_1530 ) , .p1511 ( optlc_net_1531 ) , 
    .p1512 ( optlc_net_1532 ) , .p1513 ( optlc_net_1533 ) , 
    .p1514 ( optlc_net_1534 ) , .p1515 ( optlc_net_1535 ) , 
    .p1516 ( optlc_net_1536 ) , .p1517 ( optlc_net_1537 ) , 
    .p1518 ( optlc_net_1538 ) , .p1519 ( optlc_net_1539 ) , 
    .p1520 ( optlc_net_1540 ) , .p1521 ( optlc_net_1541 ) , 
    .p1522 ( optlc_net_1542 ) , .p1523 ( optlc_net_1543 ) , 
    .p1524 ( optlc_net_1544 ) , .p1525 ( optlc_net_1545 ) , 
    .p1526 ( optlc_net_1546 ) , .p1527 ( optlc_net_1547 ) , 
    .p1528 ( optlc_net_1548 ) , .p1529 ( optlc_net_1549 ) , 
    .p1530 ( optlc_net_1550 ) , .p1531 ( optlc_net_1551 ) , 
    .p1532 ( optlc_net_1552 ) , .p1533 ( optlc_net_1553 ) , 
    .p1534 ( optlc_net_1554 ) , .p1535 ( optlc_net_1555 ) , 
    .p1536 ( optlc_net_1556 ) , .p1537 ( optlc_net_1557 ) , 
    .p1538 ( optlc_net_1558 ) , .p1539 ( optlc_net_1559 ) , 
    .p1540 ( optlc_net_1560 ) , .p1541 ( optlc_net_1561 ) , 
    .p1542 ( optlc_net_1562 ) , .p1543 ( optlc_net_1563 ) , 
    .p1544 ( optlc_net_1564 ) , .p1545 ( optlc_net_1565 ) , 
    .p1546 ( optlc_net_1566 ) , .p1547 ( optlc_net_1567 ) , 
    .p1548 ( optlc_net_1568 ) , .p1549 ( optlc_net_1569 ) , 
    .p1550 ( optlc_net_1570 ) , .p1551 ( optlc_net_1571 ) , 
    .p1552 ( optlc_net_1572 ) , .p1553 ( optlc_net_1573 ) , 
    .p1554 ( optlc_net_1574 ) , .p1555 ( optlc_net_1575 ) , 
    .p1556 ( optlc_net_1576 ) , .p1557 ( optlc_net_1577 ) , 
    .p1558 ( optlc_net_1578 ) , .p1559 ( optlc_net_1579 ) , 
    .p1560 ( optlc_net_1580 ) , .p1561 ( optlc_net_1581 ) , 
    .p1562 ( optlc_net_1582 ) , .p1563 ( optlc_net_1583 ) , 
    .p1564 ( optlc_net_1584 ) , .p1565 ( optlc_net_1585 ) , 
    .p1566 ( optlc_net_1586 ) , .p1567 ( optlc_net_1587 ) , 
    .p1568 ( optlc_net_1588 ) , .p1569 ( optlc_net_1589 ) , 
    .p1570 ( optlc_net_1590 ) , .p1571 ( optlc_net_1591 ) , 
    .p1572 ( optlc_net_1592 ) , .p1573 ( optlc_net_1593 ) , 
    .p1574 ( optlc_net_1594 ) , .p1575 ( optlc_net_1595 ) , 
    .p1576 ( optlc_net_1596 ) , .p1577 ( optlc_net_1597 ) , 
    .p1578 ( optlc_net_1598 ) , .p1579 ( optlc_net_1599 ) , 
    .p1580 ( optlc_net_1600 ) , .p1581 ( optlc_net_1601 ) , 
    .p1582 ( optlc_net_1602 ) , .p1583 ( optlc_net_1603 ) , 
    .p1584 ( optlc_net_1604 ) , .p1585 ( optlc_net_1605 ) , 
    .p1586 ( optlc_net_1606 ) , .p1587 ( optlc_net_1607 ) , 
    .p1588 ( optlc_net_1608 ) , .p1589 ( optlc_net_1609 ) , 
    .p1590 ( optlc_net_1610 ) , .p1591 ( optlc_net_1611 ) , 
    .p1592 ( optlc_net_1612 ) , .p1593 ( optlc_net_1613 ) , 
    .p1594 ( optlc_net_1614 ) , .p1595 ( optlc_net_1615 ) , 
    .p1596 ( optlc_net_1616 ) , .p1597 ( optlc_net_1617 ) , 
    .p1598 ( optlc_net_1618 ) , .p1599 ( optlc_net_1619 ) , 
    .p1600 ( optlc_net_1620 ) , .p1601 ( optlc_net_1621 ) , 
    .p1602 ( optlc_net_1622 ) , .p1603 ( optlc_net_1623 ) , 
    .p1604 ( optlc_net_1624 ) , .p1605 ( optlc_net_1625 ) , 
    .p1606 ( optlc_net_1626 ) , .p1607 ( optlc_net_1627 ) , 
    .p1608 ( optlc_net_1628 ) , .p1609 ( optlc_net_1629 ) , 
    .p1610 ( optlc_net_1630 ) , .p1611 ( optlc_net_1631 ) , 
    .p1612 ( optlc_net_1632 ) , .p1613 ( optlc_net_1633 ) , 
    .p1614 ( optlc_net_1634 ) , .p1615 ( optlc_net_1635 ) , 
    .p1616 ( optlc_net_1636 ) , .p1617 ( optlc_net_1637 ) , 
    .p1618 ( optlc_net_1638 ) , .p1619 ( optlc_net_1639 ) , 
    .p1620 ( optlc_net_1640 ) , .p1621 ( optlc_net_1641 ) , 
    .p1622 ( optlc_net_1642 ) , .p1623 ( optlc_net_1643 ) , 
    .p1624 ( optlc_net_1644 ) , .p1625 ( optlc_net_1645 ) , 
    .p1626 ( optlc_net_1646 ) , .p1627 ( optlc_net_1647 ) , 
    .p1628 ( optlc_net_1648 ) , .p1629 ( optlc_net_1649 ) , 
    .p1630 ( optlc_net_1650 ) , .p1631 ( optlc_net_1651 ) , 
    .p1632 ( optlc_net_1652 ) , .p1633 ( optlc_net_1653 ) , 
    .p1634 ( optlc_net_1654 ) , .p1635 ( optlc_net_1655 ) , 
    .p1636 ( optlc_net_1656 ) , .p1637 ( optlc_net_1657 ) , 
    .p1638 ( optlc_net_1658 ) , .p1639 ( optlc_net_1659 ) , 
    .p1640 ( optlc_net_1660 ) , .p1641 ( optlc_net_1661 ) , 
    .p1642 ( optlc_net_1662 ) , .p1643 ( optlc_net_1663 ) , 
    .p1644 ( optlc_net_1664 ) , .p1645 ( optlc_net_1665 ) , 
    .p1646 ( optlc_net_1666 ) , .p1647 ( optlc_net_1667 ) , 
    .p1648 ( optlc_net_1668 ) , .p1649 ( optlc_net_1669 ) , 
    .p1650 ( optlc_net_1670 ) , .p1651 ( optlc_net_1671 ) , 
    .p1652 ( optlc_net_1672 ) , .p1653 ( optlc_net_1673 ) , 
    .p1654 ( optlc_net_1674 ) , .p1655 ( optlc_net_1675 ) , 
    .p1656 ( optlc_net_1676 ) , .p1657 ( optlc_net_1677 ) , 
    .p1658 ( optlc_net_1678 ) , .p1659 ( optlc_net_1679 ) , 
    .p1660 ( optlc_net_1680 ) , .p1661 ( optlc_net_1681 ) , 
    .p1662 ( optlc_net_1682 ) , .p1663 ( optlc_net_1683 ) , 
    .p1664 ( optlc_net_1684 ) , .p1665 ( optlc_net_1685 ) , 
    .p1666 ( optlc_net_1686 ) , .p1667 ( optlc_net_1687 ) , 
    .p1668 ( optlc_net_1688 ) , .p1669 ( optlc_net_1689 ) , 
    .p1670 ( optlc_net_1690 ) , .p1671 ( optlc_net_1691 ) , 
    .p1672 ( optlc_net_1692 ) , .p1673 ( optlc_net_1693 ) , 
    .p1674 ( optlc_net_1694 ) , .p1675 ( optlc_net_1695 ) , 
    .p1676 ( optlc_net_1696 ) , .p1677 ( optlc_net_1697 ) , 
    .p1678 ( optlc_net_1698 ) , .p1679 ( optlc_net_1699 ) , 
    .p1680 ( optlc_net_1700 ) , .p1681 ( optlc_net_1701 ) , 
    .p1682 ( optlc_net_1702 ) , .p1683 ( optlc_net_1703 ) , 
    .p1684 ( optlc_net_1704 ) , .p1685 ( optlc_net_1705 ) , 
    .p1686 ( optlc_net_1706 ) , .p1687 ( optlc_net_1707 ) , 
    .p1688 ( optlc_net_1708 ) , .p1689 ( optlc_net_1709 ) , 
    .p1690 ( optlc_net_1710 ) , .p1691 ( optlc_net_1711 ) , 
    .p1692 ( optlc_net_1712 ) , .p1693 ( optlc_net_1713 ) , 
    .p1694 ( optlc_net_1714 ) , .p1695 ( optlc_net_1715 ) , 
    .p1696 ( optlc_net_1716 ) , .p1697 ( optlc_net_1717 ) , 
    .p1698 ( optlc_net_1718 ) , .p1699 ( optlc_net_1719 ) , 
    .p1700 ( optlc_net_1720 ) , .p1701 ( optlc_net_1721 ) , 
    .p1702 ( optlc_net_1722 ) , .p1703 ( optlc_net_1723 ) , 
    .p1704 ( optlc_net_1724 ) , .p1705 ( optlc_net_1725 ) , 
    .p1706 ( optlc_net_1726 ) , .p1707 ( optlc_net_1727 ) , 
    .p1708 ( optlc_net_1728 ) , .p1709 ( optlc_net_1729 ) , 
    .p1710 ( optlc_net_1730 ) , .p1711 ( optlc_net_1731 ) , 
    .p1712 ( optlc_net_1732 ) , .p1713 ( optlc_net_1733 ) , 
    .p1714 ( optlc_net_1734 ) , .p1715 ( optlc_net_1735 ) , 
    .p1716 ( optlc_net_1736 ) , .p1717 ( optlc_net_1737 ) , 
    .p1718 ( optlc_net_1738 ) , .p1719 ( optlc_net_1739 ) , 
    .p1720 ( optlc_net_1740 ) , .p1721 ( optlc_net_1741 ) , 
    .p1722 ( optlc_net_1742 ) , .p1723 ( optlc_net_1743 ) , 
    .p1724 ( optlc_net_1744 ) , .p1725 ( optlc_net_1745 ) , 
    .p1726 ( optlc_net_1746 ) , .p1727 ( optlc_net_1747 ) , 
    .p1728 ( optlc_net_1748 ) , .p1729 ( optlc_net_1749 ) , 
    .p1730 ( optlc_net_1750 ) , .p1731 ( optlc_net_1751 ) , 
    .p1732 ( optlc_net_1752 ) , .p1733 ( optlc_net_1753 ) , 
    .p1734 ( optlc_net_1754 ) , .p1735 ( optlc_net_1755 ) , 
    .p1736 ( optlc_net_1756 ) , .p1737 ( optlc_net_1757 ) , 
    .p1738 ( optlc_net_1758 ) , .p1739 ( optlc_net_1759 ) , 
    .p1740 ( optlc_net_1760 ) , .p1741 ( optlc_net_1761 ) , 
    .p1742 ( optlc_net_1762 ) , .p1743 ( optlc_net_1763 ) , 
    .p1744 ( optlc_net_1764 ) , .p1745 ( optlc_net_1765 ) , 
    .p1746 ( optlc_net_1766 ) , .p1747 ( optlc_net_1767 ) , 
    .p1748 ( optlc_net_1768 ) , .p1749 ( optlc_net_1769 ) , 
    .p1750 ( optlc_net_1770 ) , .p1751 ( optlc_net_1771 ) , 
    .p1752 ( optlc_net_1772 ) , .p1753 ( optlc_net_1773 ) , 
    .p1754 ( optlc_net_1774 ) , .p1755 ( optlc_net_1775 ) , 
    .p1756 ( optlc_net_1776 ) , .p1757 ( optlc_net_1777 ) , 
    .p1758 ( optlc_net_1778 ) , .p1759 ( optlc_net_1779 ) , 
    .p1760 ( optlc_net_1780 ) , .p1761 ( optlc_net_1781 ) , 
    .p1762 ( optlc_net_1782 ) , .p1763 ( optlc_net_1783 ) , 
    .p1764 ( optlc_net_1784 ) , .p1765 ( optlc_net_1785 ) , 
    .p1766 ( optlc_net_1786 ) , .p1767 ( optlc_net_1787 ) , 
    .p1768 ( optlc_net_1788 ) , .p1769 ( optlc_net_1789 ) , 
    .p1770 ( optlc_net_1790 ) , .p1771 ( optlc_net_1791 ) , 
    .p1772 ( optlc_net_1792 ) , .p1773 ( optlc_net_1793 ) , 
    .p1774 ( optlc_net_1794 ) , .p1775 ( optlc_net_1795 ) , 
    .p1776 ( optlc_net_1796 ) , .p1777 ( optlc_net_1797 ) , 
    .p1778 ( optlc_net_1798 ) , .p1779 ( optlc_net_1799 ) , 
    .p1780 ( optlc_net_1800 ) , .p1781 ( optlc_net_1801 ) , 
    .p1782 ( optlc_net_1802 ) , .p1783 ( optlc_net_1803 ) , 
    .p1784 ( optlc_net_1804 ) , .p1785 ( optlc_net_1805 ) , 
    .p1786 ( optlc_net_1806 ) , .p1787 ( optlc_net_1807 ) , 
    .p1788 ( optlc_net_1808 ) , .p1789 ( optlc_net_1809 ) , 
    .p1790 ( optlc_net_1810 ) , .p1791 ( optlc_net_1811 ) , 
    .p1792 ( optlc_net_1812 ) , .p1793 ( optlc_net_1813 ) , 
    .p1794 ( optlc_net_1814 ) , .p1795 ( optlc_net_1815 ) , 
    .p1796 ( optlc_net_1816 ) , .p1797 ( optlc_net_1817 ) , 
    .p1798 ( optlc_net_1818 ) , .p1799 ( optlc_net_1819 ) , 
    .p1800 ( optlc_net_1820 ) , .p1801 ( optlc_net_1821 ) , 
    .p1802 ( optlc_net_1822 ) , .p1803 ( optlc_net_1823 ) , 
    .p1804 ( optlc_net_1824 ) , .p1805 ( optlc_net_1825 ) , 
    .p1806 ( optlc_net_1826 ) , .p1807 ( optlc_net_1827 ) , 
    .p1808 ( optlc_net_1828 ) , .p1809 ( optlc_net_1829 ) , 
    .p1810 ( optlc_net_1830 ) , .p1811 ( optlc_net_1831 ) , 
    .p1812 ( optlc_net_1832 ) , .p1813 ( optlc_net_1833 ) , 
    .p1814 ( optlc_net_1834 ) , .p1815 ( optlc_net_1835 ) , 
    .p1816 ( optlc_net_1836 ) , .p1817 ( optlc_net_1837 ) , 
    .p1818 ( optlc_net_1838 ) , .p1819 ( optlc_net_1839 ) , 
    .p1820 ( optlc_net_1840 ) , .p1821 ( optlc_net_1841 ) , 
    .p1822 ( optlc_net_1842 ) , .p1823 ( optlc_net_1843 ) , 
    .p1824 ( optlc_net_1844 ) , .p1825 ( optlc_net_1845 ) , 
    .p1826 ( optlc_net_1846 ) , .p1827 ( optlc_net_1847 ) , 
    .p1828 ( optlc_net_1848 ) , .p1829 ( optlc_net_1849 ) , 
    .p1830 ( optlc_net_1850 ) , .p1831 ( optlc_net_1851 ) , 
    .p1832 ( optlc_net_1852 ) , .p1833 ( optlc_net_1853 ) , 
    .p1834 ( optlc_net_1854 ) , .p1835 ( optlc_net_1855 ) , 
    .p1836 ( optlc_net_1856 ) , .p1837 ( optlc_net_1857 ) , 
    .p1838 ( optlc_net_1858 ) , .p1839 ( optlc_net_1859 ) , 
    .p1840 ( optlc_net_1860 ) , .p1841 ( optlc_net_1861 ) , 
    .p1842 ( optlc_net_1862 ) , .p1843 ( optlc_net_1863 ) , 
    .p1844 ( optlc_net_1864 ) , .p1845 ( optlc_net_1865 ) , 
    .p1846 ( optlc_net_1866 ) , .p1847 ( optlc_net_1867 ) , 
    .p1848 ( optlc_net_1868 ) , .p1849 ( optlc_net_1869 ) , 
    .p1850 ( optlc_net_1870 ) , .p1851 ( optlc_net_1871 ) , 
    .p1852 ( optlc_net_1872 ) , .p1853 ( optlc_net_1873 ) , 
    .p1854 ( optlc_net_1874 ) , .p1855 ( optlc_net_1875 ) , 
    .p1856 ( optlc_net_1876 ) , .p1857 ( optlc_net_1877 ) , 
    .p1858 ( optlc_net_1878 ) , .p1859 ( optlc_net_1879 ) , 
    .p1860 ( optlc_net_1880 ) , .p1861 ( optlc_net_1881 ) , 
    .p1862 ( optlc_net_1882 ) , .p1863 ( optlc_net_1883 ) , 
    .p1864 ( optlc_net_1884 ) , .p1865 ( optlc_net_1885 ) , 
    .p1866 ( optlc_net_1886 ) , .p1867 ( optlc_net_1887 ) , 
    .p1868 ( optlc_net_1888 ) , .p1869 ( optlc_net_1889 ) , 
    .p1870 ( optlc_net_1890 ) , .p1871 ( optlc_net_1891 ) , 
    .p1872 ( optlc_net_1892 ) , .p1873 ( optlc_net_1893 ) , 
    .p1874 ( optlc_net_1894 ) , .p1875 ( optlc_net_1895 ) , 
    .p1876 ( optlc_net_1896 ) , .p1877 ( optlc_net_1897 ) , 
    .p1878 ( optlc_net_1898 ) , .p1879 ( optlc_net_1899 ) , 
    .p1880 ( optlc_net_1900 ) , .p1881 ( optlc_net_1901 ) , 
    .p1882 ( optlc_net_1902 ) , .p1883 ( optlc_net_1903 ) , 
    .p1884 ( optlc_net_1904 ) , .p1885 ( optlc_net_1905 ) , 
    .p1886 ( optlc_net_1906 ) , .p1887 ( optlc_net_1907 ) , 
    .p1888 ( optlc_net_1908 ) , .p1889 ( optlc_net_1909 ) , 
    .p1890 ( optlc_net_1910 ) , .p1891 ( optlc_net_1911 ) , 
    .p1892 ( optlc_net_1912 ) , .p1893 ( optlc_net_1913 ) , 
    .p1894 ( optlc_net_1914 ) , .p1895 ( optlc_net_1915 ) , 
    .p1896 ( optlc_net_1916 ) , .p1897 ( optlc_net_1917 ) , 
    .p1898 ( optlc_net_1918 ) , .p1899 ( optlc_net_1919 ) , 
    .p1900 ( optlc_net_1920 ) , .p1901 ( optlc_net_1921 ) , 
    .p1902 ( optlc_net_1922 ) , .p1903 ( optlc_net_1923 ) , 
    .p1904 ( optlc_net_1924 ) , .p1905 ( optlc_net_1925 ) , 
    .p1906 ( optlc_net_1926 ) , .p1907 ( optlc_net_1927 ) , 
    .p1908 ( optlc_net_1928 ) , .p1909 ( optlc_net_1929 ) , 
    .p1910 ( optlc_net_1930 ) , .p1911 ( optlc_net_1931 ) , 
    .p1912 ( optlc_net_1932 ) , .p1913 ( optlc_net_1933 ) , 
    .p1914 ( optlc_net_1934 ) , .p1915 ( optlc_net_1935 ) , 
    .p1916 ( optlc_net_1936 ) , .p1917 ( optlc_net_1937 ) , 
    .p1918 ( optlc_net_1938 ) , .p1919 ( optlc_net_1939 ) , 
    .p1920 ( optlc_net_1940 ) , .p1921 ( optlc_net_1941 ) , 
    .p1922 ( optlc_net_1942 ) , .p1923 ( optlc_net_1943 ) , 
    .p1924 ( optlc_net_1944 ) , .p1925 ( optlc_net_1945 ) , 
    .p1926 ( optlc_net_1946 ) , .p1927 ( optlc_net_1947 ) , 
    .p1928 ( optlc_net_1948 ) , .p1929 ( optlc_net_1949 ) , 
    .p1930 ( optlc_net_1950 ) , .p1931 ( optlc_net_1951 ) , 
    .p1932 ( optlc_net_1952 ) , .p1933 ( optlc_net_1953 ) , 
    .p1934 ( optlc_net_1954 ) , .p1935 ( optlc_net_1955 ) , 
    .p1936 ( optlc_net_1956 ) , .p1937 ( optlc_net_1957 ) , 
    .p1938 ( optlc_net_1958 ) , .p1939 ( optlc_net_1959 ) , 
    .p1940 ( optlc_net_1960 ) , .p1941 ( optlc_net_1961 ) , 
    .p1942 ( optlc_net_1962 ) , .p1943 ( optlc_net_1963 ) , 
    .p1944 ( optlc_net_1964 ) , .p1945 ( optlc_net_1965 ) , 
    .p1946 ( optlc_net_1966 ) , .p1947 ( optlc_net_1967 ) , 
    .p1948 ( optlc_net_1968 ) , .p1949 ( optlc_net_1969 ) , 
    .p1950 ( optlc_net_1970 ) , .p1951 ( optlc_net_1971 ) , 
    .p1952 ( optlc_net_1972 ) , .p1953 ( optlc_net_1973 ) , 
    .p1954 ( optlc_net_1974 ) , .p1955 ( optlc_net_1975 ) , 
    .p1956 ( optlc_net_1976 ) , .p1957 ( optlc_net_1977 ) , 
    .p1958 ( optlc_net_1978 ) , .p1959 ( optlc_net_1979 ) , 
    .p1960 ( optlc_net_1980 ) , .p1961 ( optlc_net_1981 ) , 
    .p1962 ( optlc_net_1982 ) , .p1963 ( optlc_net_1983 ) , 
    .p1964 ( optlc_net_1984 ) , .p1965 ( optlc_net_1985 ) , 
    .p1966 ( optlc_net_1986 ) , .p1967 ( optlc_net_1987 ) , 
    .p1968 ( optlc_net_1988 ) , .p1969 ( optlc_net_1989 ) , 
    .p1970 ( optlc_net_1990 ) , .p1971 ( optlc_net_1991 ) , 
    .p1972 ( optlc_net_1992 ) , .p1973 ( optlc_net_1993 ) , 
    .p1974 ( optlc_net_1994 ) , .p1975 ( optlc_net_1995 ) , 
    .p1976 ( optlc_net_1996 ) , .p1977 ( optlc_net_1997 ) , 
    .p1978 ( optlc_net_1998 ) , .p1979 ( optlc_net_1999 ) , 
    .p1980 ( optlc_net_2000 ) , .p1981 ( optlc_net_2001 ) , 
    .p1982 ( optlc_net_2002 ) , .p1983 ( optlc_net_2003 ) , 
    .p1984 ( optlc_net_2004 ) , .p1985 ( optlc_net_2005 ) , 
    .p1986 ( optlc_net_2006 ) , .p1987 ( optlc_net_2007 ) , 
    .p1988 ( optlc_net_2008 ) , .p1989 ( optlc_net_2009 ) , 
    .p1990 ( optlc_net_2010 ) , .p1991 ( optlc_net_2011 ) , 
    .p1992 ( optlc_net_2012 ) , .p1993 ( optlc_net_2013 ) , 
    .p1994 ( optlc_net_2014 ) , .p1995 ( optlc_net_2015 ) , 
    .p1996 ( optlc_net_2016 ) , .p1997 ( optlc_net_2017 ) , 
    .p1998 ( optlc_net_2018 ) , .p1999 ( optlc_net_2019 ) , 
    .p2000 ( optlc_net_2020 ) , .p2001 ( optlc_net_2021 ) , 
    .p2002 ( optlc_net_2022 ) , .p2003 ( optlc_net_2023 ) , 
    .p2004 ( optlc_net_2024 ) , .p2005 ( optlc_net_2025 ) , 
    .p2006 ( optlc_net_2026 ) , .p2007 ( optlc_net_2027 ) , 
    .p2008 ( optlc_net_2028 ) , .p2009 ( optlc_net_2029 ) , 
    .p2010 ( optlc_net_2030 ) , .p2011 ( optlc_net_2031 ) , 
    .p2012 ( optlc_net_2032 ) , .p2013 ( optlc_net_2033 ) , 
    .p2014 ( optlc_net_2034 ) , .p2015 ( optlc_net_2035 ) , 
    .p2016 ( optlc_net_2036 ) , .p2017 ( optlc_net_2037 ) , 
    .p2018 ( optlc_net_2038 ) , .p2019 ( optlc_net_2039 ) , 
    .p2020 ( optlc_net_2040 ) , .p2021 ( optlc_net_2041 ) , 
    .p2022 ( optlc_net_2042 ) , .p2023 ( optlc_net_2043 ) , 
    .p2024 ( optlc_net_2044 ) , .p2025 ( optlc_net_2045 ) , 
    .p2026 ( optlc_net_2046 ) , .p2027 ( optlc_net_2047 ) , 
    .p2028 ( optlc_net_2048 ) , .p2029 ( optlc_net_2049 ) , 
    .p2030 ( optlc_net_2050 ) , .p2031 ( optlc_net_2051 ) , 
    .p2032 ( optlc_net_2052 ) , .p2033 ( optlc_net_2053 ) , 
    .p2034 ( optlc_net_2054 ) , .p2035 ( optlc_net_2055 ) , 
    .p2036 ( optlc_net_2056 ) , .p2037 ( optlc_net_2057 ) , 
    .p2038 ( optlc_net_2058 ) , .p2039 ( optlc_net_2059 ) , 
    .p2040 ( optlc_net_2060 ) , .p2041 ( optlc_net_2061 ) , 
    .p2042 ( optlc_net_2062 ) , .p2043 ( optlc_net_2063 ) , 
    .p2044 ( optlc_net_2064 ) , .p2045 ( optlc_net_2065 ) , 
    .p2046 ( optlc_net_2066 ) , .p2047 ( optlc_net_2067 ) , 
    .p2048 ( optlc_net_2068 ) , .p2049 ( optlc_net_2069 ) , 
    .p2050 ( optlc_net_2070 ) , .p2051 ( optlc_net_2071 ) , 
    .p2052 ( optlc_net_2072 ) , .p2053 ( optlc_net_2073 ) , 
    .p2054 ( optlc_net_2074 ) , .p2055 ( optlc_net_2075 ) , 
    .p2056 ( optlc_net_2076 ) , .p2057 ( optlc_net_2077 ) , 
    .p2058 ( optlc_net_2078 ) , .p2059 ( optlc_net_2079 ) , 
    .p2060 ( optlc_net_2080 ) , .p2061 ( optlc_net_2081 ) , 
    .p2062 ( optlc_net_2082 ) , .p2063 ( optlc_net_2083 ) , 
    .p2064 ( optlc_net_2084 ) , .p2065 ( optlc_net_2085 ) , 
    .p2066 ( optlc_net_2086 ) , .p2067 ( optlc_net_2087 ) , 
    .p2068 ( optlc_net_2088 ) , .p2069 ( optlc_net_2089 ) , 
    .p2070 ( optlc_net_2090 ) , .p2071 ( optlc_net_2091 ) , 
    .p2072 ( optlc_net_2092 ) , .p2073 ( optlc_net_2093 ) , 
    .p2074 ( optlc_net_2094 ) , .p2075 ( optlc_net_2095 ) , 
    .p2076 ( optlc_net_2096 ) , .p2077 ( optlc_net_2097 ) , 
    .p2078 ( optlc_net_2098 ) , .p2079 ( optlc_net_2099 ) , 
    .p2080 ( optlc_net_2100 ) , .p2081 ( optlc_net_2101 ) , 
    .p2082 ( optlc_net_2102 ) , .p2083 ( optlc_net_2103 ) , 
    .p2084 ( optlc_net_2104 ) , .p2085 ( optlc_net_2105 ) , 
    .p2086 ( optlc_net_2106 ) , .p2087 ( optlc_net_2107 ) , 
    .p2088 ( optlc_net_2108 ) , .p2089 ( optlc_net_2109 ) , 
    .p2090 ( optlc_net_2110 ) , .p2091 ( optlc_net_2111 ) , 
    .p2092 ( optlc_net_2112 ) , .p2093 ( optlc_net_2113 ) , 
    .p2094 ( optlc_net_2114 ) , .p2095 ( optlc_net_2115 ) , 
    .p2096 ( optlc_net_2116 ) , .p2097 ( optlc_net_2117 ) , 
    .p2098 ( optlc_net_2118 ) , .p2099 ( optlc_net_2119 ) , 
    .p2100 ( optlc_net_2120 ) , .p2101 ( optlc_net_2121 ) , 
    .p2102 ( optlc_net_2122 ) , .p2103 ( optlc_net_2123 ) , 
    .p2104 ( optlc_net_2124 ) , .p2105 ( optlc_net_2125 ) , 
    .p2106 ( optlc_net_2126 ) , .p2107 ( optlc_net_2127 ) , 
    .p2108 ( optlc_net_2128 ) , .p2109 ( optlc_net_2129 ) , 
    .p2110 ( optlc_net_2130 ) , .p2111 ( optlc_net_2131 ) , 
    .p2112 ( optlc_net_2132 ) , .p2113 ( optlc_net_2133 ) , 
    .p2114 ( optlc_net_2134 ) , .p2115 ( optlc_net_2135 ) , 
    .p2116 ( optlc_net_2136 ) , .p2117 ( optlc_net_2137 ) , 
    .p2118 ( optlc_net_2138 ) , .p2119 ( optlc_net_2139 ) , 
    .p2120 ( optlc_net_2140 ) , .p2121 ( optlc_net_2141 ) , 
    .p2122 ( optlc_net_2142 ) , .p2123 ( optlc_net_2143 ) , 
    .p2124 ( optlc_net_2144 ) , .p2125 ( optlc_net_2145 ) , 
    .p2126 ( optlc_net_2146 ) , .p2127 ( optlc_net_2147 ) , 
    .p2128 ( optlc_net_2148 ) , .p2129 ( optlc_net_2149 ) , 
    .p2130 ( optlc_net_2150 ) , .p2131 ( optlc_net_2151 ) , 
    .p2132 ( optlc_net_2152 ) , .p2133 ( optlc_net_2153 ) , 
    .p2134 ( optlc_net_2154 ) , .p2135 ( optlc_net_2155 ) , 
    .p2136 ( optlc_net_2156 ) , .p2137 ( optlc_net_2157 ) , 
    .p2138 ( optlc_net_2158 ) , .p2139 ( optlc_net_2159 ) , 
    .p2140 ( optlc_net_2160 ) , .p2141 ( optlc_net_2161 ) , 
    .p2142 ( optlc_net_2162 ) , .p2143 ( optlc_net_2163 ) , 
    .p2144 ( optlc_net_2164 ) , .p2145 ( optlc_net_2165 ) , 
    .p2146 ( optlc_net_2166 ) , .p2147 ( optlc_net_2167 ) , 
    .p2148 ( optlc_net_2168 ) , .p2149 ( optlc_net_2169 ) , 
    .p2150 ( optlc_net_2170 ) , .p2151 ( optlc_net_2171 ) , 
    .p2152 ( optlc_net_2172 ) , .p2153 ( optlc_net_2173 ) , 
    .p2154 ( optlc_net_2174 ) , .p2155 ( optlc_net_2175 ) , 
    .p2156 ( optlc_net_2176 ) , .p2157 ( optlc_net_2177 ) , 
    .p2158 ( optlc_net_2178 ) , .p2159 ( optlc_net_2179 ) , 
    .p2160 ( optlc_net_2180 ) , .p2161 ( optlc_net_2181 ) , 
    .p2162 ( optlc_net_2182 ) , .p2163 ( optlc_net_2183 ) , 
    .p2164 ( optlc_net_2184 ) , .p2165 ( optlc_net_2185 ) , 
    .p2166 ( optlc_net_2186 ) , .p2167 ( optlc_net_2187 ) , 
    .p2168 ( optlc_net_2188 ) , .p2169 ( optlc_net_2189 ) , 
    .p2170 ( optlc_net_2190 ) , .p2171 ( optlc_net_2191 ) , 
    .p2172 ( optlc_net_2192 ) , .p2173 ( optlc_net_2193 ) , 
    .p2174 ( optlc_net_2194 ) , .p2175 ( optlc_net_2195 ) , 
    .p2176 ( optlc_net_2196 ) , .p2177 ( optlc_net_2197 ) , 
    .p2178 ( optlc_net_2198 ) , .p2179 ( optlc_net_2199 ) , 
    .p2180 ( optlc_net_2200 ) , .p2181 ( optlc_net_2201 ) , 
    .p2182 ( optlc_net_2202 ) , .p2183 ( optlc_net_2203 ) , 
    .p2184 ( optlc_net_2204 ) , .p2185 ( optlc_net_2205 ) , 
    .p2186 ( optlc_net_2206 ) , .p2187 ( optlc_net_2207 ) , 
    .p2188 ( optlc_net_2208 ) , .p2189 ( optlc_net_2209 ) , 
    .p2190 ( optlc_net_2210 ) , .p2191 ( optlc_net_2211 ) , 
    .p2192 ( optlc_net_2212 ) , .p2193 ( optlc_net_2213 ) , 
    .p2194 ( optlc_net_2214 ) , .p2195 ( optlc_net_2215 ) , 
    .p2196 ( optlc_net_2216 ) , .p2197 ( optlc_net_2217 ) , 
    .p2198 ( optlc_net_2218 ) , .p2199 ( optlc_net_2219 ) , 
    .p2200 ( optlc_net_2220 ) , .p2201 ( optlc_net_2221 ) , 
    .p2202 ( optlc_net_2222 ) , .p2203 ( optlc_net_2223 ) , 
    .p2204 ( optlc_net_2224 ) , .p2205 ( optlc_net_2225 ) , 
    .p2206 ( optlc_net_2226 ) , .p2207 ( optlc_net_2227 ) , 
    .p2208 ( optlc_net_2228 ) , .p2209 ( optlc_net_2229 ) , 
    .p2210 ( optlc_net_2230 ) , .p2211 ( optlc_net_2231 ) , 
    .p2212 ( optlc_net_2232 ) , .p2213 ( optlc_net_2233 ) , 
    .p2214 ( optlc_net_2234 ) , .p2215 ( optlc_net_2235 ) , 
    .p2216 ( optlc_net_2236 ) , .p2217 ( optlc_net_2237 ) , 
    .p2218 ( optlc_net_2238 ) , .p2219 ( optlc_net_2239 ) , 
    .p2220 ( optlc_net_2240 ) , .p2221 ( optlc_net_2241 ) , 
    .p2222 ( optlc_net_2242 ) , .p2223 ( optlc_net_2243 ) , 
    .p2224 ( optlc_net_2244 ) , .p2225 ( optlc_net_2245 ) , 
    .p2226 ( optlc_net_2246 ) , .p2227 ( optlc_net_2247 ) , 
    .p2228 ( optlc_net_2248 ) , .p2229 ( optlc_net_2249 ) , 
    .p2230 ( optlc_net_2250 ) , .p2231 ( optlc_net_2251 ) , 
    .p2232 ( optlc_net_2252 ) , .p2233 ( optlc_net_2253 ) , 
    .p2234 ( optlc_net_2254 ) , .p2235 ( optlc_net_2255 ) , 
    .p2236 ( optlc_net_2256 ) , .p2237 ( optlc_net_2257 ) , 
    .p2238 ( optlc_net_2258 ) , .p2239 ( optlc_net_2259 ) , 
    .p2240 ( optlc_net_2260 ) , .p2241 ( optlc_net_2261 ) , 
    .p2242 ( optlc_net_2262 ) , .p2243 ( optlc_net_2263 ) , 
    .p2244 ( optlc_net_2264 ) , .p2245 ( optlc_net_2265 ) , 
    .p2246 ( optlc_net_2266 ) , .p2247 ( optlc_net_2267 ) , 
    .p2248 ( optlc_net_2268 ) , .p2249 ( optlc_net_2269 ) , 
    .p2250 ( optlc_net_2270 ) , .p2251 ( optlc_net_2271 ) , 
    .p2252 ( optlc_net_2272 ) , .p2253 ( optlc_net_2273 ) , 
    .p2254 ( optlc_net_2274 ) , .p2255 ( optlc_net_2275 ) , 
    .p2256 ( optlc_net_2276 ) , .p2257 ( optlc_net_2277 ) , 
    .p2258 ( optlc_net_2278 ) , .p2259 ( optlc_net_2279 ) , 
    .p2260 ( optlc_net_2280 ) , .p2261 ( optlc_net_2281 ) , 
    .p2262 ( optlc_net_2282 ) , .p2263 ( optlc_net_2283 ) , 
    .p2264 ( optlc_net_2284 ) , .p2265 ( optlc_net_2285 ) , 
    .p2266 ( optlc_net_2286 ) , .p2267 ( optlc_net_2287 ) , 
    .p2268 ( optlc_net_2288 ) , .p2269 ( optlc_net_2289 ) , 
    .p2270 ( optlc_net_2290 ) , .p2271 ( optlc_net_2291 ) , 
    .p2272 ( optlc_net_2292 ) , .p2273 ( optlc_net_2293 ) , 
    .p2274 ( optlc_net_2294 ) , .p2275 ( optlc_net_2295 ) , 
    .p2276 ( optlc_net_2296 ) , .p2277 ( optlc_net_2297 ) , 
    .p2278 ( optlc_net_2298 ) , .p2279 ( optlc_net_2299 ) , 
    .p2280 ( optlc_net_2300 ) , .p2281 ( optlc_net_2301 ) , 
    .p2282 ( optlc_net_2302 ) , .p2283 ( optlc_net_2303 ) , 
    .p2284 ( optlc_net_2304 ) , .p2285 ( optlc_net_2305 ) , 
    .p2286 ( optlc_net_2306 ) , .p2287 ( optlc_net_2307 ) , 
    .p2288 ( optlc_net_2308 ) , .p2289 ( optlc_net_2309 ) , 
    .p2290 ( optlc_net_2310 ) , .p2291 ( optlc_net_2311 ) , 
    .p2292 ( optlc_net_2312 ) , .p2293 ( optlc_net_2313 ) , 
    .p2294 ( optlc_net_2314 ) , .p2295 ( optlc_net_2315 ) , 
    .p2296 ( optlc_net_2316 ) , .p2297 ( optlc_net_2317 ) , 
    .p2298 ( optlc_net_2318 ) , .p2299 ( optlc_net_2319 ) , 
    .p2300 ( optlc_net_2320 ) , .p2301 ( optlc_net_2321 ) , 
    .p2302 ( optlc_net_2322 ) , .p2303 ( optlc_net_2323 ) , 
    .p2304 ( optlc_net_2324 ) , .p2305 ( optlc_net_2325 ) , 
    .p2306 ( optlc_net_2326 ) , .p2307 ( optlc_net_2327 ) , 
    .p2308 ( optlc_net_2328 ) , .p2309 ( optlc_net_2329 ) , 
    .p2310 ( optlc_net_2330 ) , .p2311 ( optlc_net_2331 ) , 
    .p2312 ( optlc_net_2332 ) , .p2313 ( optlc_net_2333 ) , 
    .p2314 ( optlc_net_2334 ) , .p2315 ( optlc_net_2335 ) , 
    .p2316 ( optlc_net_2336 ) , .p2317 ( optlc_net_2337 ) , 
    .p2318 ( optlc_net_2338 ) , .p2319 ( optlc_net_2339 ) , 
    .p2320 ( optlc_net_2340 ) , .p2321 ( optlc_net_2341 ) , 
    .p2322 ( optlc_net_2342 ) , .p2323 ( optlc_net_2343 ) , 
    .p2324 ( optlc_net_2344 ) , .p2325 ( optlc_net_2345 ) , 
    .p2326 ( optlc_net_2346 ) , .p2327 ( optlc_net_2347 ) , 
    .p2328 ( optlc_net_2348 ) , .p2329 ( optlc_net_2349 ) , 
    .p2330 ( optlc_net_2350 ) , .p2331 ( optlc_net_2351 ) , 
    .p2332 ( optlc_net_2352 ) , .p2333 ( optlc_net_2353 ) , 
    .p2334 ( optlc_net_2354 ) , .p2335 ( optlc_net_2355 ) , 
    .p2336 ( optlc_net_2356 ) , .p2337 ( optlc_net_2357 ) , 
    .p2338 ( optlc_net_2358 ) , .p2339 ( optlc_net_2359 ) , 
    .p2340 ( optlc_net_2360 ) , .p2341 ( optlc_net_2361 ) , 
    .p2342 ( optlc_net_2362 ) , .p2343 ( optlc_net_2363 ) , 
    .p2344 ( optlc_net_2364 ) , .p2345 ( optlc_net_2365 ) , 
    .p2346 ( optlc_net_2366 ) , .p2347 ( optlc_net_2367 ) , 
    .p2348 ( optlc_net_2368 ) , .p2349 ( optlc_net_2369 ) , 
    .p2350 ( optlc_net_2370 ) , .p2351 ( optlc_net_2371 ) , 
    .p2352 ( optlc_net_2372 ) , .p2353 ( optlc_net_2373 ) , 
    .p2354 ( optlc_net_2374 ) , .p2355 ( optlc_net_2375 ) , 
    .p2356 ( optlc_net_2376 ) , .p2357 ( optlc_net_2377 ) , 
    .p2358 ( optlc_net_2378 ) , .p2359 ( optlc_net_2379 ) , 
    .p2360 ( optlc_net_2380 ) , .p2361 ( optlc_net_2381 ) , 
    .p2362 ( optlc_net_2382 ) , .p2363 ( optlc_net_2383 ) , 
    .p2364 ( optlc_net_2384 ) , .p2365 ( optlc_net_2385 ) , 
    .p2366 ( optlc_net_2386 ) , .p2367 ( optlc_net_2387 ) , 
    .p2368 ( optlc_net_2388 ) , .p2369 ( optlc_net_2389 ) , 
    .p2370 ( optlc_net_2390 ) , .p2371 ( optlc_net_2391 ) , 
    .p2372 ( optlc_net_2392 ) , .p2373 ( optlc_net_2393 ) , 
    .p2374 ( optlc_net_2394 ) , .p2375 ( optlc_net_2395 ) , 
    .p2376 ( optlc_net_2396 ) , .p2377 ( optlc_net_2397 ) , 
    .p2378 ( optlc_net_2398 ) , .p2379 ( optlc_net_2399 ) , 
    .p2380 ( optlc_net_2400 ) , .p2381 ( optlc_net_2401 ) , 
    .p2382 ( optlc_net_2402 ) , .p2383 ( optlc_net_2403 ) , 
    .p2384 ( optlc_net_2404 ) , .p2385 ( optlc_net_2405 ) , 
    .p2386 ( optlc_net_2406 ) , .p2387 ( optlc_net_2407 ) , 
    .p2388 ( optlc_net_2408 ) , .p2389 ( optlc_net_2409 ) , 
    .p2390 ( optlc_net_2410 ) , .p2391 ( optlc_net_2411 ) , 
    .p2392 ( optlc_net_2412 ) , .p2393 ( optlc_net_2413 ) , 
    .p2394 ( optlc_net_2414 ) , .p2395 ( optlc_net_2415 ) , 
    .p2396 ( optlc_net_2416 ) , .p2397 ( optlc_net_2417 ) , 
    .p2398 ( optlc_net_2418 ) , .p2399 ( optlc_net_2419 ) , 
    .p2400 ( optlc_net_2420 ) , .p2401 ( optlc_net_2421 ) , 
    .p2402 ( optlc_net_2422 ) , .p2403 ( optlc_net_2423 ) , 
    .p2404 ( optlc_net_2424 ) , .p2405 ( optlc_net_2425 ) , 
    .p2406 ( optlc_net_2426 ) , .p2407 ( optlc_net_2427 ) , 
    .p2408 ( optlc_net_2428 ) , .p2409 ( optlc_net_2429 ) , 
    .p2410 ( optlc_net_2430 ) , .p2411 ( optlc_net_2431 ) , 
    .p2412 ( optlc_net_2432 ) , .p2413 ( optlc_net_2433 ) , 
    .p2414 ( optlc_net_2434 ) , .p2415 ( optlc_net_2435 ) , 
    .p2416 ( optlc_net_2436 ) , .p2417 ( optlc_net_2437 ) , 
    .p2418 ( optlc_net_2438 ) , .p2419 ( optlc_net_2439 ) , 
    .p2420 ( optlc_net_2440 ) , .p2421 ( optlc_net_2441 ) , 
    .p2422 ( optlc_net_2442 ) , .p2423 ( optlc_net_2443 ) , 
    .p2424 ( optlc_net_2444 ) , .p2425 ( optlc_net_2445 ) , 
    .p2426 ( optlc_net_2446 ) , .p2427 ( optlc_net_2447 ) , 
    .p2428 ( optlc_net_2448 ) , .p2429 ( optlc_net_2449 ) , 
    .p2430 ( optlc_net_2450 ) , .p2431 ( optlc_net_2451 ) , 
    .p2432 ( optlc_net_2452 ) , .p2433 ( optlc_net_2453 ) , 
    .p2434 ( optlc_net_2454 ) , .p2435 ( optlc_net_2455 ) , 
    .p2436 ( optlc_net_2456 ) , .p2437 ( optlc_net_2457 ) , 
    .p2438 ( optlc_net_2458 ) , .p2439 ( optlc_net_2459 ) , 
    .p2440 ( optlc_net_2460 ) , .p2441 ( optlc_net_2461 ) , 
    .p2442 ( optlc_net_2462 ) , .p2443 ( optlc_net_2463 ) , 
    .p2444 ( optlc_net_2464 ) , .p2445 ( optlc_net_2465 ) , 
    .p2446 ( optlc_net_2466 ) , .p2447 ( optlc_net_2467 ) , 
    .p2448 ( optlc_net_2468 ) , .p2449 ( optlc_net_2469 ) , 
    .p2450 ( optlc_net_2470 ) , .p2451 ( optlc_net_2471 ) , 
    .p2452 ( optlc_net_2472 ) , .p2453 ( optlc_net_2473 ) , 
    .p2454 ( optlc_net_2474 ) , .p2455 ( optlc_net_2475 ) , 
    .p2456 ( optlc_net_2476 ) , .p2457 ( optlc_net_2477 ) , 
    .p2458 ( optlc_net_2478 ) , .p2459 ( optlc_net_2479 ) , 
    .p2460 ( optlc_net_2480 ) , .p2461 ( optlc_net_2481 ) , 
    .p2462 ( optlc_net_2482 ) , .p2463 ( optlc_net_2483 ) , 
    .p2464 ( optlc_net_2484 ) , .p2465 ( optlc_net_2485 ) , 
    .p2466 ( optlc_net_2486 ) , .p2467 ( optlc_net_2487 ) , 
    .p2468 ( optlc_net_2488 ) , .p2469 ( optlc_net_2489 ) , 
    .p2470 ( optlc_net_2490 ) , .p2471 ( optlc_net_2491 ) , 
    .p2472 ( optlc_net_2492 ) , .p2473 ( optlc_net_2493 ) , 
    .p2474 ( optlc_net_2494 ) , .p2475 ( optlc_net_2495 ) , 
    .p2476 ( optlc_net_2496 ) , .p2477 ( optlc_net_2497 ) , 
    .p2478 ( optlc_net_2498 ) , .p2479 ( optlc_net_2499 ) , 
    .p2480 ( optlc_net_2500 ) , .p2481 ( optlc_net_2501 ) , 
    .p2482 ( optlc_net_2502 ) , .p2483 ( optlc_net_2503 ) , 
    .p2484 ( optlc_net_2504 ) , .p2485 ( optlc_net_2505 ) , 
    .p2486 ( optlc_net_2506 ) , .p2487 ( optlc_net_2507 ) , 
    .p2488 ( optlc_net_2508 ) , .p2489 ( optlc_net_2509 ) , 
    .p2490 ( optlc_net_2510 ) , .p2491 ( optlc_net_2511 ) , 
    .p2492 ( optlc_net_2512 ) , .p2493 ( optlc_net_2513 ) , 
    .p2494 ( optlc_net_2514 ) , .p2495 ( optlc_net_2515 ) , 
    .p2496 ( optlc_net_2516 ) , .p2497 ( optlc_net_2517 ) , 
    .p2498 ( optlc_net_2518 ) , .p2499 ( optlc_net_2519 ) , 
    .p2500 ( optlc_net_2520 ) , .p2501 ( optlc_net_2521 ) , 
    .p2502 ( optlc_net_2522 ) , .p2503 ( optlc_net_2523 ) , 
    .p2504 ( optlc_net_2524 ) , .p2505 ( optlc_net_2525 ) , 
    .p2506 ( optlc_net_2526 ) , .p2507 ( optlc_net_2527 ) , 
    .p2508 ( optlc_net_2528 ) , .p2509 ( optlc_net_2529 ) , 
    .p2510 ( optlc_net_2530 ) , .p2511 ( optlc_net_2531 ) , 
    .p2512 ( optlc_net_2532 ) , .p2513 ( optlc_net_2533 ) , 
    .p2514 ( optlc_net_2534 ) , .p2515 ( optlc_net_2535 ) , 
    .p2516 ( optlc_net_2536 ) , .p2517 ( optlc_net_2537 ) , 
    .p2518 ( optlc_net_2538 ) , .p2519 ( optlc_net_2539 ) , 
    .p2520 ( optlc_net_2540 ) , .p2521 ( optlc_net_2541 ) , 
    .p2522 ( optlc_net_2542 ) , .p2523 ( optlc_net_2543 ) , 
    .p2524 ( optlc_net_2544 ) , .p2525 ( optlc_net_2545 ) , 
    .p2526 ( optlc_net_2546 ) , .p2527 ( optlc_net_2547 ) , 
    .p2528 ( optlc_net_2548 ) , .p2529 ( optlc_net_2549 ) , 
    .p2530 ( optlc_net_2550 ) , .p2531 ( optlc_net_2551 ) , 
    .p2532 ( optlc_net_2552 ) , .p2533 ( optlc_net_2553 ) , 
    .p2534 ( optlc_net_2554 ) , .p2535 ( optlc_net_2555 ) , 
    .p2536 ( optlc_net_2556 ) , .p2537 ( optlc_net_2557 ) , 
    .p2538 ( optlc_net_2558 ) , .p2539 ( optlc_net_2559 ) , 
    .p2540 ( optlc_net_2560 ) , .p2541 ( optlc_net_2561 ) , 
    .p2542 ( optlc_net_2562 ) , .p2543 ( optlc_net_2563 ) , 
    .p2544 ( optlc_net_2564 ) , .p2545 ( optlc_net_2565 ) , 
    .p2546 ( optlc_net_2566 ) , .p2547 ( optlc_net_2567 ) , 
    .p2548 ( optlc_net_2568 ) , .p2549 ( optlc_net_2569 ) , 
    .p2550 ( optlc_net_2570 ) , .p2551 ( optlc_net_2571 ) , 
    .p2552 ( optlc_net_2572 ) , .p2553 ( optlc_net_2573 ) , 
    .p2554 ( optlc_net_2574 ) , .p2555 ( optlc_net_2575 ) , 
    .p2556 ( optlc_net_2576 ) , .p2557 ( optlc_net_2577 ) , 
    .p2558 ( optlc_net_2578 ) , .p2559 ( optlc_net_2579 ) , 
    .p2560 ( optlc_net_2580 ) , .p2561 ( optlc_net_2581 ) , 
    .p2562 ( optlc_net_2582 ) , .p2563 ( optlc_net_2583 ) , 
    .p2564 ( optlc_net_2584 ) , .p2565 ( optlc_net_2585 ) , 
    .p2566 ( optlc_net_2586 ) , .p2567 ( optlc_net_2587 ) , 
    .p2568 ( optlc_net_2588 ) , .p2569 ( optlc_net_2589 ) , 
    .p2570 ( optlc_net_2590 ) , .p2571 ( optlc_net_2591 ) , 
    .p2572 ( optlc_net_2592 ) , .p2573 ( optlc_net_2593 ) , 
    .p2574 ( optlc_net_2594 ) , .p2575 ( optlc_net_2595 ) , 
    .p2576 ( optlc_net_2596 ) , .p2577 ( optlc_net_2597 ) , 
    .p2578 ( optlc_net_2598 ) , .p2579 ( optlc_net_2599 ) , 
    .p2580 ( optlc_net_2600 ) , .p2581 ( optlc_net_2601 ) , 
    .p2582 ( optlc_net_2602 ) , .p2583 ( optlc_net_2603 ) , 
    .p2584 ( optlc_net_2604 ) , .p2585 ( optlc_net_2605 ) , 
    .p2586 ( optlc_net_2606 ) , .p2587 ( optlc_net_2607 ) , 
    .p2588 ( optlc_net_2608 ) , .p2589 ( optlc_net_2609 ) , 
    .p2590 ( optlc_net_2610 ) , .p2591 ( optlc_net_2611 ) , 
    .p2592 ( optlc_net_2612 ) , .p2593 ( optlc_net_2613 ) , 
    .p2594 ( optlc_net_2614 ) , .p2595 ( optlc_net_2615 ) , 
    .p2596 ( optlc_net_2616 ) , .p2597 ( optlc_net_2617 ) , 
    .p2598 ( optlc_net_2618 ) , .p2599 ( optlc_net_2619 ) , 
    .p2600 ( optlc_net_2620 ) , .p2601 ( optlc_net_2621 ) , 
    .p2602 ( optlc_net_2622 ) , .p2603 ( optlc_net_2623 ) , 
    .p2604 ( optlc_net_2624 ) , .p2605 ( optlc_net_2625 ) , 
    .p2606 ( optlc_net_2626 ) , .p2607 ( optlc_net_2627 ) , 
    .p2608 ( optlc_net_2628 ) , .p2609 ( optlc_net_2629 ) , 
    .p2610 ( optlc_net_2630 ) , .p2611 ( optlc_net_2631 ) , 
    .p2612 ( optlc_net_2632 ) , .p2613 ( optlc_net_2633 ) , 
    .p2614 ( optlc_net_2634 ) , .p2615 ( optlc_net_2635 ) , 
    .p2616 ( optlc_net_2636 ) , .p2617 ( optlc_net_2637 ) , 
    .p2618 ( optlc_net_2638 ) , .p2619 ( optlc_net_2639 ) , 
    .p2620 ( optlc_net_2640 ) , .p2621 ( optlc_net_2641 ) , 
    .p2622 ( optlc_net_2642 ) , .p2623 ( optlc_net_2643 ) , 
    .p2624 ( optlc_net_2644 ) , .p2625 ( optlc_net_2645 ) , 
    .p2626 ( optlc_net_2646 ) , .p2627 ( optlc_net_2647 ) , 
    .p2628 ( optlc_net_2648 ) , .p2629 ( optlc_net_2649 ) , 
    .p2630 ( optlc_net_2650 ) , .p2631 ( optlc_net_2651 ) , 
    .p2632 ( optlc_net_2652 ) , .p2633 ( optlc_net_2653 ) , 
    .p2634 ( optlc_net_2654 ) , .p2635 ( optlc_net_2655 ) , 
    .p2636 ( optlc_net_2656 ) , .p2637 ( optlc_net_2657 ) , 
    .p2638 ( optlc_net_2658 ) , .p2639 ( optlc_net_2659 ) , 
    .p2640 ( optlc_net_2660 ) , .p2641 ( optlc_net_2661 ) , 
    .p2642 ( optlc_net_2662 ) , .p2643 ( optlc_net_2663 ) , 
    .p2644 ( optlc_net_2664 ) , .p2645 ( optlc_net_2665 ) , 
    .p2646 ( optlc_net_2666 ) , .p2647 ( optlc_net_2667 ) , 
    .p2648 ( optlc_net_2668 ) , .p2649 ( optlc_net_2669 ) , 
    .p2650 ( optlc_net_2670 ) , .p2651 ( optlc_net_2671 ) , 
    .p2652 ( optlc_net_2672 ) , .p2653 ( optlc_net_2673 ) , 
    .p2654 ( optlc_net_2674 ) , .p2655 ( optlc_net_2675 ) , 
    .p2656 ( optlc_net_2676 ) , .p2657 ( optlc_net_2677 ) , 
    .p2658 ( optlc_net_2678 ) , .p2659 ( optlc_net_2679 ) , 
    .p2660 ( optlc_net_2680 ) , .p2661 ( optlc_net_2681 ) , 
    .p2662 ( optlc_net_2682 ) , .p2663 ( optlc_net_2683 ) , 
    .p2664 ( optlc_net_2684 ) , .p2665 ( optlc_net_2685 ) , 
    .p2666 ( optlc_net_2686 ) , .p2667 ( optlc_net_2687 ) , 
    .p2668 ( optlc_net_2688 ) , .p2669 ( optlc_net_2689 ) , 
    .p2670 ( optlc_net_2690 ) , .p2671 ( optlc_net_2691 ) , 
    .p2672 ( optlc_net_2692 ) , .p2673 ( optlc_net_2693 ) , 
    .p2674 ( optlc_net_2694 ) , .p2675 ( optlc_net_2695 ) , 
    .p2676 ( optlc_net_2696 ) , .p2677 ( optlc_net_2697 ) , 
    .p2678 ( optlc_net_2698 ) , .p2679 ( optlc_net_2699 ) , 
    .p2680 ( optlc_net_2700 ) , .p2681 ( optlc_net_2701 ) , 
    .p2682 ( optlc_net_2702 ) , .p2683 ( optlc_net_2703 ) , 
    .p2684 ( optlc_net_2704 ) , .p2685 ( optlc_net_2705 ) , 
    .p2686 ( optlc_net_2706 ) , .p2687 ( optlc_net_2707 ) , 
    .p2688 ( optlc_net_2708 ) , .p2689 ( optlc_net_2709 ) , 
    .p2690 ( optlc_net_2710 ) , .p2691 ( optlc_net_2711 ) , 
    .p2692 ( optlc_net_2712 ) , .p2693 ( optlc_net_2713 ) , 
    .p2694 ( optlc_net_2714 ) , .p2695 ( optlc_net_2715 ) , 
    .p2696 ( optlc_net_2716 ) , .p2697 ( optlc_net_2717 ) , 
    .p2698 ( optlc_net_2718 ) , .p2699 ( optlc_net_2719 ) , 
    .p2700 ( optlc_net_2720 ) , .p2701 ( optlc_net_2721 ) , 
    .p2702 ( optlc_net_2722 ) , .p2703 ( optlc_net_2723 ) , 
    .p2704 ( optlc_net_2724 ) , .p2705 ( optlc_net_2725 ) , 
    .p2706 ( optlc_net_2726 ) , .p2707 ( optlc_net_2727 ) , 
    .p2708 ( optlc_net_2728 ) , .p2709 ( optlc_net_2729 ) , 
    .p2710 ( optlc_net_2730 ) , .p2711 ( optlc_net_2731 ) , 
    .p2712 ( optlc_net_2732 ) , .p2713 ( optlc_net_2733 ) , 
    .p2714 ( optlc_net_2734 ) , .p2715 ( optlc_net_2735 ) , 
    .p2716 ( optlc_net_2736 ) , .p2717 ( optlc_net_2737 ) , 
    .p2718 ( optlc_net_2738 ) , .p2719 ( optlc_net_2739 ) , 
    .p2720 ( optlc_net_2740 ) , .p2721 ( optlc_net_2741 ) , 
    .p2722 ( optlc_net_2742 ) , .p2723 ( optlc_net_2743 ) , 
    .p2724 ( optlc_net_2744 ) , .p2725 ( optlc_net_2745 ) , 
    .p2726 ( optlc_net_2746 ) , .p2727 ( optlc_net_2747 ) , 
    .p2728 ( optlc_net_2748 ) , .p2729 ( optlc_net_2749 ) , 
    .p2730 ( optlc_net_2750 ) , .p2731 ( optlc_net_2751 ) , 
    .p2732 ( optlc_net_2752 ) , .p2733 ( optlc_net_2753 ) , 
    .p2734 ( optlc_net_2754 ) , .p2735 ( optlc_net_2755 ) , 
    .p2736 ( optlc_net_2756 ) , .p2737 ( optlc_net_2757 ) , 
    .p2738 ( optlc_net_2758 ) , .p2739 ( optlc_net_2759 ) , 
    .p2740 ( optlc_net_2760 ) , .p2741 ( optlc_net_2761 ) , 
    .p2742 ( optlc_net_2762 ) , .p2743 ( optlc_net_2763 ) , 
    .p2744 ( optlc_net_2764 ) , .p2745 ( optlc_net_2765 ) , 
    .p2746 ( optlc_net_2766 ) , .p2747 ( optlc_net_2767 ) , 
    .p2748 ( optlc_net_2768 ) , .p2749 ( optlc_net_2769 ) , 
    .p2750 ( optlc_net_2770 ) , .p2751 ( optlc_net_2771 ) , 
    .p2752 ( optlc_net_2772 ) , .p2753 ( optlc_net_2773 ) , 
    .p2754 ( optlc_net_2774 ) , .p2755 ( optlc_net_2775 ) , 
    .p2756 ( optlc_net_2776 ) , .p2757 ( optlc_net_2777 ) , 
    .p2758 ( optlc_net_2778 ) , .p2759 ( optlc_net_2779 ) , 
    .p2760 ( optlc_net_2780 ) , .p2761 ( optlc_net_2781 ) , 
    .p2762 ( optlc_net_2782 ) , .p2763 ( optlc_net_2783 ) , 
    .p2764 ( optlc_net_2784 ) , .p2765 ( optlc_net_2785 ) , 
    .p2766 ( optlc_net_2786 ) , .p2767 ( optlc_net_2787 ) , 
    .p2768 ( optlc_net_2788 ) , .p2769 ( optlc_net_2789 ) , 
    .p2770 ( optlc_net_2790 ) , .p2771 ( optlc_net_2791 ) , 
    .p2772 ( optlc_net_2792 ) , .p2773 ( optlc_net_2793 ) , 
    .p2774 ( optlc_net_2794 ) , .p2775 ( optlc_net_2795 ) , 
    .p2776 ( optlc_net_2796 ) , .p2777 ( optlc_net_2797 ) , 
    .p2778 ( optlc_net_2798 ) , .p2779 ( optlc_net_2799 ) , 
    .p2780 ( optlc_net_2800 ) , .p2781 ( optlc_net_2801 ) , 
    .p2782 ( optlc_net_2802 ) , .p2783 ( optlc_net_2803 ) , 
    .p2784 ( optlc_net_2804 ) , .p2785 ( optlc_net_2805 ) , 
    .p2786 ( optlc_net_2806 ) , .p2787 ( optlc_net_2807 ) , 
    .p2788 ( optlc_net_2808 ) , .p2789 ( optlc_net_2809 ) , 
    .p2790 ( optlc_net_2810 ) , .p2791 ( optlc_net_2811 ) , 
    .p2792 ( optlc_net_2812 ) , .p2793 ( optlc_net_2813 ) , 
    .p2794 ( optlc_net_2814 ) , .p2795 ( optlc_net_2815 ) , 
    .p2796 ( optlc_net_2816 ) , .p2797 ( optlc_net_2817 ) , 
    .p2798 ( optlc_net_2818 ) , .p2799 ( optlc_net_2819 ) , 
    .p2800 ( optlc_net_2820 ) , .p2801 ( optlc_net_2821 ) , 
    .p2802 ( optlc_net_2822 ) , .p2803 ( optlc_net_2823 ) , 
    .p2804 ( optlc_net_2824 ) , .p2805 ( optlc_net_2825 ) , 
    .p2806 ( optlc_net_2826 ) , .p2807 ( optlc_net_2827 ) , 
    .p2808 ( optlc_net_2828 ) , .p2809 ( optlc_net_2829 ) , 
    .p2810 ( optlc_net_2830 ) , .p2811 ( optlc_net_2831 ) , 
    .p2812 ( optlc_net_2832 ) , .p2813 ( optlc_net_2833 ) , 
    .p2814 ( optlc_net_2834 ) , .p2815 ( optlc_net_2835 ) , 
    .p2816 ( optlc_net_2836 ) , .p2817 ( optlc_net_2837 ) , 
    .p2818 ( optlc_net_2838 ) , .p2819 ( optlc_net_2839 ) , 
    .p2820 ( optlc_net_2840 ) , .p2821 ( optlc_net_2841 ) , 
    .p2822 ( optlc_net_2842 ) , .p2823 ( optlc_net_2843 ) , 
    .p2824 ( optlc_net_2844 ) , .p2825 ( optlc_net_2845 ) , 
    .p2826 ( optlc_net_2846 ) , .p2827 ( optlc_net_2847 ) , 
    .p2828 ( optlc_net_2848 ) , .p2829 ( optlc_net_2849 ) , 
    .p2830 ( optlc_net_2850 ) , .p2831 ( optlc_net_2851 ) , 
    .p2832 ( optlc_net_2852 ) , .p2833 ( optlc_net_2853 ) , 
    .p2834 ( optlc_net_2854 ) , .p2835 ( optlc_net_2855 ) , 
    .p2836 ( optlc_net_2856 ) , .p2837 ( optlc_net_2857 ) , 
    .p2838 ( optlc_net_2858 ) , .p2839 ( optlc_net_2859 ) , 
    .p2840 ( optlc_net_2860 ) , .p2841 ( optlc_net_2861 ) , 
    .p2842 ( optlc_net_2862 ) , .p2843 ( optlc_net_2863 ) , 
    .p2844 ( optlc_net_2864 ) , .p2845 ( optlc_net_2865 ) , 
    .p2846 ( optlc_net_2866 ) , .p2847 ( optlc_net_2867 ) , 
    .p2848 ( optlc_net_2868 ) , .p2849 ( optlc_net_2869 ) , 
    .p2850 ( optlc_net_2870 ) , .p2851 ( optlc_net_2871 ) , 
    .p2852 ( optlc_net_2872 ) , .p2853 ( optlc_net_2873 ) , 
    .p2854 ( optlc_net_2874 ) , .p2855 ( optlc_net_2875 ) , 
    .p2856 ( optlc_net_2876 ) , .p2857 ( optlc_net_2877 ) , 
    .p2858 ( optlc_net_2878 ) , .p2859 ( optlc_net_2879 ) , 
    .p2860 ( optlc_net_2880 ) , .p2861 ( optlc_net_2881 ) , 
    .p2862 ( optlc_net_2882 ) , .p2863 ( optlc_net_2883 ) , 
    .p2864 ( optlc_net_2884 ) , .p2865 ( optlc_net_2885 ) , 
    .p2866 ( optlc_net_2886 ) , .p2867 ( optlc_net_2887 ) , 
    .p2868 ( optlc_net_2888 ) , .p2869 ( optlc_net_2889 ) , 
    .p2870 ( optlc_net_2890 ) , .p2871 ( optlc_net_2891 ) , 
    .p2872 ( optlc_net_2892 ) , .p2873 ( optlc_net_2893 ) , 
    .p2874 ( optlc_net_2894 ) , .p2875 ( optlc_net_2895 ) , 
    .p2876 ( optlc_net_2896 ) , .p2877 ( optlc_net_2897 ) , 
    .p2878 ( optlc_net_2898 ) , .p2879 ( optlc_net_2899 ) , 
    .p2880 ( optlc_net_2900 ) , .p2881 ( optlc_net_2901 ) , 
    .p2882 ( optlc_net_2902 ) , .p2883 ( optlc_net_2903 ) , 
    .p2884 ( optlc_net_2904 ) , .p2885 ( optlc_net_2905 ) , 
    .p2886 ( optlc_net_2906 ) , .p2887 ( optlc_net_2907 ) , 
    .p2888 ( optlc_net_2908 ) , .p2889 ( optlc_net_2909 ) , 
    .p2890 ( optlc_net_2910 ) , .p2891 ( optlc_net_2911 ) , 
    .p2892 ( optlc_net_2912 ) , .p2893 ( optlc_net_2913 ) , 
    .p2894 ( optlc_net_2914 ) , .p2895 ( optlc_net_2915 ) , 
    .p2896 ( optlc_net_2916 ) , .p2897 ( optlc_net_2917 ) , 
    .p2898 ( optlc_net_2918 ) , .p2899 ( optlc_net_2919 ) , 
    .p2900 ( optlc_net_2920 ) , .p2901 ( optlc_net_2921 ) , 
    .p2902 ( optlc_net_2922 ) , .p2903 ( optlc_net_2923 ) , 
    .p2904 ( optlc_net_2924 ) , .p2905 ( optlc_net_2925 ) , 
    .p2906 ( optlc_net_2926 ) , .p2907 ( optlc_net_2927 ) , 
    .p2908 ( optlc_net_2928 ) , .p2909 ( optlc_net_2929 ) , 
    .p2910 ( optlc_net_2930 ) , .p2911 ( optlc_net_2931 ) , 
    .p2912 ( optlc_net_2932 ) , .p2913 ( optlc_net_2933 ) , 
    .p2914 ( optlc_net_2934 ) , .p2915 ( optlc_net_2935 ) , 
    .p2916 ( optlc_net_2936 ) , .p2917 ( optlc_net_2937 ) , 
    .p2918 ( optlc_net_2938 ) , .p2919 ( optlc_net_2939 ) , 
    .p2920 ( optlc_net_2940 ) , .p2921 ( optlc_net_2941 ) , 
    .p2922 ( optlc_net_2942 ) , .p2923 ( optlc_net_2943 ) , 
    .p2924 ( optlc_net_2944 ) , .p2925 ( optlc_net_2945 ) , 
    .p2926 ( optlc_net_2946 ) , .p2927 ( optlc_net_2947 ) , 
    .p2928 ( optlc_net_2948 ) , .p2929 ( optlc_net_2949 ) , 
    .p2930 ( optlc_net_2950 ) , .p2931 ( optlc_net_2951 ) , 
    .p2932 ( optlc_net_2952 ) , .p2933 ( optlc_net_2953 ) , 
    .p2934 ( optlc_net_2954 ) , .p2935 ( optlc_net_2955 ) , 
    .p2936 ( optlc_net_2956 ) , .p2937 ( optlc_net_2957 ) , 
    .p2938 ( optlc_net_2958 ) , .p2939 ( optlc_net_2959 ) , 
    .p2940 ( optlc_net_2960 ) , .p2941 ( optlc_net_2961 ) , 
    .p2942 ( optlc_net_2962 ) , .p2943 ( optlc_net_2963 ) , 
    .p2944 ( optlc_net_2964 ) , .p2945 ( optlc_net_2965 ) , 
    .p2946 ( optlc_net_2966 ) , .p2947 ( optlc_net_2967 ) , 
    .p2948 ( optlc_net_2968 ) , .p2949 ( optlc_net_2969 ) , 
    .p2950 ( optlc_net_2970 ) , .p2951 ( optlc_net_2971 ) , 
    .p2952 ( optlc_net_2972 ) , .p2953 ( optlc_net_2973 ) , 
    .p2954 ( optlc_net_2974 ) , .p2955 ( optlc_net_2975 ) , 
    .p2956 ( optlc_net_2976 ) , .p2957 ( optlc_net_2977 ) , 
    .p2958 ( optlc_net_2978 ) , .p2959 ( optlc_net_2979 ) , 
    .p2960 ( optlc_net_2980 ) , .p2961 ( optlc_net_2981 ) , 
    .p2962 ( optlc_net_2982 ) , .p2963 ( optlc_net_2983 ) , 
    .p2964 ( optlc_net_2984 ) , .p2965 ( optlc_net_2985 ) , 
    .p2966 ( optlc_net_2986 ) , .p2967 ( optlc_net_2987 ) , 
    .p2968 ( optlc_net_2988 ) , .p2969 ( optlc_net_2989 ) , 
    .p2970 ( optlc_net_2990 ) , .p2971 ( optlc_net_2991 ) , 
    .p2972 ( optlc_net_2992 ) , .p2973 ( optlc_net_2993 ) , 
    .p2974 ( optlc_net_2994 ) , .p2975 ( optlc_net_2995 ) , 
    .p2976 ( optlc_net_2996 ) , .p2977 ( optlc_net_2997 ) , 
    .p2978 ( optlc_net_2998 ) , .p2979 ( optlc_net_2999 ) , 
    .p2980 ( optlc_net_3000 ) , .p2981 ( optlc_net_3001 ) , 
    .p2982 ( optlc_net_3002 ) , .p2983 ( optlc_net_3003 ) , 
    .p2984 ( optlc_net_3004 ) , .p2985 ( optlc_net_3005 ) , 
    .p2986 ( optlc_net_3006 ) , .p2987 ( optlc_net_3007 ) , 
    .p2988 ( optlc_net_3008 ) , .p2989 ( optlc_net_3009 ) , 
    .p2990 ( optlc_net_3010 ) , .p2991 ( optlc_net_3011 ) , 
    .p2992 ( optlc_net_3012 ) , .p2993 ( optlc_net_3013 ) , 
    .p2994 ( optlc_net_3014 ) , .p2995 ( optlc_net_3015 ) , 
    .p2996 ( optlc_net_3016 ) , .p2997 ( optlc_net_3017 ) , 
    .p2998 ( optlc_net_3018 ) , .p2999 ( optlc_net_3019 ) , 
    .p3000 ( optlc_net_3020 ) , .p3001 ( optlc_net_3021 ) , 
    .p3002 ( optlc_net_3022 ) , .p3003 ( optlc_net_3023 ) , 
    .p3004 ( optlc_net_3024 ) , .p3005 ( optlc_net_3025 ) , 
    .p3006 ( optlc_net_3026 ) , .p3007 ( optlc_net_3027 ) , 
    .p3008 ( optlc_net_3028 ) , .p3009 ( optlc_net_3029 ) , 
    .p3010 ( optlc_net_3030 ) , .p3011 ( optlc_net_3031 ) , 
    .p3012 ( optlc_net_3032 ) , .p3013 ( optlc_net_3033 ) , 
    .p3014 ( optlc_net_3034 ) , .p3015 ( optlc_net_3035 ) , 
    .p3016 ( optlc_net_3036 ) , .p3017 ( optlc_net_3037 ) , 
    .p3018 ( optlc_net_3038 ) , .p3019 ( optlc_net_3039 ) , 
    .p3020 ( optlc_net_3040 ) , .p3021 ( optlc_net_3041 ) , 
    .p3022 ( optlc_net_3042 ) , .p3023 ( optlc_net_3043 ) , 
    .p3024 ( optlc_net_3044 ) , .p3025 ( optlc_net_3045 ) , 
    .p3026 ( optlc_net_3046 ) , .p3027 ( optlc_net_3047 ) , 
    .p3028 ( optlc_net_3048 ) , .p3029 ( optlc_net_3049 ) , 
    .p3030 ( optlc_net_3050 ) , .p3031 ( optlc_net_3051 ) , 
    .p3032 ( optlc_net_3052 ) , .p3033 ( optlc_net_3053 ) , 
    .p3034 ( optlc_net_3054 ) , .p3035 ( optlc_net_3055 ) , 
    .p3036 ( optlc_net_3056 ) , .p3037 ( optlc_net_3057 ) , 
    .p3038 ( optlc_net_3058 ) , .p3039 ( optlc_net_3059 ) , 
    .p3040 ( optlc_net_3060 ) , .p3041 ( optlc_net_3061 ) , 
    .p3042 ( optlc_net_3062 ) , .p3043 ( optlc_net_3063 ) , 
    .p3044 ( optlc_net_3064 ) , .p3045 ( optlc_net_3065 ) , 
    .p3046 ( optlc_net_3066 ) , .p3047 ( optlc_net_3067 ) , 
    .p3048 ( optlc_net_3068 ) , .p3049 ( optlc_net_3069 ) , 
    .p3050 ( optlc_net_3070 ) , .p3051 ( optlc_net_3071 ) , 
    .p3052 ( optlc_net_3072 ) , .p3053 ( optlc_net_3073 ) , 
    .p3054 ( optlc_net_3074 ) , .p3055 ( optlc_net_3075 ) , 
    .p3056 ( optlc_net_3076 ) , .p3057 ( optlc_net_3077 ) , 
    .p3058 ( optlc_net_3078 ) , .p3059 ( optlc_net_3079 ) , 
    .p3060 ( optlc_net_3080 ) , .p3061 ( optlc_net_3081 ) , 
    .p3062 ( optlc_net_3082 ) , .p3063 ( optlc_net_3083 ) , 
    .p3064 ( optlc_net_3084 ) , .p3065 ( optlc_net_3085 ) , 
    .p3066 ( optlc_net_3086 ) , .p3067 ( optlc_net_3087 ) , 
    .p3068 ( optlc_net_3088 ) , .p3069 ( optlc_net_3089 ) , 
    .p3070 ( optlc_net_3090 ) , .p3071 ( optlc_net_3091 ) , 
    .p3072 ( optlc_net_3092 ) , .p3073 ( optlc_net_3093 ) , 
    .p3074 ( optlc_net_3094 ) , .p3075 ( optlc_net_3095 ) , 
    .p3076 ( optlc_net_3096 ) , .p3077 ( optlc_net_3097 ) , 
    .p3078 ( optlc_net_3098 ) , .p3079 ( optlc_net_3099 ) , 
    .p3080 ( optlc_net_3100 ) , .p3081 ( optlc_net_3101 ) , 
    .p3082 ( optlc_net_3102 ) , .p3083 ( optlc_net_3103 ) , 
    .p3084 ( optlc_net_3104 ) , .p3085 ( optlc_net_3105 ) , 
    .p3086 ( optlc_net_3106 ) , .p3087 ( optlc_net_3107 ) , 
    .p3088 ( optlc_net_3108 ) , .p3089 ( optlc_net_3109 ) , 
    .p3090 ( optlc_net_3110 ) , .p3091 ( optlc_net_3111 ) , 
    .p3092 ( optlc_net_3112 ) , .p3093 ( optlc_net_3113 ) , 
    .p3094 ( optlc_net_3114 ) , .p3095 ( optlc_net_3115 ) , 
    .p3096 ( optlc_net_3116 ) , .p3097 ( optlc_net_3117 ) , 
    .p3098 ( optlc_net_3118 ) , .p3099 ( optlc_net_3119 ) , 
    .p3100 ( optlc_net_3120 ) , .p3101 ( optlc_net_3121 ) , 
    .p3102 ( optlc_net_3122 ) , .p3103 ( optlc_net_3123 ) , 
    .p3104 ( optlc_net_3124 ) , .p3105 ( optlc_net_3125 ) , 
    .p3106 ( optlc_net_3126 ) , .p3107 ( optlc_net_3127 ) , 
    .p3108 ( optlc_net_3128 ) , .p3109 ( optlc_net_3129 ) , 
    .p3110 ( optlc_net_3130 ) , .p3111 ( optlc_net_3131 ) , 
    .p3112 ( optlc_net_3132 ) , .p3113 ( optlc_net_3133 ) , 
    .p3114 ( optlc_net_3134 ) , .p3115 ( optlc_net_3135 ) , 
    .p3116 ( optlc_net_3136 ) , .p3117 ( optlc_net_3137 ) , 
    .p3118 ( optlc_net_3138 ) , .p3119 ( optlc_net_3139 ) , 
    .p3120 ( optlc_net_3140 ) , .p3121 ( optlc_net_3141 ) , 
    .p3122 ( optlc_net_3142 ) , .p3123 ( optlc_net_3143 ) , 
    .p3124 ( optlc_net_3144 ) , .p3125 ( optlc_net_3145 ) , 
    .p3126 ( optlc_net_3146 ) , .p3127 ( optlc_net_3147 ) , 
    .p3128 ( optlc_net_3148 ) , .p3129 ( optlc_net_3149 ) , 
    .p3130 ( optlc_net_3150 ) , .p3131 ( optlc_net_3151 ) , 
    .p3132 ( optlc_net_3152 ) , .p3133 ( optlc_net_3153 ) , 
    .p3134 ( optlc_net_3154 ) , .p3135 ( optlc_net_3155 ) , 
    .p3136 ( optlc_net_3156 ) , .p3137 ( optlc_net_3157 ) , 
    .p3138 ( optlc_net_3158 ) , .p3139 ( optlc_net_3159 ) , 
    .p3140 ( optlc_net_3160 ) , .p3141 ( optlc_net_3161 ) , 
    .p3142 ( optlc_net_3162 ) , .p3143 ( optlc_net_3163 ) , 
    .p3144 ( optlc_net_3164 ) , .p3145 ( optlc_net_3165 ) , 
    .p3146 ( optlc_net_3166 ) , .p3147 ( optlc_net_3167 ) , 
    .p3148 ( optlc_net_3168 ) , .p3149 ( optlc_net_3169 ) , 
    .p3150 ( optlc_net_3170 ) , .p3151 ( optlc_net_3171 ) , 
    .p3152 ( optlc_net_3172 ) , .p3153 ( optlc_net_3173 ) , 
    .p3154 ( optlc_net_3174 ) , .p3155 ( optlc_net_3175 ) , 
    .p3156 ( optlc_net_3176 ) , .p3157 ( optlc_net_3177 ) , 
    .p3158 ( optlc_net_3178 ) , .p3159 ( optlc_net_3179 ) , 
    .p3160 ( optlc_net_3180 ) , .p3161 ( optlc_net_3181 ) , 
    .p3162 ( optlc_net_3182 ) , .p3163 ( optlc_net_3183 ) , 
    .p3164 ( optlc_net_3184 ) , .p3165 ( optlc_net_3185 ) , 
    .p3166 ( optlc_net_3186 ) , .p3167 ( optlc_net_3187 ) , 
    .p3168 ( optlc_net_3188 ) , .p3169 ( optlc_net_3189 ) , 
    .p3170 ( optlc_net_3190 ) , .p3171 ( optlc_net_3191 ) , 
    .p3172 ( optlc_net_3192 ) , .p3173 ( optlc_net_3193 ) , 
    .p3174 ( optlc_net_3194 ) , .p3175 ( optlc_net_3195 ) , 
    .p3176 ( optlc_net_3196 ) , .p3177 ( optlc_net_3197 ) , 
    .p3178 ( optlc_net_3198 ) , .p3179 ( optlc_net_3199 ) , 
    .p3180 ( optlc_net_3200 ) , .p3181 ( optlc_net_3201 ) , 
    .p3182 ( optlc_net_3202 ) , .p3183 ( optlc_net_3203 ) , 
    .p3184 ( optlc_net_3204 ) , .p3185 ( optlc_net_3205 ) , 
    .p3186 ( optlc_net_3206 ) , .p3187 ( optlc_net_3207 ) , 
    .p3188 ( optlc_net_3208 ) , .p3189 ( optlc_net_3209 ) , 
    .p3190 ( optlc_net_3210 ) , .p3191 ( optlc_net_3211 ) , 
    .p3192 ( optlc_net_3212 ) , .p3193 ( optlc_net_3213 ) , 
    .p3194 ( optlc_net_3214 ) , .p3195 ( optlc_net_3215 ) , 
    .p3196 ( optlc_net_3216 ) , .p3197 ( optlc_net_3217 ) , 
    .p3198 ( optlc_net_3218 ) , .p3199 ( optlc_net_3219 ) , 
    .p3200 ( optlc_net_3220 ) , .p3201 ( optlc_net_3221 ) , 
    .p3202 ( optlc_net_3222 ) , .p3203 ( optlc_net_3223 ) , 
    .p3204 ( optlc_net_3224 ) , .p3205 ( optlc_net_3225 ) , 
    .p3206 ( optlc_net_3226 ) , .p3207 ( optlc_net_3227 ) , 
    .p3208 ( optlc_net_3228 ) , .p3209 ( optlc_net_3229 ) , 
    .p3210 ( optlc_net_3230 ) , .p3211 ( optlc_net_3231 ) , 
    .p3212 ( optlc_net_3232 ) , .p3213 ( optlc_net_3233 ) , 
    .p3214 ( optlc_net_3234 ) , .p3215 ( optlc_net_3235 ) , 
    .p3216 ( optlc_net_3236 ) , .p3217 ( optlc_net_3237 ) , 
    .p3218 ( optlc_net_3238 ) , .p3219 ( optlc_net_3239 ) , 
    .p3220 ( optlc_net_3240 ) , .p3221 ( optlc_net_3241 ) , 
    .p3222 ( optlc_net_3242 ) , .p3223 ( optlc_net_3243 ) , 
    .p3224 ( optlc_net_3244 ) , .p3225 ( optlc_net_3245 ) , 
    .p3226 ( optlc_net_3246 ) , .p3227 ( optlc_net_3247 ) , 
    .p3228 ( optlc_net_3248 ) , .p3229 ( optlc_net_3249 ) , 
    .p3230 ( optlc_net_3250 ) , .p3231 ( optlc_net_3251 ) , 
    .p3232 ( optlc_net_3252 ) , .p3233 ( optlc_net_3253 ) , 
    .p3234 ( optlc_net_3254 ) , .p3235 ( optlc_net_3255 ) , 
    .p3236 ( optlc_net_3256 ) , .p3237 ( optlc_net_3257 ) , 
    .p3238 ( optlc_net_3258 ) , .p3239 ( optlc_net_3259 ) , 
    .p3240 ( optlc_net_3260 ) , .p3241 ( optlc_net_3261 ) , 
    .p3242 ( optlc_net_3262 ) , .p3243 ( optlc_net_3263 ) , 
    .p3244 ( optlc_net_3264 ) , .p3245 ( optlc_net_3265 ) , 
    .p3246 ( optlc_net_3266 ) , .p3247 ( optlc_net_3267 ) , 
    .p3248 ( optlc_net_3268 ) , .p3249 ( optlc_net_3269 ) , 
    .p3250 ( optlc_net_3270 ) , .p3251 ( optlc_net_3271 ) , 
    .p3252 ( optlc_net_3272 ) , .p3253 ( optlc_net_3273 ) , 
    .p3254 ( optlc_net_3274 ) , .p3255 ( optlc_net_3275 ) , 
    .p3256 ( optlc_net_3276 ) , .p3257 ( optlc_net_3277 ) , 
    .p3258 ( optlc_net_3278 ) , .p3259 ( optlc_net_3279 ) , 
    .p3260 ( optlc_net_3280 ) , .p3261 ( optlc_net_3281 ) , 
    .p3262 ( optlc_net_3282 ) , .p3263 ( optlc_net_3283 ) , 
    .p3264 ( optlc_net_3284 ) , .p3265 ( optlc_net_3285 ) , 
    .p3266 ( optlc_net_3286 ) , .p3267 ( optlc_net_3287 ) , 
    .p3268 ( optlc_net_3288 ) , .p3269 ( optlc_net_3289 ) , 
    .p3270 ( optlc_net_3290 ) , .p3271 ( optlc_net_3291 ) , 
    .p3272 ( optlc_net_3292 ) , .p3273 ( optlc_net_3293 ) , 
    .p3274 ( optlc_net_3294 ) , .p3275 ( optlc_net_3295 ) , 
    .p3276 ( optlc_net_3296 ) , .p3277 ( optlc_net_3297 ) , 
    .p3278 ( optlc_net_3298 ) , .p3279 ( optlc_net_3299 ) , 
    .p3280 ( optlc_net_3300 ) , .p3281 ( optlc_net_3301 ) , 
    .p3282 ( optlc_net_3302 ) , .p3283 ( optlc_net_3303 ) , 
    .p3284 ( optlc_net_3304 ) , .p3285 ( optlc_net_3305 ) , 
    .p3286 ( optlc_net_3306 ) , .p3287 ( optlc_net_3307 ) , 
    .p3288 ( optlc_net_3308 ) , .p3289 ( optlc_net_3309 ) , 
    .p3290 ( optlc_net_3310 ) , .p3291 ( optlc_net_3311 ) , 
    .p3292 ( optlc_net_3312 ) , .p3293 ( optlc_net_3313 ) , 
    .p3294 ( optlc_net_3314 ) , .p3295 ( optlc_net_3315 ) , 
    .p3296 ( optlc_net_3316 ) , .p3297 ( optlc_net_3317 ) , 
    .p3298 ( optlc_net_3318 ) , .p3299 ( optlc_net_3319 ) , 
    .p3300 ( optlc_net_3320 ) , .p3301 ( optlc_net_3321 ) , 
    .p3302 ( optlc_net_3322 ) , .p3303 ( optlc_net_3323 ) , 
    .p3304 ( optlc_net_3324 ) , .p3305 ( optlc_net_3325 ) , 
    .p3306 ( optlc_net_3326 ) , .p3307 ( optlc_net_3327 ) , 
    .p3308 ( optlc_net_3328 ) , .p3309 ( optlc_net_3329 ) , 
    .p3310 ( optlc_net_3330 ) , .p3311 ( optlc_net_3331 ) , 
    .p3312 ( optlc_net_3332 ) , .p3313 ( optlc_net_3333 ) , 
    .p3314 ( optlc_net_3334 ) , .p3315 ( optlc_net_3335 ) , 
    .p3316 ( optlc_net_3336 ) , .p3317 ( optlc_net_3337 ) , 
    .p3318 ( optlc_net_3338 ) , .p3319 ( optlc_net_3339 ) , 
    .p3320 ( optlc_net_3340 ) , .p3321 ( optlc_net_3341 ) , 
    .p3322 ( optlc_net_3342 ) , .p3323 ( optlc_net_3343 ) , 
    .p3324 ( optlc_net_3344 ) , .p3325 ( optlc_net_3345 ) , 
    .p3326 ( optlc_net_3346 ) , .p3327 ( optlc_net_3347 ) , 
    .p3328 ( optlc_net_3348 ) , .p3329 ( optlc_net_3349 ) , 
    .p3330 ( optlc_net_3350 ) , .p3331 ( optlc_net_3351 ) , 
    .p3332 ( optlc_net_3352 ) , .p3333 ( optlc_net_3353 ) , 
    .p3334 ( optlc_net_3354 ) , .p3335 ( optlc_net_3355 ) , 
    .p3336 ( optlc_net_3356 ) , .p3337 ( optlc_net_3357 ) , 
    .p3338 ( optlc_net_3358 ) , .p3339 ( optlc_net_3359 ) , 
    .p3340 ( optlc_net_3360 ) , .p3341 ( optlc_net_3361 ) , 
    .p3342 ( optlc_net_3362 ) , .p3343 ( optlc_net_3363 ) , 
    .p3344 ( optlc_net_3364 ) , .p3345 ( optlc_net_3365 ) , 
    .p3346 ( optlc_net_3366 ) , .p3347 ( optlc_net_3367 ) , 
    .p3348 ( optlc_net_3368 ) , .p3349 ( optlc_net_3369 ) , 
    .p3350 ( optlc_net_3370 ) , .p3351 ( optlc_net_3371 ) , 
    .p3352 ( optlc_net_3372 ) , .p3353 ( optlc_net_3373 ) , 
    .p3354 ( optlc_net_3374 ) , .p3355 ( optlc_net_3375 ) , 
    .p3356 ( optlc_net_3376 ) , .p3357 ( optlc_net_3377 ) , 
    .p3358 ( optlc_net_3378 ) , .p3359 ( optlc_net_3379 ) , 
    .p3360 ( optlc_net_3380 ) , .p3361 ( optlc_net_3381 ) , 
    .p3362 ( optlc_net_3382 ) , .p3363 ( optlc_net_3383 ) , 
    .p3364 ( optlc_net_3384 ) , .p3365 ( optlc_net_3385 ) , 
    .p3366 ( optlc_net_3386 ) , .p3367 ( optlc_net_3387 ) , 
    .p3368 ( optlc_net_3388 ) , .p3369 ( optlc_net_3389 ) , 
    .p3370 ( optlc_net_3390 ) , .p3371 ( optlc_net_3391 ) , 
    .p3372 ( optlc_net_3392 ) , .p3373 ( optlc_net_3393 ) , 
    .p3374 ( optlc_net_3394 ) , .p3375 ( optlc_net_3395 ) , 
    .p3376 ( optlc_net_3396 ) , .p3377 ( optlc_net_3397 ) , 
    .p3378 ( optlc_net_3398 ) , .p3379 ( optlc_net_3399 ) , 
    .p3380 ( optlc_net_3400 ) , .p3381 ( optlc_net_3401 ) , 
    .p3382 ( optlc_net_3402 ) , .p3383 ( optlc_net_3403 ) , 
    .p3384 ( optlc_net_3404 ) , .p3385 ( optlc_net_3405 ) , 
    .p3386 ( optlc_net_3406 ) , .p3387 ( optlc_net_3407 ) , 
    .p3388 ( optlc_net_3408 ) , .p3389 ( optlc_net_3409 ) , 
    .p3390 ( optlc_net_3410 ) , .p3391 ( optlc_net_3411 ) , 
    .p3392 ( optlc_net_3412 ) , .p3393 ( optlc_net_3413 ) , 
    .p3394 ( optlc_net_3414 ) , .p3395 ( optlc_net_3415 ) , 
    .p3396 ( optlc_net_3416 ) , .p3397 ( optlc_net_3417 ) , 
    .p3398 ( optlc_net_3418 ) , .p3399 ( optlc_net_3419 ) , 
    .p3400 ( optlc_net_3420 ) , .p3401 ( optlc_net_3421 ) , 
    .p3402 ( optlc_net_3422 ) , .p3403 ( optlc_net_3423 ) , 
    .p3404 ( optlc_net_3424 ) , .p3405 ( optlc_net_3425 ) , 
    .p3406 ( optlc_net_3426 ) , .p3407 ( optlc_net_3427 ) , 
    .p3408 ( optlc_net_3428 ) , .p3409 ( optlc_net_3429 ) , 
    .p3410 ( optlc_net_3430 ) , .p3411 ( optlc_net_3431 ) , 
    .p3412 ( optlc_net_3432 ) , .p3413 ( optlc_net_3433 ) , 
    .p3414 ( optlc_net_3434 ) , .p3415 ( optlc_net_3435 ) , 
    .p3416 ( optlc_net_3436 ) , .p3417 ( optlc_net_3437 ) , 
    .p3418 ( optlc_net_3438 ) , .p3419 ( optlc_net_3439 ) , 
    .p3420 ( optlc_net_3440 ) , .p3421 ( optlc_net_3441 ) , 
    .p3422 ( optlc_net_3442 ) , .p3423 ( optlc_net_3443 ) , 
    .p3424 ( optlc_net_3444 ) , .p3425 ( optlc_net_3445 ) , 
    .p3426 ( optlc_net_3446 ) , .p3427 ( optlc_net_3447 ) , 
    .p3428 ( optlc_net_3448 ) , .p3429 ( optlc_net_3449 ) , 
    .p3430 ( optlc_net_3450 ) , .p3431 ( optlc_net_3451 ) , 
    .p3432 ( optlc_net_3452 ) , .p3433 ( optlc_net_3453 ) , 
    .p3434 ( optlc_net_3454 ) , .p3435 ( optlc_net_3455 ) , 
    .p3436 ( optlc_net_3456 ) , .p3437 ( optlc_net_3457 ) , 
    .p3438 ( optlc_net_3458 ) , .p3439 ( optlc_net_3459 ) , 
    .p3440 ( optlc_net_3460 ) , .p3441 ( optlc_net_3461 ) , 
    .p3442 ( optlc_net_3462 ) , .p3443 ( optlc_net_3463 ) , 
    .p3444 ( optlc_net_3464 ) , .p3445 ( optlc_net_3465 ) , 
    .p3446 ( optlc_net_3466 ) , .p3447 ( optlc_net_3467 ) , 
    .p3448 ( optlc_net_3468 ) , .p3449 ( optlc_net_3469 ) , 
    .p3450 ( optlc_net_3470 ) , .p3451 ( optlc_net_3471 ) , 
    .p3452 ( optlc_net_3472 ) , .p3453 ( optlc_net_3473 ) , 
    .p3454 ( optlc_net_3474 ) , .p3455 ( optlc_net_3475 ) , 
    .p3456 ( optlc_net_3476 ) , .p3457 ( optlc_net_3477 ) , 
    .p3458 ( optlc_net_3478 ) , .p3459 ( optlc_net_3479 ) , 
    .p3460 ( optlc_net_3480 ) , .p3461 ( optlc_net_3481 ) , 
    .p3462 ( optlc_net_3482 ) , .p3463 ( optlc_net_3483 ) , 
    .p3464 ( optlc_net_3484 ) , .p3465 ( optlc_net_3485 ) , 
    .p3466 ( optlc_net_3486 ) , .p3467 ( optlc_net_3487 ) , 
    .p3468 ( optlc_net_3488 ) , .p3469 ( optlc_net_3489 ) , 
    .p3470 ( optlc_net_3490 ) , .p3471 ( optlc_net_3491 ) , 
    .p3472 ( optlc_net_3492 ) , .p3473 ( optlc_net_3493 ) , 
    .p3474 ( optlc_net_3494 ) , .p3475 ( optlc_net_3495 ) , 
    .p3476 ( optlc_net_3496 ) , .p3477 ( optlc_net_3497 ) , 
    .p3478 ( optlc_net_3498 ) , .p3479 ( optlc_net_3499 ) , 
    .p3480 ( optlc_net_3500 ) , .p3481 ( optlc_net_3501 ) , 
    .p3482 ( optlc_net_3502 ) , .p3483 ( optlc_net_3503 ) , 
    .p3484 ( optlc_net_3504 ) , .p3485 ( optlc_net_3505 ) , 
    .p3486 ( optlc_net_3506 ) , .p3487 ( optlc_net_3507 ) , 
    .p3488 ( optlc_net_3508 ) , .p3489 ( optlc_net_3509 ) , 
    .p3490 ( optlc_net_3510 ) , .p3491 ( optlc_net_3511 ) , 
    .p3492 ( optlc_net_3512 ) , .p3493 ( optlc_net_3513 ) , 
    .p3494 ( optlc_net_3514 ) , .p3495 ( optlc_net_3515 ) , 
    .p3496 ( optlc_net_3516 ) , .p3497 ( optlc_net_3517 ) , 
    .p3498 ( optlc_net_3518 ) , .p3499 ( optlc_net_3519 ) , 
    .p3500 ( optlc_net_3520 ) , .p3501 ( optlc_net_3521 ) , 
    .p3502 ( optlc_net_3522 ) , .p3503 ( optlc_net_3523 ) , 
    .p3504 ( optlc_net_3524 ) , .p3505 ( optlc_net_3525 ) , 
    .p3506 ( optlc_net_3526 ) , .p3507 ( optlc_net_3527 ) , 
    .p3508 ( optlc_net_3528 ) , .p3509 ( optlc_net_3529 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_0 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( io_oeb[0] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( io_oeb[1] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( io_oeb[2] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3 ( .LO ( SYNOPSYS_UNCONNECTED_5 ) , 
    .HI ( io_oeb[3] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_4 ( .LO ( SYNOPSYS_UNCONNECTED_6 ) , 
    .HI ( io_oeb[12] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_5 ( .LO ( SYNOPSYS_UNCONNECTED_7 ) , 
    .HI ( io_oeb[25] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_6 ( .LO ( SYNOPSYS_UNCONNECTED_8 ) , 
    .HI ( io_oeb[26] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_7 ( .LO ( SYNOPSYS_UNCONNECTED_9 ) , 
    .HI ( io_oeb[36] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_8 ( .LO ( SYNOPSYS_UNCONNECTED_10 ) , 
    .HI ( io_oeb[37] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_9 ( .LO ( io_oeb[11] ) , 
    .HI ( SYNOPSYS_UNCONNECTED_11 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_10 ( .LO ( io_oeb[35] ) , 
    .HI ( SYNOPSYS_UNCONNECTED_12 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_11 ( .LO ( io_out[0] ) , 
    .HI ( SYNOPSYS_UNCONNECTED_13 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_12 ( .LO ( io_out[1] ) , 
    .HI ( SYNOPSYS_UNCONNECTED_14 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_13 ( .LO ( io_out[2] ) , 
    .HI ( SYNOPSYS_UNCONNECTED_15 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_14 ( .LO ( io_out[3] ) , 
    .HI ( SYNOPSYS_UNCONNECTED_16 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_15 ( .LO ( io_out[12] ) , 
    .HI ( SYNOPSYS_UNCONNECTED_17 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_16 ( .LO ( io_out[25] ) , 
    .HI ( SYNOPSYS_UNCONNECTED_18 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_17 ( .LO ( io_out[26] ) , 
    .HI ( SYNOPSYS_UNCONNECTED_19 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_18 ( .LO ( io_out[36] ) , 
    .HI ( SYNOPSYS_UNCONNECTED_20 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_19 ( .LO ( io_out[37] ) , 
    .HI ( SYNOPSYS_UNCONNECTED_21 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_21 ( .LO ( optlc_net_20 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_22 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_23 ( .LO ( optlc_net_21 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_23 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_24 ( .LO ( optlc_net_22 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_24 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_25 ( .LO ( optlc_net_23 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_25 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_26 ( .LO ( optlc_net_24 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_26 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_27 ( .LO ( optlc_net_25 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_27 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_28 ( .LO ( optlc_net_26 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_28 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_29 ( .LO ( optlc_net_27 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_29 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_30 ( .LO ( optlc_net_28 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_30 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_31 ( .LO ( optlc_net_29 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_31 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_32 ( .LO ( optlc_net_30 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_32 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_33 ( .LO ( optlc_net_31 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_33 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_34 ( .LO ( optlc_net_32 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_34 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_35 ( .LO ( optlc_net_33 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_35 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_36 ( .LO ( optlc_net_34 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_36 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_37 ( .LO ( optlc_net_35 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_37 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_38 ( .LO ( optlc_net_36 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_38 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_39 ( .LO ( optlc_net_37 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_39 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_40 ( .LO ( optlc_net_38 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_40 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_41 ( .LO ( optlc_net_39 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_41 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_42 ( .LO ( optlc_net_40 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_42 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_43 ( .LO ( optlc_net_41 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_43 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_44 ( .LO ( optlc_net_42 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_44 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_45 ( .LO ( optlc_net_43 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_45 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_46 ( .LO ( optlc_net_44 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_46 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_47 ( .LO ( optlc_net_45 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_47 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_48 ( .LO ( optlc_net_46 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_48 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_49 ( .LO ( optlc_net_47 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_49 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_50 ( .LO ( optlc_net_48 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_50 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_51 ( .LO ( optlc_net_49 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_51 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_52 ( .LO ( optlc_net_50 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_52 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_53 ( .LO ( optlc_net_51 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_53 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_54 ( .LO ( optlc_net_52 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_54 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_55 ( .LO ( optlc_net_53 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_55 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_56 ( .LO ( optlc_net_54 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_56 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_57 ( .LO ( optlc_net_55 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_57 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_58 ( .LO ( optlc_net_56 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_58 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_59 ( .LO ( optlc_net_57 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_59 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_60 ( .LO ( optlc_net_58 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_60 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_61 ( .LO ( optlc_net_59 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_61 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_62 ( .LO ( optlc_net_60 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_62 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_63 ( .LO ( optlc_net_61 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_63 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_64 ( .LO ( optlc_net_62 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_64 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_65 ( .LO ( optlc_net_63 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_65 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_66 ( .LO ( optlc_net_64 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_66 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_67 ( .LO ( optlc_net_65 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_67 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_68 ( .LO ( optlc_net_66 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_68 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_69 ( .LO ( optlc_net_67 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_69 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_70 ( .LO ( optlc_net_68 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_70 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_71 ( .LO ( optlc_net_69 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_71 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_72 ( .LO ( optlc_net_70 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_72 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_73 ( .LO ( optlc_net_71 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_73 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_74 ( .LO ( optlc_net_72 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_74 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_75 ( .LO ( optlc_net_73 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_75 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_76 ( .LO ( optlc_net_74 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_76 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_77 ( .LO ( optlc_net_75 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_77 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_78 ( .LO ( optlc_net_76 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_78 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_79 ( .LO ( optlc_net_77 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_79 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_80 ( .LO ( optlc_net_78 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_80 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_81 ( .LO ( optlc_net_79 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_81 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_82 ( .LO ( optlc_net_80 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_82 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_83 ( .LO ( optlc_net_81 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_83 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_84 ( .LO ( optlc_net_82 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_84 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_85 ( .LO ( optlc_net_83 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_85 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_86 ( .LO ( optlc_net_84 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_86 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_87 ( .LO ( optlc_net_85 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_87 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_88 ( .LO ( optlc_net_86 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_88 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_89 ( .LO ( optlc_net_87 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_89 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_90 ( .LO ( optlc_net_88 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_90 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_91 ( .LO ( optlc_net_89 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_91 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_92 ( .LO ( optlc_net_90 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_92 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_93 ( .LO ( optlc_net_91 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_93 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_94 ( .LO ( optlc_net_92 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_94 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_95 ( .LO ( optlc_net_93 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_95 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_96 ( .LO ( optlc_net_94 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_96 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_97 ( .LO ( optlc_net_95 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_97 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_98 ( .LO ( optlc_net_96 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_98 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_99 ( .LO ( optlc_net_97 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_99 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_100 ( .LO ( optlc_net_98 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_100 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_101 ( .LO ( optlc_net_99 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_101 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_102 ( .LO ( optlc_net_100 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_102 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_103 ( .LO ( optlc_net_101 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_103 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_104 ( .LO ( optlc_net_102 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_104 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_105 ( .LO ( optlc_net_103 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_105 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_106 ( .LO ( optlc_net_104 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_106 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_107 ( .LO ( optlc_net_105 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_107 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_108 ( .LO ( optlc_net_106 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_108 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_109 ( .LO ( optlc_net_107 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_109 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_110 ( .LO ( optlc_net_108 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_110 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_111 ( .LO ( optlc_net_109 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_111 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_112 ( .LO ( optlc_net_110 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_112 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_113 ( .LO ( optlc_net_111 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_113 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_114 ( .LO ( optlc_net_112 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_114 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_115 ( .LO ( optlc_net_113 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_115 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_116 ( .LO ( optlc_net_114 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_116 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_117 ( .LO ( optlc_net_115 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_117 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_118 ( .LO ( optlc_net_116 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_118 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_119 ( .LO ( optlc_net_117 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_119 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_120 ( .LO ( optlc_net_118 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_120 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_121 ( .LO ( optlc_net_119 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_121 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_122 ( .LO ( optlc_net_120 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_122 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_123 ( .LO ( optlc_net_121 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_123 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_124 ( .LO ( optlc_net_122 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_124 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_125 ( .LO ( optlc_net_123 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_125 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_126 ( .LO ( optlc_net_124 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_126 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_127 ( .LO ( optlc_net_125 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_127 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_128 ( .LO ( optlc_net_126 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_128 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_129 ( .LO ( optlc_net_127 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_129 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_130 ( .LO ( optlc_net_128 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_130 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_131 ( .LO ( optlc_net_129 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_131 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_132 ( .LO ( optlc_net_130 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_132 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_133 ( .LO ( optlc_net_131 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_133 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_134 ( .LO ( optlc_net_132 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_134 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_135 ( .LO ( optlc_net_133 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_135 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_136 ( .LO ( optlc_net_134 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_136 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_137 ( .LO ( optlc_net_135 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_137 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_138 ( .LO ( optlc_net_136 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_138 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_139 ( .LO ( optlc_net_137 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_139 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_140 ( .LO ( optlc_net_138 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_140 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_141 ( .LO ( optlc_net_139 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_141 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_142 ( .LO ( optlc_net_140 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_142 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_143 ( .LO ( optlc_net_141 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_143 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_144 ( .LO ( optlc_net_142 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_144 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_145 ( .LO ( optlc_net_143 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_145 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_146 ( .LO ( optlc_net_144 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_146 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_147 ( .LO ( optlc_net_145 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_147 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_148 ( .LO ( optlc_net_146 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_148 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_149 ( .LO ( optlc_net_147 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_149 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_150 ( .LO ( optlc_net_148 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_150 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_151 ( .LO ( optlc_net_149 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_151 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_152 ( .LO ( optlc_net_150 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_152 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_153 ( .LO ( optlc_net_151 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_153 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_154 ( .LO ( optlc_net_152 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_154 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_155 ( .LO ( optlc_net_153 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_155 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_156 ( .LO ( optlc_net_154 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_156 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_157 ( .LO ( optlc_net_155 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_157 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_158 ( .LO ( optlc_net_156 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_158 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_159 ( .LO ( optlc_net_157 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_159 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_160 ( .LO ( optlc_net_158 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_160 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_161 ( .LO ( optlc_net_159 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_161 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_162 ( .LO ( optlc_net_160 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_162 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_163 ( .LO ( optlc_net_161 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_163 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_164 ( .LO ( optlc_net_162 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_164 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_165 ( .LO ( optlc_net_163 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_165 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_166 ( .LO ( optlc_net_164 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_166 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_167 ( .LO ( optlc_net_165 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_167 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_168 ( .LO ( optlc_net_166 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_168 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_169 ( .LO ( optlc_net_167 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_169 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_170 ( .LO ( optlc_net_168 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_170 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_171 ( .LO ( optlc_net_169 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_171 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_172 ( .LO ( optlc_net_170 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_172 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_173 ( .LO ( optlc_net_171 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_173 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_174 ( .LO ( optlc_net_172 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_174 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_175 ( .LO ( optlc_net_173 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_175 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_176 ( .LO ( optlc_net_174 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_176 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_177 ( .LO ( optlc_net_175 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_177 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_178 ( .LO ( optlc_net_176 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_178 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_179 ( .LO ( optlc_net_177 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_179 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_180 ( .LO ( optlc_net_178 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_180 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_181 ( .LO ( optlc_net_179 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_181 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_182 ( .LO ( optlc_net_180 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_182 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_183 ( .LO ( optlc_net_181 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_183 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_184 ( .LO ( optlc_net_182 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_184 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_185 ( .LO ( optlc_net_183 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_185 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_186 ( .LO ( optlc_net_184 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_186 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_187 ( .LO ( optlc_net_185 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_187 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_188 ( .LO ( optlc_net_186 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_188 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_189 ( .LO ( optlc_net_187 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_189 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_190 ( .LO ( optlc_net_188 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_190 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_191 ( .LO ( optlc_net_189 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_191 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_192 ( .LO ( optlc_net_190 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_192 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_193 ( .LO ( optlc_net_191 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_193 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_194 ( .LO ( optlc_net_192 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_194 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_195 ( .LO ( optlc_net_193 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_195 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_196 ( .LO ( optlc_net_194 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_196 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_197 ( .LO ( optlc_net_195 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_197 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_198 ( .LO ( optlc_net_196 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_198 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_199 ( .LO ( optlc_net_197 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_199 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_200 ( .LO ( optlc_net_198 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_200 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_201 ( .LO ( optlc_net_199 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_201 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_202 ( .LO ( optlc_net_200 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_202 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_203 ( .LO ( optlc_net_201 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_203 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_204 ( .LO ( optlc_net_202 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_204 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_205 ( .LO ( optlc_net_203 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_205 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_206 ( .LO ( optlc_net_204 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_206 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_207 ( .LO ( optlc_net_205 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_207 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_208 ( .LO ( optlc_net_206 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_208 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_209 ( .LO ( optlc_net_207 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_209 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_210 ( .LO ( optlc_net_208 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_210 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_211 ( .LO ( optlc_net_209 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_211 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_212 ( .LO ( optlc_net_210 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_212 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_213 ( .LO ( optlc_net_211 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_213 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_214 ( .LO ( optlc_net_212 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_214 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_215 ( .LO ( optlc_net_213 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_215 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_216 ( .LO ( optlc_net_214 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_216 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_217 ( .LO ( optlc_net_215 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_217 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_218 ( .LO ( optlc_net_216 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_218 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_219 ( .LO ( optlc_net_217 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_219 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_220 ( .LO ( optlc_net_218 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_220 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_221 ( .LO ( optlc_net_219 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_221 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_222 ( .LO ( optlc_net_220 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_222 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_223 ( .LO ( optlc_net_221 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_223 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_224 ( .LO ( optlc_net_222 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_224 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_225 ( .LO ( optlc_net_223 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_225 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_226 ( .LO ( optlc_net_224 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_226 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_227 ( .LO ( optlc_net_225 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_227 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_228 ( .LO ( optlc_net_226 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_228 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_229 ( .LO ( optlc_net_227 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_229 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_230 ( .LO ( optlc_net_228 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_230 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_231 ( .LO ( optlc_net_229 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_231 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_232 ( .LO ( optlc_net_230 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_232 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_233 ( .LO ( optlc_net_231 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_233 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_234 ( .LO ( optlc_net_232 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_234 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_235 ( .LO ( optlc_net_233 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_235 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_236 ( .LO ( optlc_net_234 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_236 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_237 ( .LO ( optlc_net_235 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_237 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_238 ( .LO ( optlc_net_236 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_238 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_239 ( .LO ( optlc_net_237 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_239 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_240 ( .LO ( optlc_net_238 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_240 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_241 ( .LO ( optlc_net_239 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_241 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_242 ( .LO ( optlc_net_240 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_242 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_243 ( .LO ( optlc_net_241 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_243 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_244 ( .LO ( optlc_net_242 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_244 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_245 ( .LO ( optlc_net_243 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_245 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_246 ( .LO ( optlc_net_244 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_246 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_247 ( .LO ( optlc_net_245 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_247 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_248 ( .LO ( optlc_net_246 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_248 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_249 ( .LO ( optlc_net_247 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_249 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_250 ( .LO ( optlc_net_248 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_250 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_251 ( .LO ( optlc_net_249 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_251 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_252 ( .LO ( optlc_net_250 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_252 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_253 ( .LO ( optlc_net_251 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_253 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_254 ( .LO ( optlc_net_252 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_254 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_255 ( .LO ( optlc_net_253 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_255 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_256 ( .LO ( optlc_net_254 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_256 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_257 ( .LO ( optlc_net_255 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_257 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_258 ( .LO ( optlc_net_256 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_258 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_259 ( .LO ( optlc_net_257 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_259 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_260 ( .LO ( optlc_net_258 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_260 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_261 ( .LO ( optlc_net_259 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_261 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_262 ( .LO ( optlc_net_260 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_262 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_263 ( .LO ( optlc_net_261 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_263 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_264 ( .LO ( optlc_net_262 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_264 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_265 ( .LO ( optlc_net_263 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_265 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_266 ( .LO ( optlc_net_264 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_266 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_267 ( .LO ( optlc_net_265 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_267 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_268 ( .LO ( optlc_net_266 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_268 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_269 ( .LO ( optlc_net_267 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_269 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_270 ( .LO ( optlc_net_268 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_270 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_271 ( .LO ( optlc_net_269 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_271 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_272 ( .LO ( optlc_net_270 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_272 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_273 ( .LO ( optlc_net_271 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_273 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_274 ( .LO ( optlc_net_272 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_274 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_275 ( .LO ( optlc_net_273 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_275 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_276 ( .LO ( optlc_net_274 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_276 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_277 ( .LO ( optlc_net_275 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_277 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_278 ( .LO ( optlc_net_276 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_278 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_279 ( .LO ( optlc_net_277 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_279 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_280 ( .LO ( optlc_net_278 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_280 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_281 ( .LO ( optlc_net_279 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_281 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_282 ( .LO ( optlc_net_280 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_282 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_283 ( .LO ( optlc_net_281 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_283 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_284 ( .LO ( optlc_net_282 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_284 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_285 ( .LO ( optlc_net_283 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_285 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_286 ( .LO ( optlc_net_284 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_286 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_287 ( .LO ( optlc_net_285 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_287 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_288 ( .LO ( optlc_net_286 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_288 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_289 ( .LO ( optlc_net_287 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_289 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_290 ( .LO ( optlc_net_288 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_290 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_291 ( .LO ( optlc_net_289 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_291 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_292 ( .LO ( optlc_net_290 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_292 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_293 ( .LO ( optlc_net_291 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_293 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_294 ( .LO ( optlc_net_292 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_294 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_295 ( .LO ( optlc_net_293 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_295 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_296 ( .LO ( optlc_net_294 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_296 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_297 ( .LO ( optlc_net_295 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_297 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_298 ( .LO ( optlc_net_296 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_298 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_299 ( .LO ( optlc_net_297 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_299 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_300 ( .LO ( optlc_net_298 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_300 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_301 ( .LO ( optlc_net_299 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_301 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_302 ( .LO ( optlc_net_300 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_302 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_303 ( .LO ( optlc_net_301 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_303 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_304 ( .LO ( optlc_net_302 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_304 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_305 ( .LO ( optlc_net_303 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_305 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_306 ( .LO ( optlc_net_304 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_306 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_307 ( .LO ( optlc_net_305 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_307 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_308 ( .LO ( optlc_net_306 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_308 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_309 ( .LO ( optlc_net_307 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_309 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_310 ( .LO ( optlc_net_308 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_310 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_311 ( .LO ( optlc_net_309 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_311 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_312 ( .LO ( optlc_net_310 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_312 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_313 ( .LO ( optlc_net_311 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_313 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_314 ( .LO ( optlc_net_312 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_314 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_315 ( .LO ( optlc_net_313 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_315 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_316 ( .LO ( optlc_net_314 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_316 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_317 ( .LO ( optlc_net_315 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_317 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_318 ( .LO ( optlc_net_316 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_318 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_319 ( .LO ( optlc_net_317 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_319 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_320 ( .LO ( optlc_net_318 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_320 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_321 ( .LO ( optlc_net_319 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_321 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_322 ( .LO ( optlc_net_320 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_322 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_323 ( .LO ( optlc_net_321 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_323 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_324 ( .LO ( optlc_net_322 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_324 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_325 ( .LO ( optlc_net_323 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_325 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_326 ( .LO ( optlc_net_324 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_326 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_327 ( .LO ( optlc_net_325 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_327 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_328 ( .LO ( optlc_net_326 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_328 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_329 ( .LO ( optlc_net_327 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_329 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_330 ( .LO ( optlc_net_328 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_330 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_331 ( .LO ( optlc_net_329 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_331 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_332 ( .LO ( optlc_net_330 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_332 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_333 ( .LO ( optlc_net_331 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_333 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_334 ( .LO ( optlc_net_332 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_334 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_335 ( .LO ( optlc_net_333 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_335 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_336 ( .LO ( optlc_net_334 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_336 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_337 ( .LO ( optlc_net_335 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_337 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_338 ( .LO ( optlc_net_336 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_338 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_339 ( .LO ( optlc_net_337 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_339 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_340 ( .LO ( optlc_net_338 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_340 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_341 ( .LO ( optlc_net_339 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_341 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_342 ( .LO ( optlc_net_340 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_342 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_343 ( .LO ( optlc_net_341 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_343 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_344 ( .LO ( optlc_net_342 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_344 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_345 ( .LO ( optlc_net_343 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_345 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_346 ( .LO ( optlc_net_344 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_346 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_347 ( .LO ( optlc_net_345 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_347 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_348 ( .LO ( optlc_net_346 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_348 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_349 ( .LO ( optlc_net_347 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_349 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_350 ( .LO ( optlc_net_348 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_350 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_351 ( .LO ( optlc_net_349 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_351 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_352 ( .LO ( optlc_net_350 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_352 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_353 ( .LO ( optlc_net_351 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_353 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_354 ( .LO ( optlc_net_352 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_354 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_355 ( .LO ( optlc_net_353 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_355 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_356 ( .LO ( optlc_net_354 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_356 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_357 ( .LO ( optlc_net_355 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_357 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_358 ( .LO ( optlc_net_356 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_358 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_359 ( .LO ( optlc_net_357 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_359 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_360 ( .LO ( optlc_net_358 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_360 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_361 ( .LO ( optlc_net_359 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_361 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_362 ( .LO ( optlc_net_360 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_362 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_363 ( .LO ( optlc_net_361 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_363 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_364 ( .LO ( optlc_net_362 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_364 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_365 ( .LO ( optlc_net_363 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_365 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_366 ( .LO ( optlc_net_364 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_366 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_367 ( .LO ( optlc_net_365 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_367 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_368 ( .LO ( optlc_net_366 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_368 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_369 ( .LO ( optlc_net_367 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_369 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_370 ( .LO ( optlc_net_368 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_370 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_371 ( .LO ( optlc_net_369 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_371 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_372 ( .LO ( optlc_net_370 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_372 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_373 ( .LO ( optlc_net_371 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_373 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_374 ( .LO ( optlc_net_372 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_374 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_375 ( .LO ( optlc_net_373 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_375 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_376 ( .LO ( optlc_net_374 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_376 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_377 ( .LO ( optlc_net_375 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_377 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_378 ( .LO ( optlc_net_376 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_378 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_379 ( .LO ( optlc_net_377 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_379 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_380 ( .LO ( optlc_net_378 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_380 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_381 ( .LO ( optlc_net_379 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_381 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_382 ( .LO ( optlc_net_380 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_382 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_383 ( .LO ( optlc_net_381 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_383 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_384 ( .LO ( optlc_net_382 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_384 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_385 ( .LO ( optlc_net_383 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_385 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_386 ( .LO ( optlc_net_384 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_386 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_387 ( .LO ( optlc_net_385 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_387 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_388 ( .LO ( optlc_net_386 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_388 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_389 ( .LO ( optlc_net_387 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_389 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_390 ( .LO ( optlc_net_388 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_390 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_391 ( .LO ( optlc_net_389 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_391 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_392 ( .LO ( optlc_net_390 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_392 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_393 ( .LO ( optlc_net_391 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_393 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_394 ( .LO ( optlc_net_392 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_394 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_395 ( .LO ( optlc_net_393 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_395 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_396 ( .LO ( optlc_net_394 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_396 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_397 ( .LO ( optlc_net_395 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_397 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_398 ( .LO ( optlc_net_396 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_398 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_399 ( .LO ( optlc_net_397 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_399 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_400 ( .LO ( optlc_net_398 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_400 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_401 ( .LO ( optlc_net_399 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_401 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_402 ( .LO ( optlc_net_400 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_402 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_403 ( .LO ( optlc_net_401 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_403 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_404 ( .LO ( optlc_net_402 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_404 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_405 ( .LO ( optlc_net_403 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_405 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_406 ( .LO ( optlc_net_404 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_406 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_407 ( .LO ( optlc_net_405 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_407 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_408 ( .LO ( optlc_net_406 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_408 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_409 ( .LO ( optlc_net_407 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_409 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_410 ( .LO ( optlc_net_408 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_410 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_411 ( .LO ( optlc_net_409 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_411 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_412 ( .LO ( optlc_net_410 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_412 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_413 ( .LO ( optlc_net_411 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_413 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_414 ( .LO ( optlc_net_412 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_414 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_415 ( .LO ( optlc_net_413 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_415 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_416 ( .LO ( optlc_net_414 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_416 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_417 ( .LO ( optlc_net_415 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_417 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_418 ( .LO ( optlc_net_416 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_418 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_419 ( .LO ( optlc_net_417 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_419 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_420 ( .LO ( optlc_net_418 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_420 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_421 ( .LO ( optlc_net_419 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_421 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_422 ( .LO ( optlc_net_420 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_422 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_423 ( .LO ( optlc_net_421 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_423 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_424 ( .LO ( optlc_net_422 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_424 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_425 ( .LO ( optlc_net_423 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_425 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_426 ( .LO ( optlc_net_424 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_426 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_427 ( .LO ( optlc_net_425 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_427 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_428 ( .LO ( optlc_net_426 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_428 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_429 ( .LO ( optlc_net_427 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_429 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_430 ( .LO ( optlc_net_428 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_430 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_431 ( .LO ( optlc_net_429 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_431 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_432 ( .LO ( optlc_net_430 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_432 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_433 ( .LO ( optlc_net_431 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_433 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_434 ( .LO ( optlc_net_432 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_434 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_435 ( .LO ( optlc_net_433 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_435 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_436 ( .LO ( optlc_net_434 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_436 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_437 ( .LO ( optlc_net_435 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_437 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_438 ( .LO ( optlc_net_436 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_438 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_439 ( .LO ( optlc_net_437 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_439 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_440 ( .LO ( optlc_net_438 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_440 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_441 ( .LO ( optlc_net_439 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_441 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_442 ( .LO ( optlc_net_440 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_442 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_443 ( .LO ( optlc_net_441 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_443 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_444 ( .LO ( optlc_net_442 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_444 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_445 ( .LO ( optlc_net_443 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_445 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_446 ( .LO ( optlc_net_444 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_446 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_447 ( .LO ( optlc_net_445 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_447 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_448 ( .LO ( optlc_net_446 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_448 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_449 ( .LO ( optlc_net_447 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_449 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_450 ( .LO ( optlc_net_448 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_450 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_451 ( .LO ( optlc_net_449 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_451 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_452 ( .LO ( optlc_net_450 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_452 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_453 ( .LO ( optlc_net_451 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_453 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_454 ( .LO ( optlc_net_452 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_454 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_455 ( .LO ( optlc_net_453 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_455 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_456 ( .LO ( optlc_net_454 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_456 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_457 ( .LO ( optlc_net_455 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_457 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_458 ( .LO ( optlc_net_456 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_458 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_459 ( .LO ( optlc_net_457 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_459 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_460 ( .LO ( optlc_net_458 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_460 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_461 ( .LO ( optlc_net_459 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_461 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_462 ( .LO ( optlc_net_460 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_462 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_463 ( .LO ( optlc_net_461 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_463 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_464 ( .LO ( optlc_net_462 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_464 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_465 ( .LO ( optlc_net_463 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_465 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_466 ( .LO ( optlc_net_464 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_466 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_467 ( .LO ( optlc_net_465 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_467 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_468 ( .LO ( optlc_net_466 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_468 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_469 ( .LO ( optlc_net_467 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_469 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_470 ( .LO ( optlc_net_468 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_470 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_471 ( .LO ( optlc_net_469 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_471 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_472 ( .LO ( optlc_net_470 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_472 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_473 ( .LO ( optlc_net_471 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_473 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_474 ( .LO ( optlc_net_472 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_474 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_475 ( .LO ( optlc_net_473 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_475 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_476 ( .LO ( optlc_net_474 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_476 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_477 ( .LO ( optlc_net_475 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_477 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_478 ( .LO ( optlc_net_476 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_478 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_479 ( .LO ( optlc_net_477 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_479 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_480 ( .LO ( optlc_net_478 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_480 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_481 ( .LO ( optlc_net_479 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_481 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_482 ( .LO ( optlc_net_480 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_482 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_483 ( .LO ( optlc_net_481 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_483 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_484 ( .LO ( optlc_net_482 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_484 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_485 ( .LO ( optlc_net_483 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_485 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_486 ( .LO ( optlc_net_484 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_486 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_487 ( .LO ( optlc_net_485 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_487 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_488 ( .LO ( optlc_net_486 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_488 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_489 ( .LO ( optlc_net_487 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_489 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_490 ( .LO ( optlc_net_488 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_490 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_491 ( .LO ( optlc_net_489 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_491 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_492 ( .LO ( optlc_net_490 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_492 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_493 ( .LO ( optlc_net_491 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_493 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_494 ( .LO ( optlc_net_492 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_494 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_495 ( .LO ( optlc_net_493 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_495 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_496 ( .LO ( optlc_net_494 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_496 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_497 ( .LO ( optlc_net_495 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_497 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_498 ( .LO ( optlc_net_496 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_498 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_499 ( .LO ( optlc_net_497 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_499 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_500 ( .LO ( optlc_net_498 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_500 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_501 ( .LO ( optlc_net_499 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_501 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_502 ( .LO ( optlc_net_500 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_502 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_503 ( .LO ( optlc_net_501 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_503 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_504 ( .LO ( optlc_net_502 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_504 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_505 ( .LO ( optlc_net_503 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_505 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_506 ( .LO ( optlc_net_504 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_506 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_507 ( .LO ( optlc_net_505 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_507 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_508 ( .LO ( optlc_net_506 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_508 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_509 ( .LO ( optlc_net_507 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_509 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_510 ( .LO ( optlc_net_508 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_510 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_511 ( .LO ( optlc_net_509 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_511 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_512 ( .LO ( optlc_net_510 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_512 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_513 ( .LO ( optlc_net_511 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_513 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_514 ( .LO ( optlc_net_512 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_514 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_515 ( .LO ( optlc_net_513 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_515 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_516 ( .LO ( optlc_net_514 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_516 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_517 ( .LO ( optlc_net_515 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_517 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_518 ( .LO ( optlc_net_516 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_518 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_519 ( .LO ( optlc_net_517 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_519 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_520 ( .LO ( optlc_net_518 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_520 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_521 ( .LO ( optlc_net_519 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_521 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_522 ( .LO ( optlc_net_520 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_522 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_523 ( .LO ( optlc_net_521 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_523 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_524 ( .LO ( optlc_net_522 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_524 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_525 ( .LO ( optlc_net_523 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_525 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_526 ( .LO ( optlc_net_524 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_526 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_527 ( .LO ( optlc_net_525 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_527 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_528 ( .LO ( optlc_net_526 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_528 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_529 ( .LO ( optlc_net_527 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_529 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_530 ( .LO ( optlc_net_528 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_530 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_531 ( .LO ( optlc_net_529 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_531 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_532 ( .LO ( optlc_net_530 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_532 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_533 ( .LO ( optlc_net_531 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_533 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_534 ( .LO ( optlc_net_532 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_534 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_535 ( .LO ( optlc_net_533 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_535 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_536 ( .LO ( optlc_net_534 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_536 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_537 ( .LO ( optlc_net_535 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_537 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_538 ( .LO ( optlc_net_536 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_538 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_539 ( .LO ( optlc_net_537 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_539 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_540 ( .LO ( optlc_net_538 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_540 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_541 ( .LO ( optlc_net_539 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_541 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_542 ( .LO ( optlc_net_540 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_542 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_543 ( .LO ( optlc_net_541 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_543 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_544 ( .LO ( optlc_net_542 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_544 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_545 ( .LO ( optlc_net_543 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_545 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_546 ( .LO ( optlc_net_544 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_546 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_547 ( .LO ( optlc_net_545 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_547 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_548 ( .LO ( optlc_net_546 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_548 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_549 ( .LO ( optlc_net_547 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_549 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_550 ( .LO ( optlc_net_548 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_550 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_551 ( .LO ( optlc_net_549 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_551 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_552 ( .LO ( optlc_net_550 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_552 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_553 ( .LO ( optlc_net_551 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_553 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_554 ( .LO ( optlc_net_552 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_554 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_555 ( .LO ( optlc_net_553 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_555 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_556 ( .LO ( optlc_net_554 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_556 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_557 ( .LO ( optlc_net_555 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_557 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_558 ( .LO ( optlc_net_556 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_558 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_559 ( .LO ( optlc_net_557 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_559 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_561 ( .LO ( optlc_net_558 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_560 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_562 ( .LO ( optlc_net_559 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_561 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_563 ( .LO ( optlc_net_560 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_562 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_564 ( .LO ( optlc_net_561 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_563 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_565 ( .LO ( optlc_net_562 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_564 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_566 ( .LO ( optlc_net_563 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_565 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_567 ( .LO ( optlc_net_564 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_566 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_568 ( .LO ( optlc_net_565 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_567 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_569 ( .LO ( optlc_net_566 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_568 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_570 ( .LO ( optlc_net_567 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_569 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_571 ( .LO ( optlc_net_568 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_570 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_572 ( .LO ( optlc_net_569 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_571 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_573 ( .LO ( optlc_net_570 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_572 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_574 ( .LO ( optlc_net_571 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_573 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_575 ( .LO ( optlc_net_572 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_574 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_576 ( .LO ( optlc_net_573 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_575 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_577 ( .LO ( optlc_net_574 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_576 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_578 ( .LO ( optlc_net_575 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_577 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_579 ( .LO ( optlc_net_576 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_578 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_580 ( .LO ( optlc_net_577 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_579 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_581 ( .LO ( optlc_net_578 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_580 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_582 ( .LO ( optlc_net_579 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_581 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_583 ( .LO ( optlc_net_580 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_582 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_584 ( .LO ( optlc_net_581 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_583 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_585 ( .LO ( optlc_net_582 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_584 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_586 ( .LO ( optlc_net_583 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_585 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_587 ( .LO ( optlc_net_584 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_586 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_588 ( .LO ( optlc_net_585 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_587 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_589 ( .LO ( optlc_net_586 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_588 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_590 ( .LO ( optlc_net_587 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_589 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_591 ( .LO ( optlc_net_588 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_590 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_592 ( .LO ( optlc_net_589 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_591 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_593 ( .LO ( optlc_net_590 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_592 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_594 ( .LO ( optlc_net_591 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_593 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_595 ( .LO ( optlc_net_592 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_594 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_596 ( .LO ( optlc_net_593 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_595 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_597 ( .LO ( optlc_net_594 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_596 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_598 ( .LO ( optlc_net_595 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_597 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_599 ( .LO ( optlc_net_596 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_598 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_600 ( .LO ( optlc_net_597 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_599 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_601 ( .LO ( optlc_net_598 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_600 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_602 ( .LO ( optlc_net_599 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_601 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_603 ( .LO ( optlc_net_600 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_602 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_604 ( .LO ( optlc_net_601 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_603 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_605 ( .LO ( optlc_net_602 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_604 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_606 ( .LO ( optlc_net_603 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_605 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_607 ( .LO ( optlc_net_604 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_606 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_608 ( .LO ( optlc_net_605 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_607 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_609 ( .LO ( optlc_net_606 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_608 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_610 ( .LO ( optlc_net_607 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_609 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_611 ( .LO ( optlc_net_608 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_610 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_612 ( .LO ( optlc_net_609 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_611 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_613 ( .LO ( optlc_net_610 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_612 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_614 ( .LO ( optlc_net_611 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_613 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_615 ( .LO ( optlc_net_612 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_614 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_616 ( .LO ( optlc_net_613 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_615 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_617 ( .LO ( optlc_net_614 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_616 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_618 ( .LO ( optlc_net_615 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_617 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_619 ( .LO ( optlc_net_616 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_618 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_620 ( .LO ( optlc_net_617 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_619 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_621 ( .LO ( optlc_net_618 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_620 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_622 ( .LO ( optlc_net_619 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_621 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_623 ( .LO ( optlc_net_620 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_622 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_624 ( .LO ( optlc_net_621 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_623 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_625 ( .LO ( optlc_net_622 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_624 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_626 ( .LO ( optlc_net_623 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_625 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_627 ( .LO ( optlc_net_624 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_626 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_628 ( .LO ( optlc_net_625 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_627 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_629 ( .LO ( optlc_net_626 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_628 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_630 ( .LO ( optlc_net_627 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_629 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_631 ( .LO ( optlc_net_628 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_630 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_632 ( .LO ( optlc_net_629 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_631 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_633 ( .LO ( optlc_net_630 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_632 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_634 ( .LO ( optlc_net_631 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_633 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_635 ( .LO ( optlc_net_632 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_634 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_636 ( .LO ( optlc_net_633 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_635 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_637 ( .LO ( optlc_net_634 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_636 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_638 ( .LO ( optlc_net_635 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_637 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_639 ( .LO ( optlc_net_636 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_638 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_640 ( .LO ( optlc_net_637 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_639 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_641 ( .LO ( optlc_net_638 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_640 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_642 ( .LO ( optlc_net_639 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_641 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_643 ( .LO ( optlc_net_640 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_642 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_644 ( .LO ( optlc_net_641 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_643 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_645 ( .LO ( optlc_net_642 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_644 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_646 ( .LO ( optlc_net_643 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_645 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_647 ( .LO ( optlc_net_644 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_646 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_648 ( .LO ( optlc_net_645 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_647 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_649 ( .LO ( optlc_net_646 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_648 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_650 ( .LO ( optlc_net_647 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_649 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_651 ( .LO ( optlc_net_648 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_650 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_652 ( .LO ( optlc_net_649 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_651 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_653 ( .LO ( optlc_net_650 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_652 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_654 ( .LO ( optlc_net_651 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_653 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_655 ( .LO ( optlc_net_652 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_654 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_656 ( .LO ( optlc_net_653 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_655 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_657 ( .LO ( optlc_net_654 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_656 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_658 ( .LO ( optlc_net_655 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_657 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_659 ( .LO ( optlc_net_656 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_658 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_660 ( .LO ( optlc_net_657 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_659 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_661 ( .LO ( optlc_net_658 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_660 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_662 ( .LO ( optlc_net_659 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_661 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_663 ( .LO ( optlc_net_660 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_662 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_664 ( .LO ( optlc_net_661 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_663 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_665 ( .LO ( optlc_net_662 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_664 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_666 ( .LO ( optlc_net_663 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_665 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_667 ( .LO ( optlc_net_664 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_666 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_668 ( .LO ( optlc_net_665 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_667 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_669 ( .LO ( optlc_net_666 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_668 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_670 ( .LO ( optlc_net_667 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_669 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_671 ( .LO ( optlc_net_668 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_670 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_672 ( .LO ( optlc_net_669 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_671 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_673 ( .LO ( optlc_net_670 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_672 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_674 ( .LO ( optlc_net_671 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_673 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_675 ( .LO ( optlc_net_672 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_674 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_676 ( .LO ( optlc_net_673 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_675 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_677 ( .LO ( optlc_net_674 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_676 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_678 ( .LO ( optlc_net_675 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_677 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_679 ( .LO ( optlc_net_676 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_678 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_680 ( .LO ( optlc_net_677 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_679 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_681 ( .LO ( optlc_net_678 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_680 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_682 ( .LO ( optlc_net_679 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_681 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_683 ( .LO ( optlc_net_680 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_682 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_684 ( .LO ( optlc_net_681 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_683 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_685 ( .LO ( optlc_net_682 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_684 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_686 ( .LO ( optlc_net_683 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_685 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_687 ( .LO ( optlc_net_684 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_686 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_688 ( .LO ( optlc_net_685 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_687 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_689 ( .LO ( optlc_net_686 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_688 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_690 ( .LO ( optlc_net_687 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_689 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_691 ( .LO ( optlc_net_688 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_690 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_692 ( .LO ( optlc_net_689 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_691 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_693 ( .LO ( optlc_net_690 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_692 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_694 ( .LO ( optlc_net_691 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_693 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_695 ( .LO ( optlc_net_692 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_694 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_696 ( .LO ( optlc_net_693 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_695 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_697 ( .LO ( optlc_net_694 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_696 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_698 ( .LO ( optlc_net_695 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_697 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_699 ( .LO ( optlc_net_696 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_698 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_700 ( .LO ( optlc_net_697 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_699 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_701 ( .LO ( optlc_net_698 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_700 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_702 ( .LO ( optlc_net_699 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_701 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_703 ( .LO ( optlc_net_700 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_702 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_704 ( .LO ( optlc_net_701 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_703 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_705 ( .LO ( optlc_net_702 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_704 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_706 ( .LO ( optlc_net_703 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_705 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_708 ( .LO ( optlc_net_704 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_706 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_709 ( .LO ( optlc_net_705 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_707 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_710 ( .LO ( optlc_net_706 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_708 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_711 ( .LO ( optlc_net_707 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_709 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_712 ( .LO ( optlc_net_708 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_710 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_713 ( .LO ( optlc_net_709 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_711 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_714 ( .LO ( optlc_net_710 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_712 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_715 ( .LO ( optlc_net_711 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_713 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_716 ( .LO ( optlc_net_712 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_714 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_717 ( .LO ( optlc_net_713 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_715 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_718 ( .LO ( optlc_net_714 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_716 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_719 ( .LO ( optlc_net_715 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_717 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_720 ( .LO ( optlc_net_716 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_718 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_721 ( .LO ( optlc_net_717 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_719 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_722 ( .LO ( optlc_net_718 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_720 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_723 ( .LO ( optlc_net_719 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_721 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_724 ( .LO ( optlc_net_720 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_722 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_725 ( .LO ( optlc_net_721 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_723 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_726 ( .LO ( optlc_net_722 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_724 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_727 ( .LO ( optlc_net_723 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_725 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_728 ( .LO ( optlc_net_724 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_726 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_729 ( .LO ( optlc_net_725 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_727 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_730 ( .LO ( optlc_net_726 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_728 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_731 ( .LO ( optlc_net_727 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_729 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_732 ( .LO ( optlc_net_728 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_730 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_733 ( .LO ( optlc_net_729 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_731 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_734 ( .LO ( optlc_net_730 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_732 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_735 ( .LO ( optlc_net_731 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_733 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_736 ( .LO ( optlc_net_732 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_734 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_737 ( .LO ( optlc_net_733 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_735 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_738 ( .LO ( optlc_net_734 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_736 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_739 ( .LO ( optlc_net_735 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_737 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_740 ( .LO ( optlc_net_736 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_738 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_741 ( .LO ( optlc_net_737 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_739 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_742 ( .LO ( optlc_net_738 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_740 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_743 ( .LO ( optlc_net_739 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_741 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_744 ( .LO ( optlc_net_740 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_742 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_745 ( .LO ( optlc_net_741 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_743 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_746 ( .LO ( optlc_net_742 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_744 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_747 ( .LO ( optlc_net_743 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_745 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_748 ( .LO ( optlc_net_744 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_746 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_749 ( .LO ( optlc_net_745 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_747 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_750 ( .LO ( optlc_net_746 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_748 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_751 ( .LO ( optlc_net_747 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_749 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_752 ( .LO ( optlc_net_748 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_750 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_753 ( .LO ( optlc_net_749 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_751 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_754 ( .LO ( optlc_net_750 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_752 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_755 ( .LO ( optlc_net_751 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_753 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_756 ( .LO ( optlc_net_752 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_754 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_757 ( .LO ( optlc_net_753 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_755 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_758 ( .LO ( optlc_net_754 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_756 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_759 ( .LO ( optlc_net_755 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_757 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_760 ( .LO ( optlc_net_756 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_758 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_761 ( .LO ( optlc_net_757 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_759 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_762 ( .LO ( optlc_net_758 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_760 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_763 ( .LO ( optlc_net_759 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_761 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_764 ( .LO ( optlc_net_760 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_762 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_765 ( .LO ( optlc_net_761 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_763 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_766 ( .LO ( optlc_net_762 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_764 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_767 ( .LO ( optlc_net_763 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_765 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_768 ( .LO ( optlc_net_764 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_766 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_769 ( .LO ( optlc_net_765 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_767 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_770 ( .LO ( optlc_net_766 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_768 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_771 ( .LO ( optlc_net_767 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_769 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_772 ( .LO ( optlc_net_768 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_770 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_773 ( .LO ( optlc_net_769 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_771 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_774 ( .LO ( optlc_net_770 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_772 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_775 ( .LO ( optlc_net_771 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_773 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_776 ( .LO ( optlc_net_772 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_774 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_778 ( .LO ( optlc_net_773 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_775 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_779 ( .LO ( optlc_net_774 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_776 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_780 ( .LO ( optlc_net_775 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_777 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_781 ( .LO ( optlc_net_776 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_778 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_782 ( .LO ( optlc_net_777 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_779 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_783 ( .LO ( optlc_net_778 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_780 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_784 ( .LO ( optlc_net_779 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_781 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_785 ( .LO ( optlc_net_780 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_782 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_786 ( .LO ( optlc_net_781 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_783 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_787 ( .LO ( optlc_net_782 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_784 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_788 ( .LO ( optlc_net_783 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_785 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_789 ( .LO ( optlc_net_784 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_786 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_790 ( .LO ( optlc_net_785 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_787 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_791 ( .LO ( optlc_net_786 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_788 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_792 ( .LO ( optlc_net_787 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_789 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_793 ( .LO ( optlc_net_788 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_790 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_794 ( .LO ( optlc_net_789 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_791 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_795 ( .LO ( optlc_net_790 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_792 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_796 ( .LO ( optlc_net_791 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_793 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_797 ( .LO ( optlc_net_792 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_794 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_798 ( .LO ( optlc_net_793 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_795 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_799 ( .LO ( optlc_net_794 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_796 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_800 ( .LO ( optlc_net_795 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_797 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_801 ( .LO ( optlc_net_796 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_798 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_802 ( .LO ( optlc_net_797 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_799 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_803 ( .LO ( optlc_net_798 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_800 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_804 ( .LO ( optlc_net_799 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_801 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_805 ( .LO ( optlc_net_800 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_802 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_806 ( .LO ( optlc_net_801 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_803 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_807 ( .LO ( optlc_net_802 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_804 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_808 ( .LO ( optlc_net_803 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_805 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_809 ( .LO ( optlc_net_804 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_806 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_810 ( .LO ( optlc_net_805 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_807 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_811 ( .LO ( optlc_net_806 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_808 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_812 ( .LO ( optlc_net_807 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_809 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_813 ( .LO ( optlc_net_808 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_810 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_814 ( .LO ( optlc_net_809 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_811 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_815 ( .LO ( optlc_net_810 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_812 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_816 ( .LO ( optlc_net_811 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_813 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_817 ( .LO ( optlc_net_812 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_814 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_818 ( .LO ( optlc_net_813 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_815 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_819 ( .LO ( optlc_net_814 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_816 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_820 ( .LO ( optlc_net_815 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_817 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_821 ( .LO ( optlc_net_816 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_818 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_822 ( .LO ( optlc_net_817 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_819 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_823 ( .LO ( optlc_net_818 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_820 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_824 ( .LO ( optlc_net_819 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_821 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_825 ( .LO ( optlc_net_820 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_822 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_826 ( .LO ( optlc_net_821 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_823 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_827 ( .LO ( optlc_net_822 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_824 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_828 ( .LO ( optlc_net_823 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_825 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_829 ( .LO ( optlc_net_824 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_826 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_830 ( .LO ( optlc_net_825 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_827 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_831 ( .LO ( optlc_net_826 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_828 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_832 ( .LO ( optlc_net_827 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_829 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_833 ( .LO ( optlc_net_828 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_830 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_835 ( .LO ( optlc_net_829 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_831 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_836 ( .LO ( optlc_net_830 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_832 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_837 ( .LO ( optlc_net_831 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_833 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_838 ( .LO ( optlc_net_832 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_834 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_839 ( .LO ( optlc_net_833 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_835 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_840 ( .LO ( optlc_net_834 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_836 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_841 ( .LO ( optlc_net_835 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_837 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_842 ( .LO ( optlc_net_836 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_838 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_843 ( .LO ( optlc_net_837 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_839 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_844 ( .LO ( optlc_net_838 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_840 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_845 ( .LO ( optlc_net_839 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_841 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_846 ( .LO ( optlc_net_840 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_842 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_847 ( .LO ( optlc_net_841 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_843 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_848 ( .LO ( optlc_net_842 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_844 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_849 ( .LO ( optlc_net_843 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_845 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_850 ( .LO ( optlc_net_844 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_846 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_851 ( .LO ( optlc_net_845 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_847 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_852 ( .LO ( optlc_net_846 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_848 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_853 ( .LO ( optlc_net_847 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_849 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_854 ( .LO ( optlc_net_848 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_850 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_856 ( .LO ( optlc_net_849 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_851 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_857 ( .LO ( optlc_net_850 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_852 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_858 ( .LO ( optlc_net_851 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_853 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_859 ( .LO ( optlc_net_852 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_854 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_860 ( .LO ( optlc_net_853 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_855 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_861 ( .LO ( optlc_net_854 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_856 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_862 ( .LO ( optlc_net_855 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_857 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_863 ( .LO ( optlc_net_856 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_858 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_864 ( .LO ( optlc_net_857 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_859 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_865 ( .LO ( optlc_net_858 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_860 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_866 ( .LO ( optlc_net_859 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_861 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_867 ( .LO ( optlc_net_860 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_862 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_868 ( .LO ( optlc_net_861 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_863 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_870 ( .LO ( optlc_net_862 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_864 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_871 ( .LO ( optlc_net_863 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_865 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_872 ( .LO ( optlc_net_864 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_866 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_873 ( .LO ( optlc_net_865 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_867 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_874 ( .LO ( optlc_net_866 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_868 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_875 ( .LO ( optlc_net_867 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_869 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_876 ( .LO ( optlc_net_868 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_870 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_877 ( .LO ( optlc_net_869 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_871 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_878 ( .LO ( optlc_net_870 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_872 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_879 ( .LO ( optlc_net_871 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_873 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_880 ( .LO ( optlc_net_872 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_874 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_881 ( .LO ( optlc_net_873 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_875 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_882 ( .LO ( optlc_net_874 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_876 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_883 ( .LO ( optlc_net_875 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_877 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_884 ( .LO ( optlc_net_876 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_878 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_885 ( .LO ( optlc_net_877 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_879 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_886 ( .LO ( optlc_net_878 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_880 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_887 ( .LO ( optlc_net_879 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_881 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_888 ( .LO ( optlc_net_880 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_882 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_889 ( .LO ( optlc_net_881 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_883 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_890 ( .LO ( optlc_net_882 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_884 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_891 ( .LO ( optlc_net_883 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_885 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_892 ( .LO ( optlc_net_884 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_886 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_893 ( .LO ( optlc_net_885 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_887 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_894 ( .LO ( optlc_net_886 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_888 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_895 ( .LO ( optlc_net_887 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_889 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_896 ( .LO ( optlc_net_888 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_890 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_897 ( .LO ( optlc_net_889 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_891 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_898 ( .LO ( optlc_net_890 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_892 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_899 ( .LO ( optlc_net_891 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_893 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_900 ( .LO ( optlc_net_892 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_894 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_901 ( .LO ( optlc_net_893 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_895 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_902 ( .LO ( optlc_net_894 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_896 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_903 ( .LO ( optlc_net_895 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_897 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_904 ( .LO ( optlc_net_896 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_898 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_905 ( .LO ( optlc_net_897 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_899 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_906 ( .LO ( optlc_net_898 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_900 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_907 ( .LO ( optlc_net_899 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_901 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_908 ( .LO ( optlc_net_900 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_902 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_909 ( .LO ( optlc_net_901 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_903 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_910 ( .LO ( optlc_net_902 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_904 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_911 ( .LO ( optlc_net_903 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_905 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_912 ( .LO ( optlc_net_904 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_906 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_913 ( .LO ( optlc_net_905 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_907 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_915 ( .LO ( optlc_net_906 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_908 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_916 ( .LO ( optlc_net_907 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_909 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_917 ( .LO ( optlc_net_908 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_910 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_918 ( .LO ( optlc_net_909 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_911 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_919 ( .LO ( optlc_net_910 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_912 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_920 ( .LO ( optlc_net_911 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_913 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_921 ( .LO ( optlc_net_912 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_914 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_922 ( .LO ( optlc_net_913 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_915 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_923 ( .LO ( optlc_net_914 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_916 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_924 ( .LO ( optlc_net_915 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_917 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_925 ( .LO ( optlc_net_916 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_918 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_926 ( .LO ( optlc_net_917 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_919 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_927 ( .LO ( optlc_net_918 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_920 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_928 ( .LO ( optlc_net_919 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_921 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_929 ( .LO ( optlc_net_920 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_922 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_930 ( .LO ( optlc_net_921 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_923 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_931 ( .LO ( optlc_net_922 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_924 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_932 ( .LO ( optlc_net_923 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_925 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_933 ( .LO ( optlc_net_924 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_926 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_934 ( .LO ( optlc_net_925 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_927 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_935 ( .LO ( optlc_net_926 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_928 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_936 ( .LO ( optlc_net_927 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_929 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_937 ( .LO ( optlc_net_928 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_930 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_938 ( .LO ( optlc_net_929 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_931 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_939 ( .LO ( optlc_net_930 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_932 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_940 ( .LO ( optlc_net_931 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_933 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_941 ( .LO ( optlc_net_932 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_934 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_942 ( .LO ( optlc_net_933 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_935 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_943 ( .LO ( optlc_net_934 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_936 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_944 ( .LO ( optlc_net_935 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_937 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_945 ( .LO ( optlc_net_936 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_938 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_946 ( .LO ( optlc_net_937 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_939 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_947 ( .LO ( optlc_net_938 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_940 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_948 ( .LO ( optlc_net_939 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_941 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_949 ( .LO ( optlc_net_940 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_942 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_950 ( .LO ( optlc_net_941 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_943 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_951 ( .LO ( optlc_net_942 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_944 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_952 ( .LO ( optlc_net_943 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_945 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_953 ( .LO ( optlc_net_944 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_946 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_954 ( .LO ( optlc_net_945 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_947 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_955 ( .LO ( optlc_net_946 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_948 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_956 ( .LO ( optlc_net_947 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_949 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_957 ( .LO ( optlc_net_948 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_950 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_958 ( .LO ( optlc_net_949 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_951 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_959 ( .LO ( optlc_net_950 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_952 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_960 ( .LO ( optlc_net_951 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_953 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_961 ( .LO ( optlc_net_952 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_954 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_962 ( .LO ( optlc_net_953 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_955 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_963 ( .LO ( optlc_net_954 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_956 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_964 ( .LO ( optlc_net_955 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_957 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_965 ( .LO ( optlc_net_956 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_958 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_966 ( .LO ( optlc_net_957 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_959 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_967 ( .LO ( optlc_net_958 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_960 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_968 ( .LO ( optlc_net_959 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_961 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_969 ( .LO ( optlc_net_960 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_962 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_970 ( .LO ( optlc_net_961 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_963 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_971 ( .LO ( optlc_net_962 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_964 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_972 ( .LO ( optlc_net_963 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_965 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_973 ( .LO ( optlc_net_964 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_966 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_974 ( .LO ( optlc_net_965 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_967 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_975 ( .LO ( optlc_net_966 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_968 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_976 ( .LO ( optlc_net_967 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_969 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_977 ( .LO ( optlc_net_968 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_970 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_978 ( .LO ( optlc_net_969 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_971 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_979 ( .LO ( optlc_net_970 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_972 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_980 ( .LO ( optlc_net_971 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_973 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_981 ( .LO ( optlc_net_972 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_974 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_982 ( .LO ( optlc_net_973 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_975 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_983 ( .LO ( optlc_net_974 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_976 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_984 ( .LO ( optlc_net_975 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_977 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_985 ( .LO ( optlc_net_976 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_978 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_986 ( .LO ( optlc_net_977 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_979 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_987 ( .LO ( optlc_net_978 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_980 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_988 ( .LO ( optlc_net_979 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_981 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_989 ( .LO ( optlc_net_980 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_982 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_990 ( .LO ( optlc_net_981 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_983 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_992 ( .LO ( optlc_net_982 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_984 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_993 ( .LO ( optlc_net_983 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_985 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_994 ( .LO ( optlc_net_984 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_986 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_995 ( .LO ( optlc_net_985 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_987 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_996 ( .LO ( optlc_net_986 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_988 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_997 ( .LO ( optlc_net_987 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_989 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_998 ( .LO ( optlc_net_988 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_990 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_999 ( .LO ( optlc_net_989 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_991 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1000 ( .LO ( optlc_net_990 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_992 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1001 ( .LO ( optlc_net_991 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_993 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1002 ( .LO ( optlc_net_992 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_994 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1003 ( .LO ( optlc_net_993 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_995 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1004 ( .LO ( optlc_net_994 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_996 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1005 ( .LO ( optlc_net_995 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_997 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1006 ( .LO ( optlc_net_996 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_998 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1007 ( .LO ( optlc_net_997 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_999 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1008 ( .LO ( optlc_net_998 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1000 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1009 ( .LO ( optlc_net_999 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1001 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1010 ( .LO ( optlc_net_1000 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1002 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1012 ( .LO ( optlc_net_1001 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1003 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1013 ( .LO ( optlc_net_1002 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1004 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1014 ( .LO ( optlc_net_1003 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1005 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1015 ( .LO ( optlc_net_1004 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1006 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1016 ( .LO ( optlc_net_1005 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1007 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1017 ( .LO ( optlc_net_1006 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1008 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1018 ( .LO ( optlc_net_1007 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1009 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1019 ( .LO ( optlc_net_1008 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1010 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1020 ( .LO ( optlc_net_1009 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1011 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1021 ( .LO ( optlc_net_1010 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1012 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1022 ( .LO ( optlc_net_1011 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1013 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1023 ( .LO ( optlc_net_1012 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1014 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1024 ( .LO ( optlc_net_1013 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1015 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1025 ( .LO ( optlc_net_1014 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1016 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1026 ( .LO ( optlc_net_1015 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1017 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1027 ( .LO ( optlc_net_1016 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1018 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1028 ( .LO ( optlc_net_1017 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1019 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1029 ( .LO ( optlc_net_1018 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1020 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1030 ( .LO ( optlc_net_1019 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1021 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1031 ( .LO ( optlc_net_1020 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1022 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1032 ( .LO ( optlc_net_1021 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1023 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1033 ( .LO ( optlc_net_1022 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1024 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1034 ( .LO ( optlc_net_1023 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1025 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1035 ( .LO ( optlc_net_1024 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1026 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1036 ( .LO ( optlc_net_1025 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1027 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1037 ( .LO ( optlc_net_1026 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1028 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1038 ( .LO ( optlc_net_1027 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1029 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1039 ( .LO ( optlc_net_1028 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1030 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1040 ( .LO ( optlc_net_1029 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1031 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1041 ( .LO ( optlc_net_1030 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1032 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1042 ( .LO ( optlc_net_1031 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1033 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1043 ( .LO ( optlc_net_1032 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1034 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1044 ( .LO ( optlc_net_1033 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1035 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1045 ( .LO ( optlc_net_1034 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1036 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1046 ( .LO ( optlc_net_1035 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1037 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1047 ( .LO ( optlc_net_1036 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1038 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1048 ( .LO ( optlc_net_1037 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1039 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1049 ( .LO ( optlc_net_1038 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1040 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1050 ( .LO ( optlc_net_1039 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1041 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1051 ( .LO ( optlc_net_1040 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1042 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1052 ( .LO ( optlc_net_1041 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1043 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1053 ( .LO ( optlc_net_1042 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1044 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1054 ( .LO ( optlc_net_1043 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1045 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1055 ( .LO ( optlc_net_1044 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1046 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1056 ( .LO ( optlc_net_1045 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1047 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1057 ( .LO ( optlc_net_1046 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1048 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1058 ( .LO ( optlc_net_1047 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1049 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1059 ( .LO ( optlc_net_1048 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1050 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1060 ( .LO ( optlc_net_1049 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1051 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1061 ( .LO ( optlc_net_1050 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1052 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1062 ( .LO ( optlc_net_1051 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1053 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1063 ( .LO ( optlc_net_1052 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1054 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1064 ( .LO ( optlc_net_1053 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1055 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1065 ( .LO ( optlc_net_1054 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1056 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1066 ( .LO ( optlc_net_1055 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1057 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1067 ( .LO ( optlc_net_1056 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1058 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1068 ( .LO ( optlc_net_1057 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1059 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1069 ( .LO ( optlc_net_1058 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1060 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1070 ( .LO ( optlc_net_1059 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1061 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1071 ( .LO ( optlc_net_1060 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1062 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1072 ( .LO ( optlc_net_1061 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1063 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1073 ( .LO ( optlc_net_1062 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1064 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1074 ( .LO ( optlc_net_1063 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1065 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1075 ( .LO ( optlc_net_1064 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1066 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1076 ( .LO ( optlc_net_1065 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1067 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1077 ( .LO ( optlc_net_1066 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1068 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1078 ( .LO ( optlc_net_1067 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1069 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1079 ( .LO ( optlc_net_1068 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1070 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1080 ( .LO ( optlc_net_1069 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1071 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1081 ( .LO ( optlc_net_1070 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1072 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1082 ( .LO ( optlc_net_1071 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1073 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1083 ( .LO ( optlc_net_1072 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1074 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1084 ( .LO ( optlc_net_1073 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1075 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1085 ( .LO ( optlc_net_1074 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1076 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1086 ( .LO ( optlc_net_1075 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1077 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1087 ( .LO ( optlc_net_1076 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1078 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1088 ( .LO ( optlc_net_1077 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1079 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1089 ( .LO ( optlc_net_1078 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1080 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1090 ( .LO ( optlc_net_1079 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1081 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1091 ( .LO ( optlc_net_1080 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1082 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1092 ( .LO ( optlc_net_1081 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1083 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1093 ( .LO ( optlc_net_1082 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1084 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1094 ( .LO ( optlc_net_1083 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1085 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1095 ( .LO ( optlc_net_1084 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1086 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1096 ( .LO ( optlc_net_1085 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1087 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1098 ( .LO ( optlc_net_1086 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1088 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1099 ( .LO ( optlc_net_1087 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1089 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1100 ( .LO ( optlc_net_1088 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1090 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1101 ( .LO ( optlc_net_1089 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1091 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1102 ( .LO ( optlc_net_1090 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1092 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1103 ( .LO ( optlc_net_1091 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1093 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1104 ( .LO ( optlc_net_1092 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1094 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1105 ( .LO ( optlc_net_1093 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1095 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1106 ( .LO ( optlc_net_1094 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1096 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1107 ( .LO ( optlc_net_1095 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1097 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1108 ( .LO ( optlc_net_1096 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1098 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1109 ( .LO ( optlc_net_1097 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1099 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1110 ( .LO ( optlc_net_1098 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1100 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1111 ( .LO ( optlc_net_1099 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1101 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1112 ( .LO ( optlc_net_1100 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1102 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1113 ( .LO ( optlc_net_1101 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1103 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1114 ( .LO ( optlc_net_1102 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1104 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1115 ( .LO ( optlc_net_1103 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1105 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1116 ( .LO ( optlc_net_1104 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1106 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1117 ( .LO ( optlc_net_1105 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1107 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1119 ( .LO ( optlc_net_1106 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1108 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1120 ( .LO ( optlc_net_1107 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1109 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1121 ( .LO ( optlc_net_1108 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1110 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1122 ( .LO ( optlc_net_1109 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1111 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1123 ( .LO ( optlc_net_1110 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1112 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1125 ( .LO ( optlc_net_1111 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1113 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1126 ( .LO ( optlc_net_1112 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1114 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1127 ( .LO ( optlc_net_1113 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1115 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1128 ( .LO ( optlc_net_1114 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1116 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1129 ( .LO ( optlc_net_1115 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1117 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1130 ( .LO ( optlc_net_1116 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1118 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1131 ( .LO ( optlc_net_1117 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1119 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1132 ( .LO ( optlc_net_1118 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1120 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1133 ( .LO ( optlc_net_1119 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1121 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1134 ( .LO ( optlc_net_1120 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1122 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1135 ( .LO ( optlc_net_1121 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1123 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1136 ( .LO ( optlc_net_1122 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1124 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1137 ( .LO ( optlc_net_1123 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1125 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1138 ( .LO ( optlc_net_1124 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1126 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1139 ( .LO ( optlc_net_1125 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1127 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1140 ( .LO ( optlc_net_1126 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1128 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1141 ( .LO ( optlc_net_1127 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1129 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1142 ( .LO ( optlc_net_1128 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1130 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1143 ( .LO ( optlc_net_1129 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1131 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1144 ( .LO ( optlc_net_1130 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1132 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1145 ( .LO ( optlc_net_1131 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1133 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1146 ( .LO ( optlc_net_1132 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1134 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1148 ( .LO ( optlc_net_1133 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1135 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1149 ( .LO ( optlc_net_1134 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1136 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1150 ( .LO ( optlc_net_1135 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1137 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1151 ( .LO ( optlc_net_1136 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1138 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1152 ( .LO ( optlc_net_1137 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1139 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1153 ( .LO ( optlc_net_1138 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1140 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1154 ( .LO ( optlc_net_1139 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1141 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1156 ( .LO ( optlc_net_1140 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1142 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1158 ( .LO ( optlc_net_1141 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1143 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1159 ( .LO ( optlc_net_1142 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1144 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1160 ( .LO ( optlc_net_1143 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1145 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1161 ( .LO ( optlc_net_1144 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1146 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1162 ( .LO ( optlc_net_1145 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1147 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1163 ( .LO ( optlc_net_1146 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1148 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1164 ( .LO ( optlc_net_1147 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1149 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1165 ( .LO ( optlc_net_1148 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1150 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1166 ( .LO ( optlc_net_1149 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1151 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1167 ( .LO ( optlc_net_1150 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1152 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1168 ( .LO ( optlc_net_1151 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1153 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1169 ( .LO ( optlc_net_1152 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1154 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1170 ( .LO ( optlc_net_1153 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1155 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1171 ( .LO ( optlc_net_1154 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1156 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1172 ( .LO ( optlc_net_1155 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1157 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1174 ( .LO ( optlc_net_1156 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1158 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1175 ( .LO ( optlc_net_1157 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1159 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1176 ( .LO ( optlc_net_1158 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1160 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1177 ( .LO ( optlc_net_1159 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1161 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1178 ( .LO ( optlc_net_1160 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1162 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1179 ( .LO ( optlc_net_1161 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1163 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1180 ( .LO ( optlc_net_1162 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1164 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1181 ( .LO ( optlc_net_1163 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1165 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1182 ( .LO ( optlc_net_1164 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1166 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1183 ( .LO ( optlc_net_1165 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1167 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1184 ( .LO ( optlc_net_1166 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1168 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1185 ( .LO ( optlc_net_1167 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1169 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1186 ( .LO ( optlc_net_1168 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1170 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1187 ( .LO ( optlc_net_1169 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1171 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1188 ( .LO ( optlc_net_1170 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1172 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1189 ( .LO ( optlc_net_1171 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1173 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1190 ( .LO ( optlc_net_1172 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1174 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1191 ( .LO ( optlc_net_1173 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1175 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1192 ( .LO ( optlc_net_1174 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1176 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1193 ( .LO ( optlc_net_1175 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1177 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1194 ( .LO ( optlc_net_1176 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1178 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1195 ( .LO ( optlc_net_1177 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1179 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1196 ( .LO ( optlc_net_1178 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1180 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1197 ( .LO ( optlc_net_1179 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1181 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1198 ( .LO ( optlc_net_1180 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1182 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1199 ( .LO ( optlc_net_1181 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1183 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1200 ( .LO ( optlc_net_1182 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1184 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1201 ( .LO ( optlc_net_1183 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1185 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1202 ( .LO ( optlc_net_1184 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1186 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1203 ( .LO ( optlc_net_1185 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1187 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1204 ( .LO ( optlc_net_1186 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1188 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1205 ( .LO ( optlc_net_1187 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1189 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1206 ( .LO ( optlc_net_1188 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1190 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1207 ( .LO ( optlc_net_1189 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1191 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1208 ( .LO ( optlc_net_1190 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1192 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1209 ( .LO ( optlc_net_1191 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1193 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1210 ( .LO ( optlc_net_1192 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1194 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1211 ( .LO ( optlc_net_1193 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1195 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1213 ( .LO ( optlc_net_1194 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1196 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1214 ( .LO ( optlc_net_1195 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1197 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1215 ( .LO ( optlc_net_1196 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1198 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1216 ( .LO ( optlc_net_1197 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1199 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1217 ( .LO ( optlc_net_1198 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1200 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1219 ( .LO ( optlc_net_1199 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1201 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1220 ( .LO ( optlc_net_1200 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1202 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1222 ( .LO ( optlc_net_1201 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1203 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1223 ( .LO ( optlc_net_1202 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1204 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1224 ( .LO ( optlc_net_1203 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1205 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1225 ( .LO ( optlc_net_1204 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1206 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1226 ( .LO ( optlc_net_1205 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1207 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1227 ( .LO ( optlc_net_1206 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1208 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1228 ( .LO ( optlc_net_1207 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1209 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1229 ( .LO ( optlc_net_1208 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1210 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1230 ( .LO ( optlc_net_1209 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1211 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1232 ( .LO ( optlc_net_1210 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1212 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1233 ( .LO ( optlc_net_1211 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1213 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1234 ( .LO ( optlc_net_1212 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1214 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1235 ( .LO ( optlc_net_1213 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1215 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1236 ( .LO ( optlc_net_1214 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1216 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1237 ( .LO ( optlc_net_1215 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1217 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1238 ( .LO ( optlc_net_1216 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1218 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1239 ( .LO ( optlc_net_1217 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1219 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1240 ( .LO ( optlc_net_1218 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1220 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1241 ( .LO ( optlc_net_1219 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1221 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1242 ( .LO ( optlc_net_1220 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1222 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1243 ( .LO ( optlc_net_1221 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1223 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1244 ( .LO ( optlc_net_1222 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1224 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1246 ( .LO ( optlc_net_1223 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1225 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1247 ( .LO ( optlc_net_1224 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1226 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1248 ( .LO ( optlc_net_1225 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1227 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1249 ( .LO ( optlc_net_1226 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1228 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1250 ( .LO ( optlc_net_1227 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1229 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1251 ( .LO ( optlc_net_1228 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1230 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1252 ( .LO ( optlc_net_1229 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1231 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1254 ( .LO ( optlc_net_1230 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1232 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1255 ( .LO ( optlc_net_1231 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1233 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1256 ( .LO ( optlc_net_1232 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1234 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1257 ( .LO ( optlc_net_1233 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1235 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1258 ( .LO ( optlc_net_1234 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1236 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1259 ( .LO ( optlc_net_1235 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1237 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1261 ( .LO ( optlc_net_1236 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1238 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1262 ( .LO ( optlc_net_1237 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1239 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1263 ( .LO ( optlc_net_1238 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1240 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1264 ( .LO ( optlc_net_1239 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1241 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1266 ( .LO ( optlc_net_1240 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1242 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1267 ( .LO ( optlc_net_1241 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1243 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1268 ( .LO ( optlc_net_1242 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1244 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1269 ( .LO ( optlc_net_1243 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1245 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1271 ( .LO ( optlc_net_1244 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1246 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1272 ( .LO ( optlc_net_1245 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1247 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1273 ( .LO ( optlc_net_1246 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1248 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1274 ( .LO ( optlc_net_1247 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1249 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1275 ( .LO ( optlc_net_1248 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1250 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1277 ( .LO ( optlc_net_1249 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1251 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1278 ( .LO ( optlc_net_1250 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1252 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1279 ( .LO ( optlc_net_1251 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1253 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1280 ( .LO ( optlc_net_1252 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1254 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1281 ( .LO ( optlc_net_1253 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1255 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1282 ( .LO ( optlc_net_1254 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1256 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1284 ( .LO ( optlc_net_1255 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1257 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1285 ( .LO ( optlc_net_1256 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1258 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1286 ( .LO ( optlc_net_1257 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1259 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1287 ( .LO ( optlc_net_1258 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1260 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1289 ( .LO ( optlc_net_1259 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1261 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1290 ( .LO ( optlc_net_1260 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1262 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1291 ( .LO ( optlc_net_1261 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1263 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1292 ( .LO ( optlc_net_1262 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1264 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1293 ( .LO ( optlc_net_1263 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1265 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1294 ( .LO ( optlc_net_1264 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1266 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1295 ( .LO ( optlc_net_1265 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1267 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1296 ( .LO ( optlc_net_1266 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1268 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1297 ( .LO ( optlc_net_1267 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1269 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1298 ( .LO ( optlc_net_1268 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1270 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1299 ( .LO ( optlc_net_1269 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1271 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1300 ( .LO ( optlc_net_1270 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1272 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1301 ( .LO ( optlc_net_1271 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1273 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1302 ( .LO ( optlc_net_1272 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1274 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1304 ( .LO ( optlc_net_1273 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1275 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1305 ( .LO ( optlc_net_1274 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1276 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1306 ( .LO ( optlc_net_1275 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1277 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1307 ( .LO ( optlc_net_1276 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1278 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1308 ( .LO ( optlc_net_1277 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1279 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1309 ( .LO ( optlc_net_1278 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1280 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1311 ( .LO ( optlc_net_1279 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1281 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1312 ( .LO ( optlc_net_1280 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1282 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1313 ( .LO ( optlc_net_1281 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1283 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1314 ( .LO ( optlc_net_1282 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1284 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1315 ( .LO ( optlc_net_1283 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1285 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1316 ( .LO ( optlc_net_1284 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1286 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1317 ( .LO ( optlc_net_1285 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1287 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1318 ( .LO ( optlc_net_1286 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1288 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1320 ( .LO ( optlc_net_1287 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1289 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1321 ( .LO ( optlc_net_1288 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1290 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1322 ( .LO ( optlc_net_1289 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1291 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1323 ( .LO ( optlc_net_1290 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1292 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1324 ( .LO ( optlc_net_1291 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1293 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1326 ( .LO ( optlc_net_1292 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1294 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1327 ( .LO ( optlc_net_1293 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1295 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1328 ( .LO ( optlc_net_1294 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1296 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1329 ( .LO ( optlc_net_1295 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1297 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1331 ( .LO ( optlc_net_1296 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1298 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1332 ( .LO ( optlc_net_1297 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1299 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1333 ( .LO ( optlc_net_1298 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1300 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1334 ( .LO ( optlc_net_1299 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1301 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1335 ( .LO ( optlc_net_1300 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1302 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1336 ( .LO ( optlc_net_1301 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1303 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1337 ( .LO ( optlc_net_1302 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1304 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1338 ( .LO ( optlc_net_1303 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1305 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1339 ( .LO ( optlc_net_1304 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1306 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1340 ( .LO ( optlc_net_1305 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1307 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1341 ( .LO ( optlc_net_1306 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1308 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1342 ( .LO ( optlc_net_1307 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1309 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1344 ( .LO ( optlc_net_1308 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1310 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1345 ( .LO ( optlc_net_1309 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1311 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1346 ( .LO ( optlc_net_1310 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1312 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1347 ( .LO ( optlc_net_1311 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1313 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1349 ( .LO ( optlc_net_1312 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1314 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1350 ( .LO ( optlc_net_1313 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1315 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1351 ( .LO ( optlc_net_1314 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1316 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1353 ( .LO ( optlc_net_1315 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1317 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1355 ( .LO ( optlc_net_1316 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1318 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1357 ( .LO ( optlc_net_1317 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1319 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1358 ( .LO ( optlc_net_1318 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1320 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1360 ( .LO ( optlc_net_1319 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1321 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1361 ( .LO ( optlc_net_1320 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1322 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1362 ( .LO ( optlc_net_1321 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1323 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1363 ( .LO ( optlc_net_1322 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1324 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1364 ( .LO ( optlc_net_1323 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1325 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1365 ( .LO ( optlc_net_1324 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1326 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1366 ( .LO ( optlc_net_1325 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1327 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1368 ( .LO ( optlc_net_1326 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1328 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1369 ( .LO ( optlc_net_1327 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1329 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1370 ( .LO ( optlc_net_1328 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1330 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1372 ( .LO ( optlc_net_1329 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1331 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1374 ( .LO ( optlc_net_1330 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1332 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1375 ( .LO ( optlc_net_1331 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1333 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1376 ( .LO ( optlc_net_1332 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1334 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1377 ( .LO ( optlc_net_1333 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1335 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1378 ( .LO ( optlc_net_1334 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1336 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1379 ( .LO ( optlc_net_1335 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1337 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1380 ( .LO ( optlc_net_1336 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1338 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1382 ( .LO ( optlc_net_1337 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1339 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1383 ( .LO ( optlc_net_1338 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1340 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1384 ( .LO ( optlc_net_1339 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1341 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1385 ( .LO ( optlc_net_1340 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1342 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1386 ( .LO ( optlc_net_1341 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1343 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1387 ( .LO ( optlc_net_1342 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1344 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1388 ( .LO ( optlc_net_1343 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1345 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1389 ( .LO ( optlc_net_1344 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1346 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1390 ( .LO ( optlc_net_1345 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1347 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1391 ( .LO ( optlc_net_1346 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1348 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1392 ( .LO ( optlc_net_1347 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1349 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1394 ( .LO ( optlc_net_1348 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1350 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1396 ( .LO ( optlc_net_1349 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1351 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1398 ( .LO ( optlc_net_1350 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1352 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1399 ( .LO ( optlc_net_1351 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1353 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1400 ( .LO ( optlc_net_1352 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1354 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1401 ( .LO ( optlc_net_1353 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1355 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1402 ( .LO ( optlc_net_1354 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1356 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1404 ( .LO ( optlc_net_1355 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1357 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1405 ( .LO ( optlc_net_1356 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1358 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1407 ( .LO ( optlc_net_1357 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1359 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1409 ( .LO ( optlc_net_1358 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1360 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1410 ( .LO ( optlc_net_1359 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1361 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1411 ( .LO ( optlc_net_1360 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1362 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1412 ( .LO ( optlc_net_1361 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1363 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1413 ( .LO ( optlc_net_1362 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1364 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1414 ( .LO ( optlc_net_1363 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1365 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1415 ( .LO ( optlc_net_1364 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1366 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1416 ( .LO ( optlc_net_1365 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1367 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1418 ( .LO ( optlc_net_1366 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1368 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1420 ( .LO ( optlc_net_1367 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1369 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1422 ( .LO ( optlc_net_1368 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1370 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1423 ( .LO ( optlc_net_1369 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1371 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1425 ( .LO ( optlc_net_1370 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1372 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1426 ( .LO ( optlc_net_1371 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1373 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1427 ( .LO ( optlc_net_1372 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1374 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1428 ( .LO ( optlc_net_1373 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1375 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1429 ( .LO ( optlc_net_1374 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1376 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1430 ( .LO ( optlc_net_1375 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1377 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1431 ( .LO ( optlc_net_1376 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1378 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1432 ( .LO ( optlc_net_1377 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1379 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1434 ( .LO ( optlc_net_1378 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1380 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1435 ( .LO ( optlc_net_1379 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1381 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1436 ( .LO ( optlc_net_1380 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1382 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1438 ( .LO ( optlc_net_1381 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1383 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1440 ( .LO ( optlc_net_1382 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1384 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1441 ( .LO ( optlc_net_1383 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1385 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1443 ( .LO ( optlc_net_1384 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1386 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1444 ( .LO ( optlc_net_1385 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1387 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1445 ( .LO ( optlc_net_1386 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1388 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1447 ( .LO ( optlc_net_1387 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1389 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1449 ( .LO ( optlc_net_1388 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1390 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1450 ( .LO ( optlc_net_1389 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1391 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1451 ( .LO ( optlc_net_1390 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1392 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1452 ( .LO ( optlc_net_1391 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1393 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1453 ( .LO ( optlc_net_1392 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1394 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1455 ( .LO ( optlc_net_1393 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1395 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1457 ( .LO ( optlc_net_1394 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1396 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1458 ( .LO ( optlc_net_1395 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1397 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1459 ( .LO ( optlc_net_1396 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1398 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1460 ( .LO ( optlc_net_1397 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1399 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1461 ( .LO ( optlc_net_1398 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1400 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1463 ( .LO ( optlc_net_1399 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1401 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1464 ( .LO ( optlc_net_1400 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1402 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1465 ( .LO ( optlc_net_1401 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1403 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1467 ( .LO ( optlc_net_1402 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1404 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1468 ( .LO ( optlc_net_1403 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1405 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1469 ( .LO ( optlc_net_1404 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1406 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1471 ( .LO ( optlc_net_1405 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1407 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1472 ( .LO ( optlc_net_1406 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1408 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1474 ( .LO ( optlc_net_1407 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1409 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1475 ( .LO ( optlc_net_1408 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1410 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1477 ( .LO ( optlc_net_1409 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1411 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1478 ( .LO ( optlc_net_1410 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1412 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1479 ( .LO ( optlc_net_1411 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1413 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1480 ( .LO ( optlc_net_1412 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1414 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1482 ( .LO ( optlc_net_1413 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1415 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1484 ( .LO ( optlc_net_1414 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1416 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1486 ( .LO ( optlc_net_1415 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1417 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1488 ( .LO ( optlc_net_1416 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1418 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1489 ( .LO ( optlc_net_1417 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1419 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1490 ( .LO ( optlc_net_1418 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1420 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1491 ( .LO ( optlc_net_1419 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1421 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1493 ( .LO ( optlc_net_1420 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1422 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1494 ( .LO ( optlc_net_1421 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1423 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1495 ( .LO ( optlc_net_1422 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1424 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1497 ( .LO ( optlc_net_1423 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1425 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1498 ( .LO ( optlc_net_1424 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1426 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1500 ( .LO ( optlc_net_1425 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1427 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1501 ( .LO ( optlc_net_1426 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1428 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1502 ( .LO ( optlc_net_1427 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1429 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1503 ( .LO ( optlc_net_1428 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1430 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1504 ( .LO ( optlc_net_1429 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1431 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1505 ( .LO ( optlc_net_1430 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1432 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1507 ( .LO ( optlc_net_1431 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1433 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1508 ( .LO ( optlc_net_1432 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1434 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1510 ( .LO ( optlc_net_1433 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1435 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1511 ( .LO ( optlc_net_1434 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1436 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1512 ( .LO ( optlc_net_1435 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1437 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1514 ( .LO ( optlc_net_1436 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1438 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1515 ( .LO ( optlc_net_1437 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1439 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1516 ( .LO ( optlc_net_1438 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1440 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1517 ( .LO ( optlc_net_1439 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1441 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1519 ( .LO ( optlc_net_1440 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1442 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1521 ( .LO ( optlc_net_1441 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1443 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1522 ( .LO ( optlc_net_1442 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1444 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1523 ( .LO ( optlc_net_1443 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1445 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1525 ( .LO ( optlc_net_1444 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1446 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1526 ( .LO ( optlc_net_1445 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1447 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1527 ( .LO ( optlc_net_1446 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1448 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1528 ( .LO ( optlc_net_1447 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1449 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1529 ( .LO ( optlc_net_1448 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1450 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1530 ( .LO ( optlc_net_1449 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1451 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1531 ( .LO ( optlc_net_1450 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1452 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1533 ( .LO ( optlc_net_1451 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1453 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1534 ( .LO ( optlc_net_1452 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1454 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1535 ( .LO ( optlc_net_1453 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1455 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1536 ( .LO ( optlc_net_1454 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1456 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1538 ( .LO ( optlc_net_1455 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1457 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1539 ( .LO ( optlc_net_1456 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1458 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1541 ( .LO ( optlc_net_1457 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1459 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1542 ( .LO ( optlc_net_1458 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1460 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1543 ( .LO ( optlc_net_1459 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1461 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1544 ( .LO ( optlc_net_1460 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1462 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1546 ( .LO ( optlc_net_1461 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1463 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1548 ( .LO ( optlc_net_1462 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1464 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1550 ( .LO ( optlc_net_1463 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1465 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1551 ( .LO ( optlc_net_1464 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1466 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1552 ( .LO ( optlc_net_1465 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1467 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1553 ( .LO ( optlc_net_1466 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1468 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1555 ( .LO ( optlc_net_1467 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1469 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1557 ( .LO ( optlc_net_1468 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1470 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1558 ( .LO ( optlc_net_1469 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1471 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1559 ( .LO ( optlc_net_1470 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1472 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1561 ( .LO ( optlc_net_1471 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1473 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1562 ( .LO ( optlc_net_1472 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1474 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1563 ( .LO ( optlc_net_1473 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1475 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1564 ( .LO ( optlc_net_1474 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1476 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1565 ( .LO ( optlc_net_1475 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1477 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1566 ( .LO ( optlc_net_1476 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1478 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1567 ( .LO ( optlc_net_1477 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1479 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1569 ( .LO ( optlc_net_1478 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1480 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1570 ( .LO ( optlc_net_1479 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1481 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1572 ( .LO ( optlc_net_1480 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1482 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1574 ( .LO ( optlc_net_1481 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1483 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1575 ( .LO ( optlc_net_1482 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1484 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1577 ( .LO ( optlc_net_1483 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1485 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1579 ( .LO ( optlc_net_1484 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1486 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1580 ( .LO ( optlc_net_1485 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1487 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1581 ( .LO ( optlc_net_1486 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1488 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1582 ( .LO ( optlc_net_1487 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1489 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1583 ( .LO ( optlc_net_1488 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1490 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1584 ( .LO ( optlc_net_1489 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1491 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1586 ( .LO ( optlc_net_1490 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1492 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1588 ( .LO ( optlc_net_1491 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1493 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1589 ( .LO ( optlc_net_1492 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1494 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1590 ( .LO ( optlc_net_1493 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1495 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1592 ( .LO ( optlc_net_1494 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1496 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1593 ( .LO ( optlc_net_1495 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1497 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1595 ( .LO ( optlc_net_1496 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1498 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1597 ( .LO ( optlc_net_1497 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1499 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1598 ( .LO ( optlc_net_1498 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1500 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1600 ( .LO ( optlc_net_1499 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1501 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1601 ( .LO ( optlc_net_1500 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1502 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1602 ( .LO ( optlc_net_1501 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1503 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1603 ( .LO ( optlc_net_1502 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1504 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1604 ( .LO ( optlc_net_1503 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1505 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1606 ( .LO ( optlc_net_1504 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1506 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1607 ( .LO ( optlc_net_1505 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1507 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1608 ( .LO ( optlc_net_1506 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1508 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1610 ( .LO ( optlc_net_1507 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1509 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1612 ( .LO ( optlc_net_1508 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1510 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1613 ( .LO ( optlc_net_1509 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1511 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1614 ( .LO ( optlc_net_1510 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1512 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1616 ( .LO ( optlc_net_1511 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1513 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1618 ( .LO ( optlc_net_1512 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1514 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1620 ( .LO ( optlc_net_1513 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1515 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1621 ( .LO ( optlc_net_1514 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1516 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1622 ( .LO ( optlc_net_1515 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1517 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1623 ( .LO ( optlc_net_1516 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1518 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1625 ( .LO ( optlc_net_1517 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1519 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1627 ( .LO ( optlc_net_1518 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1520 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1629 ( .LO ( optlc_net_1519 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1521 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1630 ( .LO ( optlc_net_1520 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1522 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1631 ( .LO ( optlc_net_1521 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1523 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1633 ( .LO ( optlc_net_1522 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1524 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1635 ( .LO ( optlc_net_1523 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1525 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1636 ( .LO ( optlc_net_1524 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1526 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1637 ( .LO ( optlc_net_1525 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1527 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1639 ( .LO ( optlc_net_1526 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1528 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1641 ( .LO ( optlc_net_1527 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1529 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1642 ( .LO ( optlc_net_1528 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1530 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1644 ( .LO ( optlc_net_1529 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1531 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1645 ( .LO ( optlc_net_1530 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1532 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1646 ( .LO ( optlc_net_1531 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1533 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1647 ( .LO ( optlc_net_1532 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1534 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1648 ( .LO ( optlc_net_1533 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1535 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1650 ( .LO ( optlc_net_1534 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1536 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1651 ( .LO ( optlc_net_1535 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1537 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1652 ( .LO ( optlc_net_1536 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1538 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1653 ( .LO ( optlc_net_1537 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1539 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1655 ( .LO ( optlc_net_1538 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1540 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1656 ( .LO ( optlc_net_1539 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1541 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1658 ( .LO ( optlc_net_1540 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1542 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1660 ( .LO ( optlc_net_1541 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1543 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1662 ( .LO ( optlc_net_1542 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1544 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1664 ( .LO ( optlc_net_1543 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1545 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1665 ( .LO ( optlc_net_1544 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1546 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1667 ( .LO ( optlc_net_1545 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1547 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1668 ( .LO ( optlc_net_1546 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1548 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1670 ( .LO ( optlc_net_1547 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1549 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1671 ( .LO ( optlc_net_1548 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1550 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1673 ( .LO ( optlc_net_1549 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1551 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1674 ( .LO ( optlc_net_1550 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1552 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1676 ( .LO ( optlc_net_1551 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1553 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1678 ( .LO ( optlc_net_1552 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1554 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1679 ( .LO ( optlc_net_1553 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1555 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1680 ( .LO ( optlc_net_1554 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1556 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1681 ( .LO ( optlc_net_1555 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1557 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1683 ( .LO ( optlc_net_1556 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1558 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1685 ( .LO ( optlc_net_1557 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1559 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1686 ( .LO ( optlc_net_1558 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1560 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1688 ( .LO ( optlc_net_1559 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1561 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1689 ( .LO ( optlc_net_1560 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1562 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1690 ( .LO ( optlc_net_1561 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1563 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1691 ( .LO ( optlc_net_1562 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1564 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1693 ( .LO ( optlc_net_1563 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1565 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1694 ( .LO ( optlc_net_1564 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1566 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1695 ( .LO ( optlc_net_1565 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1567 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1696 ( .LO ( optlc_net_1566 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1568 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1698 ( .LO ( optlc_net_1567 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1569 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1700 ( .LO ( optlc_net_1568 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1570 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1701 ( .LO ( optlc_net_1569 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1571 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1703 ( .LO ( optlc_net_1570 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1572 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1704 ( .LO ( optlc_net_1571 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1573 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1705 ( .LO ( optlc_net_1572 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1574 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1707 ( .LO ( optlc_net_1573 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1575 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1709 ( .LO ( optlc_net_1574 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1576 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1711 ( .LO ( optlc_net_1575 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1577 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1713 ( .LO ( optlc_net_1576 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1578 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1715 ( .LO ( optlc_net_1577 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1579 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1717 ( .LO ( optlc_net_1578 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1580 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1719 ( .LO ( optlc_net_1579 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1581 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1720 ( .LO ( optlc_net_1580 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1582 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1721 ( .LO ( optlc_net_1581 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1583 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1723 ( .LO ( optlc_net_1582 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1584 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1725 ( .LO ( optlc_net_1583 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1585 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1727 ( .LO ( optlc_net_1584 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1586 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1729 ( .LO ( optlc_net_1585 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1587 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1730 ( .LO ( optlc_net_1586 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1588 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1732 ( .LO ( optlc_net_1587 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1589 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1734 ( .LO ( optlc_net_1588 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1590 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1735 ( .LO ( optlc_net_1589 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1591 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1736 ( .LO ( optlc_net_1590 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1592 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1738 ( .LO ( optlc_net_1591 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1593 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1740 ( .LO ( optlc_net_1592 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1594 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1742 ( .LO ( optlc_net_1593 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1595 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1743 ( .LO ( optlc_net_1594 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1596 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1745 ( .LO ( optlc_net_1595 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1597 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1746 ( .LO ( optlc_net_1596 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1598 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1747 ( .LO ( optlc_net_1597 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1599 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1748 ( .LO ( optlc_net_1598 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1600 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1750 ( .LO ( optlc_net_1599 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1601 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1752 ( .LO ( optlc_net_1600 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1602 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1754 ( .LO ( optlc_net_1601 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1603 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1755 ( .LO ( optlc_net_1602 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1604 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1757 ( .LO ( optlc_net_1603 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1605 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1759 ( .LO ( optlc_net_1604 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1606 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1760 ( .LO ( optlc_net_1605 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1607 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1762 ( .LO ( optlc_net_1606 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1608 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1763 ( .LO ( optlc_net_1607 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1609 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1764 ( .LO ( optlc_net_1608 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1610 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1765 ( .LO ( optlc_net_1609 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1611 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1767 ( .LO ( optlc_net_1610 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1612 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1768 ( .LO ( optlc_net_1611 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1613 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1769 ( .LO ( optlc_net_1612 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1614 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1770 ( .LO ( optlc_net_1613 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1615 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1772 ( .LO ( optlc_net_1614 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1616 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1774 ( .LO ( optlc_net_1615 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1617 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1776 ( .LO ( optlc_net_1616 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1618 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1778 ( .LO ( optlc_net_1617 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1619 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1780 ( .LO ( optlc_net_1618 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1620 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1781 ( .LO ( optlc_net_1619 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1621 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1782 ( .LO ( optlc_net_1620 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1622 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1783 ( .LO ( optlc_net_1621 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1623 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1785 ( .LO ( optlc_net_1622 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1624 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1786 ( .LO ( optlc_net_1623 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1625 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1787 ( .LO ( optlc_net_1624 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1626 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1788 ( .LO ( optlc_net_1625 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1627 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1789 ( .LO ( optlc_net_1626 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1628 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1790 ( .LO ( optlc_net_1627 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1629 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1791 ( .LO ( optlc_net_1628 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1630 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1792 ( .LO ( optlc_net_1629 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1631 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1793 ( .LO ( optlc_net_1630 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1632 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1794 ( .LO ( optlc_net_1631 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1633 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1796 ( .LO ( optlc_net_1632 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1634 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1798 ( .LO ( optlc_net_1633 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1635 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1800 ( .LO ( optlc_net_1634 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1636 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1802 ( .LO ( optlc_net_1635 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1637 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1804 ( .LO ( optlc_net_1636 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1638 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1806 ( .LO ( optlc_net_1637 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1639 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1807 ( .LO ( optlc_net_1638 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1640 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1808 ( .LO ( optlc_net_1639 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1641 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1810 ( .LO ( optlc_net_1640 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1642 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1811 ( .LO ( optlc_net_1641 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1643 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1812 ( .LO ( optlc_net_1642 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1644 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1813 ( .LO ( optlc_net_1643 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1645 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1814 ( .LO ( optlc_net_1644 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1646 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1815 ( .LO ( optlc_net_1645 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1647 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1816 ( .LO ( optlc_net_1646 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1648 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1817 ( .LO ( optlc_net_1647 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1649 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1818 ( .LO ( optlc_net_1648 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1650 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1819 ( .LO ( optlc_net_1649 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1651 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1820 ( .LO ( optlc_net_1650 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1652 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1821 ( .LO ( optlc_net_1651 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1653 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1822 ( .LO ( optlc_net_1652 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1654 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1823 ( .LO ( optlc_net_1653 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1655 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1824 ( .LO ( optlc_net_1654 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1656 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1825 ( .LO ( optlc_net_1655 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1657 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1826 ( .LO ( optlc_net_1656 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1658 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1827 ( .LO ( optlc_net_1657 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1659 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1828 ( .LO ( optlc_net_1658 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1660 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1829 ( .LO ( optlc_net_1659 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1661 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1830 ( .LO ( optlc_net_1660 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1662 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1831 ( .LO ( optlc_net_1661 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1663 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1832 ( .LO ( optlc_net_1662 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1664 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1833 ( .LO ( optlc_net_1663 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1665 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1834 ( .LO ( optlc_net_1664 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1666 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1835 ( .LO ( optlc_net_1665 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1667 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1836 ( .LO ( optlc_net_1666 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1668 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1837 ( .LO ( optlc_net_1667 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1669 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1838 ( .LO ( optlc_net_1668 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1670 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1839 ( .LO ( optlc_net_1669 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1671 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1840 ( .LO ( optlc_net_1670 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1672 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1841 ( .LO ( optlc_net_1671 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1673 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1842 ( .LO ( optlc_net_1672 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1674 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1843 ( .LO ( optlc_net_1673 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1675 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1844 ( .LO ( optlc_net_1674 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1676 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1845 ( .LO ( optlc_net_1675 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1677 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1846 ( .LO ( optlc_net_1676 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1678 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1847 ( .LO ( optlc_net_1677 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1679 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1848 ( .LO ( optlc_net_1678 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1680 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1849 ( .LO ( optlc_net_1679 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1681 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1850 ( .LO ( optlc_net_1680 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1682 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1851 ( .LO ( optlc_net_1681 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1683 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1852 ( .LO ( optlc_net_1682 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1684 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1853 ( .LO ( optlc_net_1683 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1685 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1854 ( .LO ( optlc_net_1684 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1686 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1855 ( .LO ( optlc_net_1685 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1687 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1856 ( .LO ( optlc_net_1686 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1688 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1857 ( .LO ( optlc_net_1687 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1689 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1858 ( .LO ( optlc_net_1688 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1690 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1859 ( .LO ( optlc_net_1689 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1691 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1860 ( .LO ( optlc_net_1690 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1692 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1861 ( .LO ( optlc_net_1691 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1693 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1862 ( .LO ( optlc_net_1692 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1694 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1863 ( .LO ( optlc_net_1693 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1695 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1864 ( .LO ( optlc_net_1694 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1696 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1865 ( .LO ( optlc_net_1695 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1697 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1866 ( .LO ( optlc_net_1696 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1698 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1867 ( .LO ( optlc_net_1697 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1699 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1868 ( .LO ( optlc_net_1698 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1700 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1869 ( .LO ( optlc_net_1699 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1701 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1870 ( .LO ( optlc_net_1700 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1702 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1871 ( .LO ( optlc_net_1701 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1703 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1872 ( .LO ( optlc_net_1702 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1704 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1873 ( .LO ( optlc_net_1703 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1705 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1874 ( .LO ( optlc_net_1704 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1706 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1875 ( .LO ( optlc_net_1705 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1707 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1876 ( .LO ( optlc_net_1706 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1708 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1877 ( .LO ( optlc_net_1707 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1709 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1878 ( .LO ( optlc_net_1708 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1710 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1879 ( .LO ( optlc_net_1709 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1711 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1880 ( .LO ( optlc_net_1710 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1712 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1881 ( .LO ( optlc_net_1711 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1713 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1883 ( .LO ( optlc_net_1712 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1714 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1884 ( .LO ( optlc_net_1713 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1715 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1885 ( .LO ( optlc_net_1714 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1716 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1886 ( .LO ( optlc_net_1715 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1717 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1887 ( .LO ( optlc_net_1716 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1718 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1888 ( .LO ( optlc_net_1717 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1719 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1889 ( .LO ( optlc_net_1718 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1720 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1890 ( .LO ( optlc_net_1719 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1721 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1891 ( .LO ( optlc_net_1720 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1722 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1892 ( .LO ( optlc_net_1721 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1723 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1893 ( .LO ( optlc_net_1722 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1724 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1894 ( .LO ( optlc_net_1723 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1725 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1895 ( .LO ( optlc_net_1724 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1726 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1896 ( .LO ( optlc_net_1725 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1727 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1897 ( .LO ( optlc_net_1726 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1728 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1898 ( .LO ( optlc_net_1727 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1729 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1899 ( .LO ( optlc_net_1728 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1730 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1900 ( .LO ( optlc_net_1729 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1731 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1901 ( .LO ( optlc_net_1730 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1732 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1902 ( .LO ( optlc_net_1731 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1733 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1903 ( .LO ( optlc_net_1732 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1734 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1904 ( .LO ( optlc_net_1733 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1735 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1905 ( .LO ( optlc_net_1734 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1736 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1906 ( .LO ( optlc_net_1735 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1737 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1907 ( .LO ( optlc_net_1736 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1738 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1908 ( .LO ( optlc_net_1737 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1739 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1909 ( .LO ( optlc_net_1738 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1740 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1910 ( .LO ( optlc_net_1739 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1741 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1911 ( .LO ( optlc_net_1740 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1742 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1912 ( .LO ( optlc_net_1741 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1743 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1913 ( .LO ( optlc_net_1742 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1744 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1914 ( .LO ( optlc_net_1743 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1745 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1915 ( .LO ( optlc_net_1744 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1746 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1917 ( .LO ( optlc_net_1745 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1747 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1918 ( .LO ( optlc_net_1746 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1748 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1919 ( .LO ( optlc_net_1747 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1749 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1920 ( .LO ( optlc_net_1748 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1750 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1921 ( .LO ( optlc_net_1749 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1751 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1922 ( .LO ( optlc_net_1750 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1752 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1923 ( .LO ( optlc_net_1751 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1753 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1924 ( .LO ( optlc_net_1752 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1754 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1925 ( .LO ( optlc_net_1753 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1755 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1926 ( .LO ( optlc_net_1754 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1756 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1927 ( .LO ( optlc_net_1755 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1757 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1928 ( .LO ( optlc_net_1756 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1758 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1929 ( .LO ( optlc_net_1757 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1759 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1930 ( .LO ( optlc_net_1758 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1760 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1931 ( .LO ( optlc_net_1759 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1761 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1932 ( .LO ( optlc_net_1760 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1762 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1933 ( .LO ( optlc_net_1761 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1763 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1934 ( .LO ( optlc_net_1762 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1764 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1935 ( .LO ( optlc_net_1763 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1765 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1936 ( .LO ( optlc_net_1764 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1766 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1937 ( .LO ( optlc_net_1765 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1767 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1938 ( .LO ( optlc_net_1766 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1768 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1939 ( .LO ( optlc_net_1767 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1769 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1941 ( .LO ( optlc_net_1768 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1770 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1942 ( .LO ( optlc_net_1769 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1771 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1943 ( .LO ( optlc_net_1770 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1772 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1944 ( .LO ( optlc_net_1771 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1773 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1945 ( .LO ( optlc_net_1772 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1774 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1947 ( .LO ( optlc_net_1773 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1775 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1948 ( .LO ( optlc_net_1774 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1776 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1950 ( .LO ( optlc_net_1775 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1777 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1951 ( .LO ( optlc_net_1776 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1778 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1952 ( .LO ( optlc_net_1777 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1779 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1954 ( .LO ( optlc_net_1778 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1780 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1955 ( .LO ( optlc_net_1779 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1781 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1957 ( .LO ( optlc_net_1780 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1782 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1959 ( .LO ( optlc_net_1781 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1783 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1960 ( .LO ( optlc_net_1782 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1784 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1961 ( .LO ( optlc_net_1783 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1785 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1962 ( .LO ( optlc_net_1784 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1786 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1963 ( .LO ( optlc_net_1785 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1787 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1964 ( .LO ( optlc_net_1786 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1788 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1965 ( .LO ( optlc_net_1787 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1789 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1966 ( .LO ( optlc_net_1788 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1790 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1967 ( .LO ( optlc_net_1789 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1791 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1968 ( .LO ( optlc_net_1790 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1792 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1969 ( .LO ( optlc_net_1791 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1793 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1970 ( .LO ( optlc_net_1792 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1794 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1971 ( .LO ( optlc_net_1793 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1795 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1973 ( .LO ( optlc_net_1794 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1796 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1974 ( .LO ( optlc_net_1795 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1797 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1975 ( .LO ( optlc_net_1796 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1798 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1977 ( .LO ( optlc_net_1797 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1799 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1979 ( .LO ( optlc_net_1798 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1800 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1980 ( .LO ( optlc_net_1799 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1801 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1982 ( .LO ( optlc_net_1800 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1802 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1983 ( .LO ( optlc_net_1801 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1803 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1984 ( .LO ( optlc_net_1802 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1804 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1985 ( .LO ( optlc_net_1803 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1805 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1986 ( .LO ( optlc_net_1804 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1806 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1987 ( .LO ( optlc_net_1805 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1807 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1989 ( .LO ( optlc_net_1806 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1808 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1990 ( .LO ( optlc_net_1807 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1809 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1991 ( .LO ( optlc_net_1808 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1810 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1992 ( .LO ( optlc_net_1809 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1811 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1993 ( .LO ( optlc_net_1810 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1812 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1995 ( .LO ( optlc_net_1811 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1813 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1996 ( .LO ( optlc_net_1812 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1814 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1998 ( .LO ( optlc_net_1813 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1815 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_1999 ( .LO ( optlc_net_1814 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1816 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2001 ( .LO ( optlc_net_1815 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1817 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2003 ( .LO ( optlc_net_1816 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1818 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2005 ( .LO ( optlc_net_1817 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1819 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2006 ( .LO ( optlc_net_1818 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1820 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2008 ( .LO ( optlc_net_1819 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1821 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2009 ( .LO ( optlc_net_1820 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1822 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2011 ( .LO ( optlc_net_1821 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1823 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2012 ( .LO ( optlc_net_1822 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1824 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2013 ( .LO ( optlc_net_1823 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1825 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2014 ( .LO ( optlc_net_1824 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1826 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2015 ( .LO ( optlc_net_1825 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1827 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2016 ( .LO ( optlc_net_1826 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1828 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2017 ( .LO ( optlc_net_1827 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1829 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2018 ( .LO ( optlc_net_1828 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1830 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2020 ( .LO ( optlc_net_1829 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1831 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2022 ( .LO ( optlc_net_1830 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1832 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2024 ( .LO ( optlc_net_1831 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1833 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2026 ( .LO ( optlc_net_1832 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1834 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2028 ( .LO ( optlc_net_1833 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1835 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2029 ( .LO ( optlc_net_1834 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1836 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2030 ( .LO ( optlc_net_1835 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1837 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2032 ( .LO ( optlc_net_1836 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1838 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2034 ( .LO ( optlc_net_1837 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1839 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2036 ( .LO ( optlc_net_1838 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1840 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2037 ( .LO ( optlc_net_1839 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1841 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2038 ( .LO ( optlc_net_1840 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1842 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2040 ( .LO ( optlc_net_1841 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1843 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2042 ( .LO ( optlc_net_1842 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1844 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2044 ( .LO ( optlc_net_1843 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1845 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2046 ( .LO ( optlc_net_1844 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1846 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2048 ( .LO ( optlc_net_1845 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1847 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2049 ( .LO ( optlc_net_1846 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1848 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2051 ( .LO ( optlc_net_1847 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1849 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2053 ( .LO ( optlc_net_1848 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1850 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2054 ( .LO ( optlc_net_1849 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1851 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2056 ( .LO ( optlc_net_1850 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1852 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2057 ( .LO ( optlc_net_1851 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1853 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2058 ( .LO ( optlc_net_1852 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1854 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2059 ( .LO ( optlc_net_1853 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1855 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2060 ( .LO ( optlc_net_1854 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1856 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2062 ( .LO ( optlc_net_1855 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1857 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2064 ( .LO ( optlc_net_1856 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1858 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2065 ( .LO ( optlc_net_1857 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1859 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2066 ( .LO ( optlc_net_1858 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1860 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2067 ( .LO ( optlc_net_1859 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1861 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2068 ( .LO ( optlc_net_1860 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1862 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2070 ( .LO ( optlc_net_1861 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1863 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2072 ( .LO ( optlc_net_1862 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1864 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2073 ( .LO ( optlc_net_1863 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1865 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2074 ( .LO ( optlc_net_1864 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1866 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2075 ( .LO ( optlc_net_1865 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1867 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2077 ( .LO ( optlc_net_1866 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1868 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2078 ( .LO ( optlc_net_1867 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1869 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2080 ( .LO ( optlc_net_1868 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1870 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2081 ( .LO ( optlc_net_1869 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1871 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2083 ( .LO ( optlc_net_1870 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1872 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2085 ( .LO ( optlc_net_1871 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1873 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2086 ( .LO ( optlc_net_1872 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1874 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2088 ( .LO ( optlc_net_1873 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1875 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2089 ( .LO ( optlc_net_1874 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1876 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2091 ( .LO ( optlc_net_1875 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1877 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2092 ( .LO ( optlc_net_1876 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1878 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2093 ( .LO ( optlc_net_1877 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1879 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2094 ( .LO ( optlc_net_1878 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1880 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2096 ( .LO ( optlc_net_1879 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1881 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2098 ( .LO ( optlc_net_1880 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1882 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2100 ( .LO ( optlc_net_1881 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1883 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2101 ( .LO ( optlc_net_1882 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1884 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2102 ( .LO ( optlc_net_1883 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1885 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2103 ( .LO ( optlc_net_1884 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1886 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2105 ( .LO ( optlc_net_1885 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1887 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2107 ( .LO ( optlc_net_1886 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1888 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2109 ( .LO ( optlc_net_1887 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1889 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2111 ( .LO ( optlc_net_1888 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1890 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2112 ( .LO ( optlc_net_1889 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1891 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2113 ( .LO ( optlc_net_1890 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1892 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2114 ( .LO ( optlc_net_1891 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1893 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2116 ( .LO ( optlc_net_1892 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1894 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2118 ( .LO ( optlc_net_1893 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1895 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2120 ( .LO ( optlc_net_1894 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1896 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2122 ( .LO ( optlc_net_1895 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1897 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2124 ( .LO ( optlc_net_1896 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1898 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2126 ( .LO ( optlc_net_1897 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1899 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2128 ( .LO ( optlc_net_1898 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1900 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2129 ( .LO ( optlc_net_1899 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1901 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2130 ( .LO ( optlc_net_1900 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1902 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2131 ( .LO ( optlc_net_1901 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1903 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2133 ( .LO ( optlc_net_1902 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1904 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2135 ( .LO ( optlc_net_1903 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1905 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2136 ( .LO ( optlc_net_1904 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1906 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2137 ( .LO ( optlc_net_1905 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1907 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2138 ( .LO ( optlc_net_1906 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1908 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2140 ( .LO ( optlc_net_1907 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1909 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2141 ( .LO ( optlc_net_1908 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1910 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2143 ( .LO ( optlc_net_1909 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1911 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2144 ( .LO ( optlc_net_1910 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1912 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2146 ( .LO ( optlc_net_1911 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1913 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2148 ( .LO ( optlc_net_1912 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1914 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2150 ( .LO ( optlc_net_1913 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1915 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2151 ( .LO ( optlc_net_1914 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1916 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2152 ( .LO ( optlc_net_1915 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1917 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2153 ( .LO ( optlc_net_1916 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1918 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2154 ( .LO ( optlc_net_1917 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1919 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2155 ( .LO ( optlc_net_1918 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1920 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2157 ( .LO ( optlc_net_1919 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1921 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2159 ( .LO ( optlc_net_1920 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1922 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2161 ( .LO ( optlc_net_1921 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1923 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2162 ( .LO ( optlc_net_1922 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1924 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2164 ( .LO ( optlc_net_1923 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1925 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2166 ( .LO ( optlc_net_1924 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1926 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2167 ( .LO ( optlc_net_1925 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1927 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2169 ( .LO ( optlc_net_1926 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1928 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2171 ( .LO ( optlc_net_1927 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1929 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2173 ( .LO ( optlc_net_1928 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1930 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2174 ( .LO ( optlc_net_1929 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1931 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2175 ( .LO ( optlc_net_1930 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1932 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2176 ( .LO ( optlc_net_1931 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1933 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2177 ( .LO ( optlc_net_1932 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1934 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2178 ( .LO ( optlc_net_1933 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1935 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2180 ( .LO ( optlc_net_1934 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1936 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2182 ( .LO ( optlc_net_1935 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1937 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2184 ( .LO ( optlc_net_1936 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1938 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2185 ( .LO ( optlc_net_1937 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1939 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2186 ( .LO ( optlc_net_1938 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1940 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2188 ( .LO ( optlc_net_1939 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1941 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2189 ( .LO ( optlc_net_1940 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1942 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2190 ( .LO ( optlc_net_1941 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1943 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2191 ( .LO ( optlc_net_1942 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1944 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2193 ( .LO ( optlc_net_1943 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1945 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2194 ( .LO ( optlc_net_1944 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1946 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2195 ( .LO ( optlc_net_1945 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1947 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2197 ( .LO ( optlc_net_1946 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1948 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2199 ( .LO ( optlc_net_1947 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1949 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2200 ( .LO ( optlc_net_1948 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1950 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2201 ( .LO ( optlc_net_1949 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1951 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2202 ( .LO ( optlc_net_1950 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1952 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2204 ( .LO ( optlc_net_1951 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1953 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2206 ( .LO ( optlc_net_1952 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1954 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2207 ( .LO ( optlc_net_1953 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1955 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2209 ( .LO ( optlc_net_1954 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1956 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2210 ( .LO ( optlc_net_1955 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1957 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2212 ( .LO ( optlc_net_1956 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1958 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2214 ( .LO ( optlc_net_1957 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1959 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2215 ( .LO ( optlc_net_1958 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1960 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2217 ( .LO ( optlc_net_1959 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1961 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2218 ( .LO ( optlc_net_1960 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1962 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2220 ( .LO ( optlc_net_1961 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1963 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2222 ( .LO ( optlc_net_1962 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1964 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2224 ( .LO ( optlc_net_1963 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1965 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2225 ( .LO ( optlc_net_1964 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1966 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2226 ( .LO ( optlc_net_1965 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1967 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2227 ( .LO ( optlc_net_1966 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1968 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2229 ( .LO ( optlc_net_1967 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1969 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2231 ( .LO ( optlc_net_1968 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1970 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2233 ( .LO ( optlc_net_1969 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1971 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2235 ( .LO ( optlc_net_1970 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1972 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2236 ( .LO ( optlc_net_1971 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1973 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2237 ( .LO ( optlc_net_1972 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1974 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2238 ( .LO ( optlc_net_1973 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1975 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2239 ( .LO ( optlc_net_1974 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1976 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2240 ( .LO ( optlc_net_1975 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1977 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2242 ( .LO ( optlc_net_1976 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1978 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2243 ( .LO ( optlc_net_1977 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1979 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2245 ( .LO ( optlc_net_1978 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1980 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2247 ( .LO ( optlc_net_1979 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1981 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2248 ( .LO ( optlc_net_1980 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1982 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2250 ( .LO ( optlc_net_1981 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1983 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2251 ( .LO ( optlc_net_1982 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1984 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2253 ( .LO ( optlc_net_1983 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1985 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2254 ( .LO ( optlc_net_1984 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1986 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2255 ( .LO ( optlc_net_1985 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1987 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2256 ( .LO ( optlc_net_1986 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1988 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2257 ( .LO ( optlc_net_1987 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1989 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2258 ( .LO ( optlc_net_1988 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1990 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2259 ( .LO ( optlc_net_1989 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1991 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2260 ( .LO ( optlc_net_1990 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1992 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2261 ( .LO ( optlc_net_1991 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1993 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2262 ( .LO ( optlc_net_1992 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1994 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2263 ( .LO ( optlc_net_1993 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1995 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2264 ( .LO ( optlc_net_1994 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1996 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2265 ( .LO ( optlc_net_1995 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1997 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2266 ( .LO ( optlc_net_1996 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1998 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2267 ( .LO ( optlc_net_1997 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_1999 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2268 ( .LO ( optlc_net_1998 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2000 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2269 ( .LO ( optlc_net_1999 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2001 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2270 ( .LO ( optlc_net_2000 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2002 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2271 ( .LO ( optlc_net_2001 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2003 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2272 ( .LO ( optlc_net_2002 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2004 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2273 ( .LO ( optlc_net_2003 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2005 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2274 ( .LO ( optlc_net_2004 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2006 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2275 ( .LO ( optlc_net_2005 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2007 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2276 ( .LO ( optlc_net_2006 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2008 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2277 ( .LO ( optlc_net_2007 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2009 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2278 ( .LO ( optlc_net_2008 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2010 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2279 ( .LO ( optlc_net_2009 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2011 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2280 ( .LO ( optlc_net_2010 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2012 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2281 ( .LO ( optlc_net_2011 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2013 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2282 ( .LO ( optlc_net_2012 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2014 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2283 ( .LO ( optlc_net_2013 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2015 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2284 ( .LO ( optlc_net_2014 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2016 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2285 ( .LO ( optlc_net_2015 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2017 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2286 ( .LO ( optlc_net_2016 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2018 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2287 ( .LO ( optlc_net_2017 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2019 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2288 ( .LO ( optlc_net_2018 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2020 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2289 ( .LO ( optlc_net_2019 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2021 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2290 ( .LO ( optlc_net_2020 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2022 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2291 ( .LO ( optlc_net_2021 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2023 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2292 ( .LO ( optlc_net_2022 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2024 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2293 ( .LO ( optlc_net_2023 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2025 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2294 ( .LO ( optlc_net_2024 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2026 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2295 ( .LO ( optlc_net_2025 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2027 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2296 ( .LO ( optlc_net_2026 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2028 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2297 ( .LO ( optlc_net_2027 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2029 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2298 ( .LO ( optlc_net_2028 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2030 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2299 ( .LO ( optlc_net_2029 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2031 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2300 ( .LO ( optlc_net_2030 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2032 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2301 ( .LO ( optlc_net_2031 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2033 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2302 ( .LO ( optlc_net_2032 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2034 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2303 ( .LO ( optlc_net_2033 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2035 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2304 ( .LO ( optlc_net_2034 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2036 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2305 ( .LO ( optlc_net_2035 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2037 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2306 ( .LO ( optlc_net_2036 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2038 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2307 ( .LO ( optlc_net_2037 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2039 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2308 ( .LO ( optlc_net_2038 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2040 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2309 ( .LO ( optlc_net_2039 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2041 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2310 ( .LO ( optlc_net_2040 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2042 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2311 ( .LO ( optlc_net_2041 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2043 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2312 ( .LO ( optlc_net_2042 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2044 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2313 ( .LO ( optlc_net_2043 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2045 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2314 ( .LO ( optlc_net_2044 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2046 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2315 ( .LO ( optlc_net_2045 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2047 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2316 ( .LO ( optlc_net_2046 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2048 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2317 ( .LO ( optlc_net_2047 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2049 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2318 ( .LO ( optlc_net_2048 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2050 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2319 ( .LO ( optlc_net_2049 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2051 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2320 ( .LO ( optlc_net_2050 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2052 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2321 ( .LO ( optlc_net_2051 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2053 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2322 ( .LO ( optlc_net_2052 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2054 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2323 ( .LO ( optlc_net_2053 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2055 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2324 ( .LO ( optlc_net_2054 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2056 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2325 ( .LO ( optlc_net_2055 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2057 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2326 ( .LO ( optlc_net_2056 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2058 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2327 ( .LO ( optlc_net_2057 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2059 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2328 ( .LO ( optlc_net_2058 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2060 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2329 ( .LO ( optlc_net_2059 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2061 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2330 ( .LO ( optlc_net_2060 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2062 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2331 ( .LO ( optlc_net_2061 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2063 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2332 ( .LO ( optlc_net_2062 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2064 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2333 ( .LO ( optlc_net_2063 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2065 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2334 ( .LO ( optlc_net_2064 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2066 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2335 ( .LO ( optlc_net_2065 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2067 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2336 ( .LO ( optlc_net_2066 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2068 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2337 ( .LO ( optlc_net_2067 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2069 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2338 ( .LO ( optlc_net_2068 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2070 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2339 ( .LO ( optlc_net_2069 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2071 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2340 ( .LO ( optlc_net_2070 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2072 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2341 ( .LO ( optlc_net_2071 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2073 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2342 ( .LO ( optlc_net_2072 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2074 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2343 ( .LO ( optlc_net_2073 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2075 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2344 ( .LO ( optlc_net_2074 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2076 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2345 ( .LO ( optlc_net_2075 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2077 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2346 ( .LO ( optlc_net_2076 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2078 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2347 ( .LO ( optlc_net_2077 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2079 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2348 ( .LO ( optlc_net_2078 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2080 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2349 ( .LO ( optlc_net_2079 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2081 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2350 ( .LO ( optlc_net_2080 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2082 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2351 ( .LO ( optlc_net_2081 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2083 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2352 ( .LO ( optlc_net_2082 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2084 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2353 ( .LO ( optlc_net_2083 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2085 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2354 ( .LO ( optlc_net_2084 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2086 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2355 ( .LO ( optlc_net_2085 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2087 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2356 ( .LO ( optlc_net_2086 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2088 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2357 ( .LO ( optlc_net_2087 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2089 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2358 ( .LO ( optlc_net_2088 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2090 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2359 ( .LO ( optlc_net_2089 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2091 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2360 ( .LO ( optlc_net_2090 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2092 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2361 ( .LO ( optlc_net_2091 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2093 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2362 ( .LO ( optlc_net_2092 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2094 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2363 ( .LO ( optlc_net_2093 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2095 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2364 ( .LO ( optlc_net_2094 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2096 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2365 ( .LO ( optlc_net_2095 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2097 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2366 ( .LO ( optlc_net_2096 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2098 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2367 ( .LO ( optlc_net_2097 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2099 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2368 ( .LO ( optlc_net_2098 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2100 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2369 ( .LO ( optlc_net_2099 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2101 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2370 ( .LO ( optlc_net_2100 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2102 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2371 ( .LO ( optlc_net_2101 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2103 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2372 ( .LO ( optlc_net_2102 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2104 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2373 ( .LO ( optlc_net_2103 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2105 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2374 ( .LO ( optlc_net_2104 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2106 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2375 ( .LO ( optlc_net_2105 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2107 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2376 ( .LO ( optlc_net_2106 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2108 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2377 ( .LO ( optlc_net_2107 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2109 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2378 ( .LO ( optlc_net_2108 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2110 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2379 ( .LO ( optlc_net_2109 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2111 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2380 ( .LO ( optlc_net_2110 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2112 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2381 ( .LO ( optlc_net_2111 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2113 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2382 ( .LO ( optlc_net_2112 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2114 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2384 ( .LO ( optlc_net_2113 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2115 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2385 ( .LO ( optlc_net_2114 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2116 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2386 ( .LO ( optlc_net_2115 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2117 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2387 ( .LO ( optlc_net_2116 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2118 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2389 ( .LO ( optlc_net_2117 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2119 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2390 ( .LO ( optlc_net_2118 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2120 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2391 ( .LO ( optlc_net_2119 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2121 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2392 ( .LO ( optlc_net_2120 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2122 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2393 ( .LO ( optlc_net_2121 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2123 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2395 ( .LO ( optlc_net_2122 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2124 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2397 ( .LO ( optlc_net_2123 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2125 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2398 ( .LO ( optlc_net_2124 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2126 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2399 ( .LO ( optlc_net_2125 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2127 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2400 ( .LO ( optlc_net_2126 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2128 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2402 ( .LO ( optlc_net_2127 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2129 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2403 ( .LO ( optlc_net_2128 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2130 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2405 ( .LO ( optlc_net_2129 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2131 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2407 ( .LO ( optlc_net_2130 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2132 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2408 ( .LO ( optlc_net_2131 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2133 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2410 ( .LO ( optlc_net_2132 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2134 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2412 ( .LO ( optlc_net_2133 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2135 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2413 ( .LO ( optlc_net_2134 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2136 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2415 ( .LO ( optlc_net_2135 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2137 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2416 ( .LO ( optlc_net_2136 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2138 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2418 ( .LO ( optlc_net_2137 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2139 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2420 ( .LO ( optlc_net_2138 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2140 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2421 ( .LO ( optlc_net_2139 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2141 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2422 ( .LO ( optlc_net_2140 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2142 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2423 ( .LO ( optlc_net_2141 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2143 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2424 ( .LO ( optlc_net_2142 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2144 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2425 ( .LO ( optlc_net_2143 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2145 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2426 ( .LO ( optlc_net_2144 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2146 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2428 ( .LO ( optlc_net_2145 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2147 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2430 ( .LO ( optlc_net_2146 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2148 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2431 ( .LO ( optlc_net_2147 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2149 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2433 ( .LO ( optlc_net_2148 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2150 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2434 ( .LO ( optlc_net_2149 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2151 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2435 ( .LO ( optlc_net_2150 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2152 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2437 ( .LO ( optlc_net_2151 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2153 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2438 ( .LO ( optlc_net_2152 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2154 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2439 ( .LO ( optlc_net_2153 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2155 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2441 ( .LO ( optlc_net_2154 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2156 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2442 ( .LO ( optlc_net_2155 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2157 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2443 ( .LO ( optlc_net_2156 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2158 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2444 ( .LO ( optlc_net_2157 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2159 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2446 ( .LO ( optlc_net_2158 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2160 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2447 ( .LO ( optlc_net_2159 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2161 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2449 ( .LO ( optlc_net_2160 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2162 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2450 ( .LO ( optlc_net_2161 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2163 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2452 ( .LO ( optlc_net_2162 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2164 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2454 ( .LO ( optlc_net_2163 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2165 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2455 ( .LO ( optlc_net_2164 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2166 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2456 ( .LO ( optlc_net_2165 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2167 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2457 ( .LO ( optlc_net_2166 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2168 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2459 ( .LO ( optlc_net_2167 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2169 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2460 ( .LO ( optlc_net_2168 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2170 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2462 ( .LO ( optlc_net_2169 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2171 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2464 ( .LO ( optlc_net_2170 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2172 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2465 ( .LO ( optlc_net_2171 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2173 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2467 ( .LO ( optlc_net_2172 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2174 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2468 ( .LO ( optlc_net_2173 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2175 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2470 ( .LO ( optlc_net_2174 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2176 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2472 ( .LO ( optlc_net_2175 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2177 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2473 ( .LO ( optlc_net_2176 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2178 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2474 ( .LO ( optlc_net_2177 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2179 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2475 ( .LO ( optlc_net_2178 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2180 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2476 ( .LO ( optlc_net_2179 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2181 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2478 ( .LO ( optlc_net_2180 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2182 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2480 ( .LO ( optlc_net_2181 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2183 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2482 ( .LO ( optlc_net_2182 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2184 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2484 ( .LO ( optlc_net_2183 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2185 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2485 ( .LO ( optlc_net_2184 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2186 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2486 ( .LO ( optlc_net_2185 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2187 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2487 ( .LO ( optlc_net_2186 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2188 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2488 ( .LO ( optlc_net_2187 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2189 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2490 ( .LO ( optlc_net_2188 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2190 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2492 ( .LO ( optlc_net_2189 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2191 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2494 ( .LO ( optlc_net_2190 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2192 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2495 ( .LO ( optlc_net_2191 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2193 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2496 ( .LO ( optlc_net_2192 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2194 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2497 ( .LO ( optlc_net_2193 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2195 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2498 ( .LO ( optlc_net_2194 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2196 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2500 ( .LO ( optlc_net_2195 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2197 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2501 ( .LO ( optlc_net_2196 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2198 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2503 ( .LO ( optlc_net_2197 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2199 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2504 ( .LO ( optlc_net_2198 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2200 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2505 ( .LO ( optlc_net_2199 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2201 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2506 ( .LO ( optlc_net_2200 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2202 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2507 ( .LO ( optlc_net_2201 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2203 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2509 ( .LO ( optlc_net_2202 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2204 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2511 ( .LO ( optlc_net_2203 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2205 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2512 ( .LO ( optlc_net_2204 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2206 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2514 ( .LO ( optlc_net_2205 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2207 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2515 ( .LO ( optlc_net_2206 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2208 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2517 ( .LO ( optlc_net_2207 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2209 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2518 ( .LO ( optlc_net_2208 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2210 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2519 ( .LO ( optlc_net_2209 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2211 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2521 ( .LO ( optlc_net_2210 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2212 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2522 ( .LO ( optlc_net_2211 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2213 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2523 ( .LO ( optlc_net_2212 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2214 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2525 ( .LO ( optlc_net_2213 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2215 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2527 ( .LO ( optlc_net_2214 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2216 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2528 ( .LO ( optlc_net_2215 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2217 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2529 ( .LO ( optlc_net_2216 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2218 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2530 ( .LO ( optlc_net_2217 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2219 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2531 ( .LO ( optlc_net_2218 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2220 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2532 ( .LO ( optlc_net_2219 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2221 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2533 ( .LO ( optlc_net_2220 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2222 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2534 ( .LO ( optlc_net_2221 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2223 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2536 ( .LO ( optlc_net_2222 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2224 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2537 ( .LO ( optlc_net_2223 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2225 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2539 ( .LO ( optlc_net_2224 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2226 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2540 ( .LO ( optlc_net_2225 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2227 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2541 ( .LO ( optlc_net_2226 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2228 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2543 ( .LO ( optlc_net_2227 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2229 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2544 ( .LO ( optlc_net_2228 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2230 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2546 ( .LO ( optlc_net_2229 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2231 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2547 ( .LO ( optlc_net_2230 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2232 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2548 ( .LO ( optlc_net_2231 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2233 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2549 ( .LO ( optlc_net_2232 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2234 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2550 ( .LO ( optlc_net_2233 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2235 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2551 ( .LO ( optlc_net_2234 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2236 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2552 ( .LO ( optlc_net_2235 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2237 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2553 ( .LO ( optlc_net_2236 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2238 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2554 ( .LO ( optlc_net_2237 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2239 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2556 ( .LO ( optlc_net_2238 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2240 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2557 ( .LO ( optlc_net_2239 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2241 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2558 ( .LO ( optlc_net_2240 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2242 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2559 ( .LO ( optlc_net_2241 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2243 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2560 ( .LO ( optlc_net_2242 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2244 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2562 ( .LO ( optlc_net_2243 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2245 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2563 ( .LO ( optlc_net_2244 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2246 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2564 ( .LO ( optlc_net_2245 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2247 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2566 ( .LO ( optlc_net_2246 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2248 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2568 ( .LO ( optlc_net_2247 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2249 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2569 ( .LO ( optlc_net_2248 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2250 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2570 ( .LO ( optlc_net_2249 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2251 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2571 ( .LO ( optlc_net_2250 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2252 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2572 ( .LO ( optlc_net_2251 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2253 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2573 ( .LO ( optlc_net_2252 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2254 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2574 ( .LO ( optlc_net_2253 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2255 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2575 ( .LO ( optlc_net_2254 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2256 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2577 ( .LO ( optlc_net_2255 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2257 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2578 ( .LO ( optlc_net_2256 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2258 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2579 ( .LO ( optlc_net_2257 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2259 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2580 ( .LO ( optlc_net_2258 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2260 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2582 ( .LO ( optlc_net_2259 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2261 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2584 ( .LO ( optlc_net_2260 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2262 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2586 ( .LO ( optlc_net_2261 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2263 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2588 ( .LO ( optlc_net_2262 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2264 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2589 ( .LO ( optlc_net_2263 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2265 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2590 ( .LO ( optlc_net_2264 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2266 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2591 ( .LO ( optlc_net_2265 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2267 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2592 ( .LO ( optlc_net_2266 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2268 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2593 ( .LO ( optlc_net_2267 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2269 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2595 ( .LO ( optlc_net_2268 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2270 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2596 ( .LO ( optlc_net_2269 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2271 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2598 ( .LO ( optlc_net_2270 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2272 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2599 ( .LO ( optlc_net_2271 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2273 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2600 ( .LO ( optlc_net_2272 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2274 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2601 ( .LO ( optlc_net_2273 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2275 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2603 ( .LO ( optlc_net_2274 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2276 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2604 ( .LO ( optlc_net_2275 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2277 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2605 ( .LO ( optlc_net_2276 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2278 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2606 ( .LO ( optlc_net_2277 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2279 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2607 ( .LO ( optlc_net_2278 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2280 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2608 ( .LO ( optlc_net_2279 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2281 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2609 ( .LO ( optlc_net_2280 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2282 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2610 ( .LO ( optlc_net_2281 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2283 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2611 ( .LO ( optlc_net_2282 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2284 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2613 ( .LO ( optlc_net_2283 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2285 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2614 ( .LO ( optlc_net_2284 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2286 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2615 ( .LO ( optlc_net_2285 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2287 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2617 ( .LO ( optlc_net_2286 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2288 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2619 ( .LO ( optlc_net_2287 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2289 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2620 ( .LO ( optlc_net_2288 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2290 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2621 ( .LO ( optlc_net_2289 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2291 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2622 ( .LO ( optlc_net_2290 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2292 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2623 ( .LO ( optlc_net_2291 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2293 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2624 ( .LO ( optlc_net_2292 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2294 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2625 ( .LO ( optlc_net_2293 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2295 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2626 ( .LO ( optlc_net_2294 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2296 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2627 ( .LO ( optlc_net_2295 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2297 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2628 ( .LO ( optlc_net_2296 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2298 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2629 ( .LO ( optlc_net_2297 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2299 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2630 ( .LO ( optlc_net_2298 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2300 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2631 ( .LO ( optlc_net_2299 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2301 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2632 ( .LO ( optlc_net_2300 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2302 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2633 ( .LO ( optlc_net_2301 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2303 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2634 ( .LO ( optlc_net_2302 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2304 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2635 ( .LO ( optlc_net_2303 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2305 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2636 ( .LO ( optlc_net_2304 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2306 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2637 ( .LO ( optlc_net_2305 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2307 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2638 ( .LO ( optlc_net_2306 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2308 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2639 ( .LO ( optlc_net_2307 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2309 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2640 ( .LO ( optlc_net_2308 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2310 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2641 ( .LO ( optlc_net_2309 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2311 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2642 ( .LO ( optlc_net_2310 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2312 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2643 ( .LO ( optlc_net_2311 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2313 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2644 ( .LO ( optlc_net_2312 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2314 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2645 ( .LO ( optlc_net_2313 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2315 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2646 ( .LO ( optlc_net_2314 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2316 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2647 ( .LO ( optlc_net_2315 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2317 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2648 ( .LO ( optlc_net_2316 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2318 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2649 ( .LO ( optlc_net_2317 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2319 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2650 ( .LO ( optlc_net_2318 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2320 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2651 ( .LO ( optlc_net_2319 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2321 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2652 ( .LO ( optlc_net_2320 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2322 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2653 ( .LO ( optlc_net_2321 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2323 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2654 ( .LO ( optlc_net_2322 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2324 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2655 ( .LO ( optlc_net_2323 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2325 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2656 ( .LO ( optlc_net_2324 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2326 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2657 ( .LO ( optlc_net_2325 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2327 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2658 ( .LO ( optlc_net_2326 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2328 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2659 ( .LO ( optlc_net_2327 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2329 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2660 ( .LO ( optlc_net_2328 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2330 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2661 ( .LO ( optlc_net_2329 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2331 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2662 ( .LO ( optlc_net_2330 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2332 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2663 ( .LO ( optlc_net_2331 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2333 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2664 ( .LO ( optlc_net_2332 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2334 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2665 ( .LO ( optlc_net_2333 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2335 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2666 ( .LO ( optlc_net_2334 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2336 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2667 ( .LO ( optlc_net_2335 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2337 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2668 ( .LO ( optlc_net_2336 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2338 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2669 ( .LO ( optlc_net_2337 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2339 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2670 ( .LO ( optlc_net_2338 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2340 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2671 ( .LO ( optlc_net_2339 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2341 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2672 ( .LO ( optlc_net_2340 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2342 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2673 ( .LO ( optlc_net_2341 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2343 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2674 ( .LO ( optlc_net_2342 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2344 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2675 ( .LO ( optlc_net_2343 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2345 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2676 ( .LO ( optlc_net_2344 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2346 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2677 ( .LO ( optlc_net_2345 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2347 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2678 ( .LO ( optlc_net_2346 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2348 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2679 ( .LO ( optlc_net_2347 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2349 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2680 ( .LO ( optlc_net_2348 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2350 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2681 ( .LO ( optlc_net_2349 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2351 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2682 ( .LO ( optlc_net_2350 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2352 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2683 ( .LO ( optlc_net_2351 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2353 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2684 ( .LO ( optlc_net_2352 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2354 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2685 ( .LO ( optlc_net_2353 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2355 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2686 ( .LO ( optlc_net_2354 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2356 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2687 ( .LO ( optlc_net_2355 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2357 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2688 ( .LO ( optlc_net_2356 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2358 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2689 ( .LO ( optlc_net_2357 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2359 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2690 ( .LO ( optlc_net_2358 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2360 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2691 ( .LO ( optlc_net_2359 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2361 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2692 ( .LO ( optlc_net_2360 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2362 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2693 ( .LO ( optlc_net_2361 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2363 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2694 ( .LO ( optlc_net_2362 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2364 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2695 ( .LO ( optlc_net_2363 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2365 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2696 ( .LO ( optlc_net_2364 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2366 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2697 ( .LO ( optlc_net_2365 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2367 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2698 ( .LO ( optlc_net_2366 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2368 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2699 ( .LO ( optlc_net_2367 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2369 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2700 ( .LO ( optlc_net_2368 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2370 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2701 ( .LO ( optlc_net_2369 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2371 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2702 ( .LO ( optlc_net_2370 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2372 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2703 ( .LO ( optlc_net_2371 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2373 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2704 ( .LO ( optlc_net_2372 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2374 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2705 ( .LO ( optlc_net_2373 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2375 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2706 ( .LO ( optlc_net_2374 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2376 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2707 ( .LO ( optlc_net_2375 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2377 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2708 ( .LO ( optlc_net_2376 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2378 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2709 ( .LO ( optlc_net_2377 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2379 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2710 ( .LO ( optlc_net_2378 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2380 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2711 ( .LO ( optlc_net_2379 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2381 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2712 ( .LO ( optlc_net_2380 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2382 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2713 ( .LO ( optlc_net_2381 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2383 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2714 ( .LO ( optlc_net_2382 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2384 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2715 ( .LO ( optlc_net_2383 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2385 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2716 ( .LO ( optlc_net_2384 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2386 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2717 ( .LO ( optlc_net_2385 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2387 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2718 ( .LO ( optlc_net_2386 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2388 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2719 ( .LO ( optlc_net_2387 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2389 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2720 ( .LO ( optlc_net_2388 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2390 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2721 ( .LO ( optlc_net_2389 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2391 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2722 ( .LO ( optlc_net_2390 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2392 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2723 ( .LO ( optlc_net_2391 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2393 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2724 ( .LO ( optlc_net_2392 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2394 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2725 ( .LO ( optlc_net_2393 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2395 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2726 ( .LO ( optlc_net_2394 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2396 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2727 ( .LO ( optlc_net_2395 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2397 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2728 ( .LO ( optlc_net_2396 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2398 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2729 ( .LO ( optlc_net_2397 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2399 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2730 ( .LO ( optlc_net_2398 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2400 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2731 ( .LO ( optlc_net_2399 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2401 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2732 ( .LO ( optlc_net_2400 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2402 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2733 ( .LO ( optlc_net_2401 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2403 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2734 ( .LO ( optlc_net_2402 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2404 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2735 ( .LO ( optlc_net_2403 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2405 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2736 ( .LO ( optlc_net_2404 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2406 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2737 ( .LO ( optlc_net_2405 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2407 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2738 ( .LO ( optlc_net_2406 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2408 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2740 ( .LO ( optlc_net_2407 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2409 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2741 ( .LO ( optlc_net_2408 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2410 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2742 ( .LO ( optlc_net_2409 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2411 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2743 ( .LO ( optlc_net_2410 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2412 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2744 ( .LO ( optlc_net_2411 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2413 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2745 ( .LO ( optlc_net_2412 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2414 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2746 ( .LO ( optlc_net_2413 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2415 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2748 ( .LO ( optlc_net_2414 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2416 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2749 ( .LO ( optlc_net_2415 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2417 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2750 ( .LO ( optlc_net_2416 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2418 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2751 ( .LO ( optlc_net_2417 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2419 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2752 ( .LO ( optlc_net_2418 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2420 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2753 ( .LO ( optlc_net_2419 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2421 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2754 ( .LO ( optlc_net_2420 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2422 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2755 ( .LO ( optlc_net_2421 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2423 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2757 ( .LO ( optlc_net_2422 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2424 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2758 ( .LO ( optlc_net_2423 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2425 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2759 ( .LO ( optlc_net_2424 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2426 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2760 ( .LO ( optlc_net_2425 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2427 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2761 ( .LO ( optlc_net_2426 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2428 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2763 ( .LO ( optlc_net_2427 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2429 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2765 ( .LO ( optlc_net_2428 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2430 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2767 ( .LO ( optlc_net_2429 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2431 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2768 ( .LO ( optlc_net_2430 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2432 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2769 ( .LO ( optlc_net_2431 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2433 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2770 ( .LO ( optlc_net_2432 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2434 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2771 ( .LO ( optlc_net_2433 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2435 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2772 ( .LO ( optlc_net_2434 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2436 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2773 ( .LO ( optlc_net_2435 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2437 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2775 ( .LO ( optlc_net_2436 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2438 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2777 ( .LO ( optlc_net_2437 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2439 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2779 ( .LO ( optlc_net_2438 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2440 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2780 ( .LO ( optlc_net_2439 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2441 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2781 ( .LO ( optlc_net_2440 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2442 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2783 ( .LO ( optlc_net_2441 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2443 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2785 ( .LO ( optlc_net_2442 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2444 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2786 ( .LO ( optlc_net_2443 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2445 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2788 ( .LO ( optlc_net_2444 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2446 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2789 ( .LO ( optlc_net_2445 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2447 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2791 ( .LO ( optlc_net_2446 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2448 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2792 ( .LO ( optlc_net_2447 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2449 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2793 ( .LO ( optlc_net_2448 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2450 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2794 ( .LO ( optlc_net_2449 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2451 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2795 ( .LO ( optlc_net_2450 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2452 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2796 ( .LO ( optlc_net_2451 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2453 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2798 ( .LO ( optlc_net_2452 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2454 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2799 ( .LO ( optlc_net_2453 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2455 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2800 ( .LO ( optlc_net_2454 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2456 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2801 ( .LO ( optlc_net_2455 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2457 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2802 ( .LO ( optlc_net_2456 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2458 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2804 ( .LO ( optlc_net_2457 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2459 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2806 ( .LO ( optlc_net_2458 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2460 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2808 ( .LO ( optlc_net_2459 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2461 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2810 ( .LO ( optlc_net_2460 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2462 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2811 ( .LO ( optlc_net_2461 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2463 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2813 ( .LO ( optlc_net_2462 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2464 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2815 ( .LO ( optlc_net_2463 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2465 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2817 ( .LO ( optlc_net_2464 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2466 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2819 ( .LO ( optlc_net_2465 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2467 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2820 ( .LO ( optlc_net_2466 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2468 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2821 ( .LO ( optlc_net_2467 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2469 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2822 ( .LO ( optlc_net_2468 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2470 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2823 ( .LO ( optlc_net_2469 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2471 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2825 ( .LO ( optlc_net_2470 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2472 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2827 ( .LO ( optlc_net_2471 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2473 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2828 ( .LO ( optlc_net_2472 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2474 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2830 ( .LO ( optlc_net_2473 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2475 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2832 ( .LO ( optlc_net_2474 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2476 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2834 ( .LO ( optlc_net_2475 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2477 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2835 ( .LO ( optlc_net_2476 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2478 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2836 ( .LO ( optlc_net_2477 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2479 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2837 ( .LO ( optlc_net_2478 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2480 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2838 ( .LO ( optlc_net_2479 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2481 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2840 ( .LO ( optlc_net_2480 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2482 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2841 ( .LO ( optlc_net_2481 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2483 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2842 ( .LO ( optlc_net_2482 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2484 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2844 ( .LO ( optlc_net_2483 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2485 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2845 ( .LO ( optlc_net_2484 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2486 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2847 ( .LO ( optlc_net_2485 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2487 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2849 ( .LO ( optlc_net_2486 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2488 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2851 ( .LO ( optlc_net_2487 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2489 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2852 ( .LO ( optlc_net_2488 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2490 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2853 ( .LO ( optlc_net_2489 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2491 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2854 ( .LO ( optlc_net_2490 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2492 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2855 ( .LO ( optlc_net_2491 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2493 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2856 ( .LO ( optlc_net_2492 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2494 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2858 ( .LO ( optlc_net_2493 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2495 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2859 ( .LO ( optlc_net_2494 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2496 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2861 ( .LO ( optlc_net_2495 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2497 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2862 ( .LO ( optlc_net_2496 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2498 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2863 ( .LO ( optlc_net_2497 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2499 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2864 ( .LO ( optlc_net_2498 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2500 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2865 ( .LO ( optlc_net_2499 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2501 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2867 ( .LO ( optlc_net_2500 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2502 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2868 ( .LO ( optlc_net_2501 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2503 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2869 ( .LO ( optlc_net_2502 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2504 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2870 ( .LO ( optlc_net_2503 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2505 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2871 ( .LO ( optlc_net_2504 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2506 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2872 ( .LO ( optlc_net_2505 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2507 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2873 ( .LO ( optlc_net_2506 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2508 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2874 ( .LO ( optlc_net_2507 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2509 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2876 ( .LO ( optlc_net_2508 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2510 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2877 ( .LO ( optlc_net_2509 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2511 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2878 ( .LO ( optlc_net_2510 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2512 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2879 ( .LO ( optlc_net_2511 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2513 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2880 ( .LO ( optlc_net_2512 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2514 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2881 ( .LO ( optlc_net_2513 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2515 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2883 ( .LO ( optlc_net_2514 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2516 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2885 ( .LO ( optlc_net_2515 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2517 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2887 ( .LO ( optlc_net_2516 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2518 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2889 ( .LO ( optlc_net_2517 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2519 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2890 ( .LO ( optlc_net_2518 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2520 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2891 ( .LO ( optlc_net_2519 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2521 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2893 ( .LO ( optlc_net_2520 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2522 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2894 ( .LO ( optlc_net_2521 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2523 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2895 ( .LO ( optlc_net_2522 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2524 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2896 ( .LO ( optlc_net_2523 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2525 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2898 ( .LO ( optlc_net_2524 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2526 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2900 ( .LO ( optlc_net_2525 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2527 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2901 ( .LO ( optlc_net_2526 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2528 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2903 ( .LO ( optlc_net_2527 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2529 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2904 ( .LO ( optlc_net_2528 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2530 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2905 ( .LO ( optlc_net_2529 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2531 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2906 ( .LO ( optlc_net_2530 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2532 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2908 ( .LO ( optlc_net_2531 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2533 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2910 ( .LO ( optlc_net_2532 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2534 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2912 ( .LO ( optlc_net_2533 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2535 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2914 ( .LO ( optlc_net_2534 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2536 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2916 ( .LO ( optlc_net_2535 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2537 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2917 ( .LO ( optlc_net_2536 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2538 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2918 ( .LO ( optlc_net_2537 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2539 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2919 ( .LO ( optlc_net_2538 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2540 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2920 ( .LO ( optlc_net_2539 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2541 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2921 ( .LO ( optlc_net_2540 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2542 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2922 ( .LO ( optlc_net_2541 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2543 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2924 ( .LO ( optlc_net_2542 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2544 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2925 ( .LO ( optlc_net_2543 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2545 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2926 ( .LO ( optlc_net_2544 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2546 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2927 ( .LO ( optlc_net_2545 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2547 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2928 ( .LO ( optlc_net_2546 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2548 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2929 ( .LO ( optlc_net_2547 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2549 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2930 ( .LO ( optlc_net_2548 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2550 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2931 ( .LO ( optlc_net_2549 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2551 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2932 ( .LO ( optlc_net_2550 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2552 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2933 ( .LO ( optlc_net_2551 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2553 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2934 ( .LO ( optlc_net_2552 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2554 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2935 ( .LO ( optlc_net_2553 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2555 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2936 ( .LO ( optlc_net_2554 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2556 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2937 ( .LO ( optlc_net_2555 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2557 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2938 ( .LO ( optlc_net_2556 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2558 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2939 ( .LO ( optlc_net_2557 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2559 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2940 ( .LO ( optlc_net_2558 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2560 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2941 ( .LO ( optlc_net_2559 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2561 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2942 ( .LO ( optlc_net_2560 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2562 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2943 ( .LO ( optlc_net_2561 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2563 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2944 ( .LO ( optlc_net_2562 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2564 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2945 ( .LO ( optlc_net_2563 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2565 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2946 ( .LO ( optlc_net_2564 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2566 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2947 ( .LO ( optlc_net_2565 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2567 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2948 ( .LO ( optlc_net_2566 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2568 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2949 ( .LO ( optlc_net_2567 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2569 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2950 ( .LO ( optlc_net_2568 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2570 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2951 ( .LO ( optlc_net_2569 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2571 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2952 ( .LO ( optlc_net_2570 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2572 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2953 ( .LO ( optlc_net_2571 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2573 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2954 ( .LO ( optlc_net_2572 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2574 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2955 ( .LO ( optlc_net_2573 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2575 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2956 ( .LO ( optlc_net_2574 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2576 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2957 ( .LO ( optlc_net_2575 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2577 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2958 ( .LO ( optlc_net_2576 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2578 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2959 ( .LO ( optlc_net_2577 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2579 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2960 ( .LO ( optlc_net_2578 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2580 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2961 ( .LO ( optlc_net_2579 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2581 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2962 ( .LO ( optlc_net_2580 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2582 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2963 ( .LO ( optlc_net_2581 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2583 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2964 ( .LO ( optlc_net_2582 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2584 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2965 ( .LO ( optlc_net_2583 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2585 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2966 ( .LO ( optlc_net_2584 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2586 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2967 ( .LO ( optlc_net_2585 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2587 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2968 ( .LO ( optlc_net_2586 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2588 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2969 ( .LO ( optlc_net_2587 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2589 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2970 ( .LO ( optlc_net_2588 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2590 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2971 ( .LO ( optlc_net_2589 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2591 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2972 ( .LO ( optlc_net_2590 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2592 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2973 ( .LO ( optlc_net_2591 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2593 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2974 ( .LO ( optlc_net_2592 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2594 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2975 ( .LO ( optlc_net_2593 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2595 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2976 ( .LO ( optlc_net_2594 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2596 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2977 ( .LO ( optlc_net_2595 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2597 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2978 ( .LO ( optlc_net_2596 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2598 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2979 ( .LO ( optlc_net_2597 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2599 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2980 ( .LO ( optlc_net_2598 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2600 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2981 ( .LO ( optlc_net_2599 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2601 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2982 ( .LO ( optlc_net_2600 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2602 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2983 ( .LO ( optlc_net_2601 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2603 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2984 ( .LO ( optlc_net_2602 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2604 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2985 ( .LO ( optlc_net_2603 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2605 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2986 ( .LO ( optlc_net_2604 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2606 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2987 ( .LO ( optlc_net_2605 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2607 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2988 ( .LO ( optlc_net_2606 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2608 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2989 ( .LO ( optlc_net_2607 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2609 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2990 ( .LO ( optlc_net_2608 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2610 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2991 ( .LO ( optlc_net_2609 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2611 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2992 ( .LO ( optlc_net_2610 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2612 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2993 ( .LO ( optlc_net_2611 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2613 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2994 ( .LO ( optlc_net_2612 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2614 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2995 ( .LO ( optlc_net_2613 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2615 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2996 ( .LO ( optlc_net_2614 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2616 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2997 ( .LO ( optlc_net_2615 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2617 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2998 ( .LO ( optlc_net_2616 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2618 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_2999 ( .LO ( optlc_net_2617 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2619 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3000 ( .LO ( optlc_net_2618 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2620 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3001 ( .LO ( optlc_net_2619 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2621 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3003 ( .LO ( optlc_net_2620 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2622 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3004 ( .LO ( optlc_net_2621 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2623 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3005 ( .LO ( optlc_net_2622 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2624 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3006 ( .LO ( optlc_net_2623 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2625 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3007 ( .LO ( optlc_net_2624 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2626 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3009 ( .LO ( optlc_net_2625 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2627 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3010 ( .LO ( optlc_net_2626 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2628 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3012 ( .LO ( optlc_net_2627 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2629 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3013 ( .LO ( optlc_net_2628 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2630 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3015 ( .LO ( optlc_net_2629 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2631 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3016 ( .LO ( optlc_net_2630 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2632 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3017 ( .LO ( optlc_net_2631 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2633 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3019 ( .LO ( optlc_net_2632 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2634 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3020 ( .LO ( optlc_net_2633 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2635 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3022 ( .LO ( optlc_net_2634 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2636 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3023 ( .LO ( optlc_net_2635 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2637 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3024 ( .LO ( optlc_net_2636 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2638 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3026 ( .LO ( optlc_net_2637 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2639 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3027 ( .LO ( optlc_net_2638 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2640 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3029 ( .LO ( optlc_net_2639 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2641 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3030 ( .LO ( optlc_net_2640 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2642 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3031 ( .LO ( optlc_net_2641 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2643 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3033 ( .LO ( optlc_net_2642 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2644 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3034 ( .LO ( optlc_net_2643 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2645 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3035 ( .LO ( optlc_net_2644 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2646 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3037 ( .LO ( optlc_net_2645 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2647 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3038 ( .LO ( optlc_net_2646 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2648 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3039 ( .LO ( optlc_net_2647 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2649 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3040 ( .LO ( optlc_net_2648 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2650 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3041 ( .LO ( optlc_net_2649 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2651 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3043 ( .LO ( optlc_net_2650 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2652 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3044 ( .LO ( optlc_net_2651 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2653 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3045 ( .LO ( optlc_net_2652 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2654 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3047 ( .LO ( optlc_net_2653 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2655 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3049 ( .LO ( optlc_net_2654 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2656 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3050 ( .LO ( optlc_net_2655 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2657 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3051 ( .LO ( optlc_net_2656 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2658 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3052 ( .LO ( optlc_net_2657 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2659 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3053 ( .LO ( optlc_net_2658 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2660 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3054 ( .LO ( optlc_net_2659 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2661 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3055 ( .LO ( optlc_net_2660 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2662 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3056 ( .LO ( optlc_net_2661 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2663 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3057 ( .LO ( optlc_net_2662 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2664 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3059 ( .LO ( optlc_net_2663 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2665 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3060 ( .LO ( optlc_net_2664 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2666 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3061 ( .LO ( optlc_net_2665 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2667 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3062 ( .LO ( optlc_net_2666 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2668 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3064 ( .LO ( optlc_net_2667 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2669 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3065 ( .LO ( optlc_net_2668 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2670 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3066 ( .LO ( optlc_net_2669 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2671 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3068 ( .LO ( optlc_net_2670 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2672 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3070 ( .LO ( optlc_net_2671 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2673 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3071 ( .LO ( optlc_net_2672 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2674 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3072 ( .LO ( optlc_net_2673 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2675 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3074 ( .LO ( optlc_net_2674 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2676 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3075 ( .LO ( optlc_net_2675 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2677 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3076 ( .LO ( optlc_net_2676 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2678 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3077 ( .LO ( optlc_net_2677 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2679 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3078 ( .LO ( optlc_net_2678 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2680 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3079 ( .LO ( optlc_net_2679 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2681 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3080 ( .LO ( optlc_net_2680 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2682 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3082 ( .LO ( optlc_net_2681 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2683 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3084 ( .LO ( optlc_net_2682 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2684 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3085 ( .LO ( optlc_net_2683 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2685 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3086 ( .LO ( optlc_net_2684 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2686 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3087 ( .LO ( optlc_net_2685 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2687 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3088 ( .LO ( optlc_net_2686 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2688 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3089 ( .LO ( optlc_net_2687 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2689 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3091 ( .LO ( optlc_net_2688 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2690 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3093 ( .LO ( optlc_net_2689 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2691 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3094 ( .LO ( optlc_net_2690 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2692 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3095 ( .LO ( optlc_net_2691 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2693 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3096 ( .LO ( optlc_net_2692 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2694 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3097 ( .LO ( optlc_net_2693 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2695 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3098 ( .LO ( optlc_net_2694 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2696 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3100 ( .LO ( optlc_net_2695 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2697 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3101 ( .LO ( optlc_net_2696 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2698 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3102 ( .LO ( optlc_net_2697 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2699 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3103 ( .LO ( optlc_net_2698 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2700 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3104 ( .LO ( optlc_net_2699 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2701 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3106 ( .LO ( optlc_net_2700 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2702 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3108 ( .LO ( optlc_net_2701 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2703 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3110 ( .LO ( optlc_net_2702 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2704 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3112 ( .LO ( optlc_net_2703 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2705 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3114 ( .LO ( optlc_net_2704 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2706 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3115 ( .LO ( optlc_net_2705 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2707 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3116 ( .LO ( optlc_net_2706 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2708 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3117 ( .LO ( optlc_net_2707 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2709 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3118 ( .LO ( optlc_net_2708 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2710 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3119 ( .LO ( optlc_net_2709 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2711 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3120 ( .LO ( optlc_net_2710 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2712 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3122 ( .LO ( optlc_net_2711 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2713 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3123 ( .LO ( optlc_net_2712 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2714 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3125 ( .LO ( optlc_net_2713 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2715 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3126 ( .LO ( optlc_net_2714 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2716 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3127 ( .LO ( optlc_net_2715 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2717 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3128 ( .LO ( optlc_net_2716 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2718 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3129 ( .LO ( optlc_net_2717 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2719 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3131 ( .LO ( optlc_net_2718 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2720 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3132 ( .LO ( optlc_net_2719 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2721 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3133 ( .LO ( optlc_net_2720 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2722 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3135 ( .LO ( optlc_net_2721 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2723 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3136 ( .LO ( optlc_net_2722 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2724 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3137 ( .LO ( optlc_net_2723 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2725 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3138 ( .LO ( optlc_net_2724 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2726 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3139 ( .LO ( optlc_net_2725 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2727 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3140 ( .LO ( optlc_net_2726 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2728 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3141 ( .LO ( optlc_net_2727 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2729 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3143 ( .LO ( optlc_net_2728 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2730 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3144 ( .LO ( optlc_net_2729 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2731 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3145 ( .LO ( optlc_net_2730 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2732 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3146 ( .LO ( optlc_net_2731 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2733 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3147 ( .LO ( optlc_net_2732 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2734 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3148 ( .LO ( optlc_net_2733 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2735 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3149 ( .LO ( optlc_net_2734 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2736 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3150 ( .LO ( optlc_net_2735 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2737 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3151 ( .LO ( optlc_net_2736 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2738 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3152 ( .LO ( optlc_net_2737 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2739 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3153 ( .LO ( optlc_net_2738 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2740 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3154 ( .LO ( optlc_net_2739 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2741 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3155 ( .LO ( optlc_net_2740 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2742 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3156 ( .LO ( optlc_net_2741 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2743 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3157 ( .LO ( optlc_net_2742 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2744 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3158 ( .LO ( optlc_net_2743 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2745 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3159 ( .LO ( optlc_net_2744 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2746 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3160 ( .LO ( optlc_net_2745 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2747 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3161 ( .LO ( optlc_net_2746 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2748 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3162 ( .LO ( optlc_net_2747 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2749 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3163 ( .LO ( optlc_net_2748 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2750 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3164 ( .LO ( optlc_net_2749 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2751 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3165 ( .LO ( optlc_net_2750 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2752 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3166 ( .LO ( optlc_net_2751 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2753 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3167 ( .LO ( optlc_net_2752 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2754 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3168 ( .LO ( optlc_net_2753 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2755 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3169 ( .LO ( optlc_net_2754 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2756 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3170 ( .LO ( optlc_net_2755 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2757 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3171 ( .LO ( optlc_net_2756 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2758 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3172 ( .LO ( optlc_net_2757 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2759 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3173 ( .LO ( optlc_net_2758 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2760 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3174 ( .LO ( optlc_net_2759 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2761 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3175 ( .LO ( optlc_net_2760 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2762 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3176 ( .LO ( optlc_net_2761 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2763 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3177 ( .LO ( optlc_net_2762 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2764 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3178 ( .LO ( optlc_net_2763 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2765 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3179 ( .LO ( optlc_net_2764 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2766 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3180 ( .LO ( optlc_net_2765 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2767 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3181 ( .LO ( optlc_net_2766 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2768 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3182 ( .LO ( optlc_net_2767 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2769 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3183 ( .LO ( optlc_net_2768 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2770 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3184 ( .LO ( optlc_net_2769 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2771 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3185 ( .LO ( optlc_net_2770 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2772 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3186 ( .LO ( optlc_net_2771 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2773 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3187 ( .LO ( optlc_net_2772 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2774 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3188 ( .LO ( optlc_net_2773 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2775 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3189 ( .LO ( optlc_net_2774 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2776 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3190 ( .LO ( optlc_net_2775 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2777 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3191 ( .LO ( optlc_net_2776 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2778 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3192 ( .LO ( optlc_net_2777 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2779 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3193 ( .LO ( optlc_net_2778 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2780 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3194 ( .LO ( optlc_net_2779 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2781 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3195 ( .LO ( optlc_net_2780 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2782 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3196 ( .LO ( optlc_net_2781 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2783 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3197 ( .LO ( optlc_net_2782 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2784 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3198 ( .LO ( optlc_net_2783 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2785 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3199 ( .LO ( optlc_net_2784 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2786 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3200 ( .LO ( optlc_net_2785 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2787 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3201 ( .LO ( optlc_net_2786 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2788 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3202 ( .LO ( optlc_net_2787 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2789 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3203 ( .LO ( optlc_net_2788 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2790 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3204 ( .LO ( optlc_net_2789 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2791 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3205 ( .LO ( optlc_net_2790 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2792 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3206 ( .LO ( optlc_net_2791 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2793 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3207 ( .LO ( optlc_net_2792 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2794 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3208 ( .LO ( optlc_net_2793 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2795 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3209 ( .LO ( optlc_net_2794 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2796 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3211 ( .LO ( optlc_net_2795 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2797 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3212 ( .LO ( optlc_net_2796 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2798 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3213 ( .LO ( optlc_net_2797 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2799 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3214 ( .LO ( optlc_net_2798 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2800 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3216 ( .LO ( optlc_net_2799 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2801 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3217 ( .LO ( optlc_net_2800 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2802 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3218 ( .LO ( optlc_net_2801 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2803 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3219 ( .LO ( optlc_net_2802 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2804 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3221 ( .LO ( optlc_net_2803 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2805 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3222 ( .LO ( optlc_net_2804 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2806 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3223 ( .LO ( optlc_net_2805 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2807 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3224 ( .LO ( optlc_net_2806 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2808 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3225 ( .LO ( optlc_net_2807 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2809 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3226 ( .LO ( optlc_net_2808 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2810 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3227 ( .LO ( optlc_net_2809 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2811 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3228 ( .LO ( optlc_net_2810 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2812 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3230 ( .LO ( optlc_net_2811 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2813 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3231 ( .LO ( optlc_net_2812 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2814 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3232 ( .LO ( optlc_net_2813 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2815 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3233 ( .LO ( optlc_net_2814 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2816 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3234 ( .LO ( optlc_net_2815 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2817 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3235 ( .LO ( optlc_net_2816 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2818 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3236 ( .LO ( optlc_net_2817 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2819 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3238 ( .LO ( optlc_net_2818 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2820 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3239 ( .LO ( optlc_net_2819 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2821 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3240 ( .LO ( optlc_net_2820 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2822 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3241 ( .LO ( optlc_net_2821 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2823 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3242 ( .LO ( optlc_net_2822 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2824 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3243 ( .LO ( optlc_net_2823 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2825 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3244 ( .LO ( optlc_net_2824 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2826 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3245 ( .LO ( optlc_net_2825 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2827 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3246 ( .LO ( optlc_net_2826 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2828 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3247 ( .LO ( optlc_net_2827 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2829 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3249 ( .LO ( optlc_net_2828 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2830 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3251 ( .LO ( optlc_net_2829 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2831 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3252 ( .LO ( optlc_net_2830 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2832 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3253 ( .LO ( optlc_net_2831 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2833 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3254 ( .LO ( optlc_net_2832 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2834 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3255 ( .LO ( optlc_net_2833 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2835 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3256 ( .LO ( optlc_net_2834 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2836 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3257 ( .LO ( optlc_net_2835 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2837 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3258 ( .LO ( optlc_net_2836 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2838 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3259 ( .LO ( optlc_net_2837 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2839 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3260 ( .LO ( optlc_net_2838 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2840 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3261 ( .LO ( optlc_net_2839 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2841 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3262 ( .LO ( optlc_net_2840 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2842 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3264 ( .LO ( optlc_net_2841 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2843 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3265 ( .LO ( optlc_net_2842 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2844 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3266 ( .LO ( optlc_net_2843 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2845 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3267 ( .LO ( optlc_net_2844 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2846 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3268 ( .LO ( optlc_net_2845 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2847 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3269 ( .LO ( optlc_net_2846 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2848 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3270 ( .LO ( optlc_net_2847 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2849 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3271 ( .LO ( optlc_net_2848 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2850 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3272 ( .LO ( optlc_net_2849 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2851 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3273 ( .LO ( optlc_net_2850 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2852 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3274 ( .LO ( optlc_net_2851 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2853 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3275 ( .LO ( optlc_net_2852 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2854 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3277 ( .LO ( optlc_net_2853 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2855 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3278 ( .LO ( optlc_net_2854 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2856 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3279 ( .LO ( optlc_net_2855 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2857 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3281 ( .LO ( optlc_net_2856 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2858 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3282 ( .LO ( optlc_net_2857 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2859 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3283 ( .LO ( optlc_net_2858 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2860 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3284 ( .LO ( optlc_net_2859 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2861 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3286 ( .LO ( optlc_net_2860 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2862 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3287 ( .LO ( optlc_net_2861 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2863 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3288 ( .LO ( optlc_net_2862 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2864 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3289 ( .LO ( optlc_net_2863 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2865 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3290 ( .LO ( optlc_net_2864 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2866 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3292 ( .LO ( optlc_net_2865 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2867 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3293 ( .LO ( optlc_net_2866 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2868 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3294 ( .LO ( optlc_net_2867 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2869 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3296 ( .LO ( optlc_net_2868 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2870 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3297 ( .LO ( optlc_net_2869 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2871 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3298 ( .LO ( optlc_net_2870 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2872 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3299 ( .LO ( optlc_net_2871 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2873 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3300 ( .LO ( optlc_net_2872 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2874 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3302 ( .LO ( optlc_net_2873 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2875 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3304 ( .LO ( optlc_net_2874 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2876 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3305 ( .LO ( optlc_net_2875 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2877 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3306 ( .LO ( optlc_net_2876 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2878 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3307 ( .LO ( optlc_net_2877 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2879 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3308 ( .LO ( optlc_net_2878 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2880 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3309 ( .LO ( optlc_net_2879 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2881 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3310 ( .LO ( optlc_net_2880 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2882 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3311 ( .LO ( optlc_net_2881 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2883 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3312 ( .LO ( optlc_net_2882 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2884 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3314 ( .LO ( optlc_net_2883 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2885 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3315 ( .LO ( optlc_net_2884 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2886 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3316 ( .LO ( optlc_net_2885 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2887 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3317 ( .LO ( optlc_net_2886 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2888 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3318 ( .LO ( optlc_net_2887 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2889 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3319 ( .LO ( optlc_net_2888 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2890 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3320 ( .LO ( optlc_net_2889 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2891 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3321 ( .LO ( optlc_net_2890 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2892 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3322 ( .LO ( optlc_net_2891 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2893 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3323 ( .LO ( optlc_net_2892 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2894 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3324 ( .LO ( optlc_net_2893 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2895 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3325 ( .LO ( optlc_net_2894 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2896 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3326 ( .LO ( optlc_net_2895 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2897 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3327 ( .LO ( optlc_net_2896 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2898 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3328 ( .LO ( optlc_net_2897 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2899 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3329 ( .LO ( optlc_net_2898 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2900 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3330 ( .LO ( optlc_net_2899 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2901 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3331 ( .LO ( optlc_net_2900 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2902 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3332 ( .LO ( optlc_net_2901 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2903 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3333 ( .LO ( optlc_net_2902 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2904 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3334 ( .LO ( optlc_net_2903 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2905 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3335 ( .LO ( optlc_net_2904 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2906 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3336 ( .LO ( optlc_net_2905 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2907 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3337 ( .LO ( optlc_net_2906 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2908 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3338 ( .LO ( optlc_net_2907 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2909 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3339 ( .LO ( optlc_net_2908 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2910 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3340 ( .LO ( optlc_net_2909 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2911 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3341 ( .LO ( optlc_net_2910 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2912 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3342 ( .LO ( optlc_net_2911 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2913 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3343 ( .LO ( optlc_net_2912 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2914 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3344 ( .LO ( optlc_net_2913 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2915 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3345 ( .LO ( optlc_net_2914 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2916 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3346 ( .LO ( optlc_net_2915 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2917 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3347 ( .LO ( optlc_net_2916 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2918 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3348 ( .LO ( optlc_net_2917 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2919 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3349 ( .LO ( optlc_net_2918 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2920 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3350 ( .LO ( optlc_net_2919 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2921 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3351 ( .LO ( optlc_net_2920 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2922 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3352 ( .LO ( optlc_net_2921 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2923 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3353 ( .LO ( optlc_net_2922 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2924 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3354 ( .LO ( optlc_net_2923 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2925 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3355 ( .LO ( optlc_net_2924 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2926 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3356 ( .LO ( optlc_net_2925 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2927 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3357 ( .LO ( optlc_net_2926 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2928 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3358 ( .LO ( optlc_net_2927 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2929 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3359 ( .LO ( optlc_net_2928 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2930 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3360 ( .LO ( optlc_net_2929 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2931 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3361 ( .LO ( optlc_net_2930 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2932 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3362 ( .LO ( optlc_net_2931 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2933 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3363 ( .LO ( optlc_net_2932 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2934 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3364 ( .LO ( optlc_net_2933 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2935 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3365 ( .LO ( optlc_net_2934 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2936 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3366 ( .LO ( optlc_net_2935 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2937 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3367 ( .LO ( optlc_net_2936 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2938 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3368 ( .LO ( optlc_net_2937 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2939 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3369 ( .LO ( optlc_net_2938 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2940 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3370 ( .LO ( optlc_net_2939 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2941 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3371 ( .LO ( optlc_net_2940 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2942 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3372 ( .LO ( optlc_net_2941 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2943 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3374 ( .LO ( optlc_net_2942 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2944 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3375 ( .LO ( optlc_net_2943 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2945 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3377 ( .LO ( optlc_net_2944 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2946 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3378 ( .LO ( optlc_net_2945 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2947 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3379 ( .LO ( optlc_net_2946 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2948 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3380 ( .LO ( optlc_net_2947 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2949 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3381 ( .LO ( optlc_net_2948 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2950 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3382 ( .LO ( optlc_net_2949 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2951 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3383 ( .LO ( optlc_net_2950 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2952 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3384 ( .LO ( optlc_net_2951 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2953 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3386 ( .LO ( optlc_net_2952 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2954 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3387 ( .LO ( optlc_net_2953 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2955 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3389 ( .LO ( optlc_net_2954 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2956 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3390 ( .LO ( optlc_net_2955 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2957 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3392 ( .LO ( optlc_net_2956 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2958 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3393 ( .LO ( optlc_net_2957 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2959 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3395 ( .LO ( optlc_net_2958 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2960 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3396 ( .LO ( optlc_net_2959 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2961 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3397 ( .LO ( optlc_net_2960 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2962 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3398 ( .LO ( optlc_net_2961 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2963 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3399 ( .LO ( optlc_net_2962 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2964 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3400 ( .LO ( optlc_net_2963 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2965 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3402 ( .LO ( optlc_net_2964 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2966 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3403 ( .LO ( optlc_net_2965 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2967 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3404 ( .LO ( optlc_net_2966 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2968 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3405 ( .LO ( optlc_net_2967 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2969 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3406 ( .LO ( optlc_net_2968 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2970 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3407 ( .LO ( optlc_net_2969 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2971 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3408 ( .LO ( optlc_net_2970 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2972 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3409 ( .LO ( optlc_net_2971 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2973 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3410 ( .LO ( optlc_net_2972 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2974 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3411 ( .LO ( optlc_net_2973 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2975 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3412 ( .LO ( optlc_net_2974 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2976 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3413 ( .LO ( optlc_net_2975 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2977 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3414 ( .LO ( optlc_net_2976 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2978 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3415 ( .LO ( optlc_net_2977 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2979 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3416 ( .LO ( optlc_net_2978 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2980 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3417 ( .LO ( optlc_net_2979 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2981 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3418 ( .LO ( optlc_net_2980 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2982 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3419 ( .LO ( optlc_net_2981 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2983 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3420 ( .LO ( optlc_net_2982 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2984 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3421 ( .LO ( optlc_net_2983 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2985 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3422 ( .LO ( optlc_net_2984 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2986 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3424 ( .LO ( optlc_net_2985 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2987 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3425 ( .LO ( optlc_net_2986 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2988 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3427 ( .LO ( optlc_net_2987 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2989 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3428 ( .LO ( optlc_net_2988 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2990 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3429 ( .LO ( optlc_net_2989 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2991 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3430 ( .LO ( optlc_net_2990 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2992 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3431 ( .LO ( optlc_net_2991 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2993 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3433 ( .LO ( optlc_net_2992 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2994 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3434 ( .LO ( optlc_net_2993 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2995 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3435 ( .LO ( optlc_net_2994 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2996 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3436 ( .LO ( optlc_net_2995 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2997 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3437 ( .LO ( optlc_net_2996 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2998 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3438 ( .LO ( optlc_net_2997 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_2999 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3439 ( .LO ( optlc_net_2998 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3000 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3440 ( .LO ( optlc_net_2999 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3001 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3441 ( .LO ( optlc_net_3000 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3002 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3443 ( .LO ( optlc_net_3001 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3003 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3444 ( .LO ( optlc_net_3002 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3004 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3445 ( .LO ( optlc_net_3003 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3005 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3446 ( .LO ( optlc_net_3004 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3006 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3447 ( .LO ( optlc_net_3005 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3007 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3448 ( .LO ( optlc_net_3006 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3008 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3449 ( .LO ( optlc_net_3007 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3009 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3451 ( .LO ( optlc_net_3008 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3010 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3453 ( .LO ( optlc_net_3009 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3011 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3454 ( .LO ( optlc_net_3010 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3012 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3455 ( .LO ( optlc_net_3011 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3013 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3457 ( .LO ( optlc_net_3012 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3014 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3458 ( .LO ( optlc_net_3013 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3015 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3459 ( .LO ( optlc_net_3014 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3016 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3460 ( .LO ( optlc_net_3015 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3017 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3461 ( .LO ( optlc_net_3016 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3018 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3462 ( .LO ( optlc_net_3017 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3019 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3463 ( .LO ( optlc_net_3018 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3020 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3464 ( .LO ( optlc_net_3019 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3021 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3465 ( .LO ( optlc_net_3020 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3022 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3466 ( .LO ( optlc_net_3021 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3023 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3467 ( .LO ( optlc_net_3022 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3024 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3468 ( .LO ( optlc_net_3023 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3025 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3469 ( .LO ( optlc_net_3024 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3026 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3470 ( .LO ( optlc_net_3025 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3027 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3471 ( .LO ( optlc_net_3026 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3028 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3472 ( .LO ( optlc_net_3027 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3029 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3473 ( .LO ( optlc_net_3028 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3030 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3474 ( .LO ( optlc_net_3029 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3031 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3475 ( .LO ( optlc_net_3030 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3032 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3476 ( .LO ( optlc_net_3031 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3033 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3477 ( .LO ( optlc_net_3032 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3034 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3478 ( .LO ( optlc_net_3033 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3035 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3479 ( .LO ( optlc_net_3034 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3036 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3480 ( .LO ( optlc_net_3035 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3037 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3481 ( .LO ( optlc_net_3036 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3038 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3482 ( .LO ( optlc_net_3037 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3039 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3483 ( .LO ( optlc_net_3038 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3040 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3484 ( .LO ( optlc_net_3039 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3041 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3485 ( .LO ( optlc_net_3040 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3042 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3486 ( .LO ( optlc_net_3041 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3043 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3487 ( .LO ( optlc_net_3042 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3044 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3488 ( .LO ( optlc_net_3043 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3045 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3489 ( .LO ( optlc_net_3044 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3046 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3490 ( .LO ( optlc_net_3045 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3047 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3491 ( .LO ( optlc_net_3046 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3048 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3492 ( .LO ( optlc_net_3047 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3049 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3493 ( .LO ( optlc_net_3048 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3050 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3494 ( .LO ( optlc_net_3049 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3051 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3495 ( .LO ( optlc_net_3050 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3052 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3496 ( .LO ( optlc_net_3051 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3053 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3497 ( .LO ( optlc_net_3052 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3054 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3498 ( .LO ( optlc_net_3053 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3055 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3499 ( .LO ( optlc_net_3054 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3056 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3500 ( .LO ( optlc_net_3055 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3057 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3501 ( .LO ( optlc_net_3056 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3058 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3502 ( .LO ( optlc_net_3057 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3059 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3503 ( .LO ( optlc_net_3058 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3060 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3504 ( .LO ( optlc_net_3059 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3061 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3505 ( .LO ( optlc_net_3060 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3062 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3506 ( .LO ( optlc_net_3061 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3063 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3507 ( .LO ( optlc_net_3062 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3064 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3508 ( .LO ( optlc_net_3063 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3065 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3509 ( .LO ( optlc_net_3064 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3066 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3511 ( .LO ( optlc_net_3065 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3067 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3512 ( .LO ( optlc_net_3066 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3068 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3513 ( .LO ( optlc_net_3067 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3069 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3514 ( .LO ( optlc_net_3068 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3070 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3515 ( .LO ( optlc_net_3069 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3071 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3516 ( .LO ( optlc_net_3070 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3072 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3517 ( .LO ( optlc_net_3071 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3073 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3518 ( .LO ( optlc_net_3072 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3074 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3519 ( .LO ( optlc_net_3073 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3075 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3520 ( .LO ( optlc_net_3074 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3076 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3521 ( .LO ( optlc_net_3075 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3077 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3522 ( .LO ( optlc_net_3076 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3078 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3523 ( .LO ( optlc_net_3077 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3079 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3524 ( .LO ( optlc_net_3078 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3080 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3525 ( .LO ( optlc_net_3079 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3081 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3526 ( .LO ( optlc_net_3080 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3082 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3527 ( .LO ( optlc_net_3081 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3083 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3529 ( .LO ( optlc_net_3082 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3084 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3530 ( .LO ( optlc_net_3083 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3085 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3531 ( .LO ( optlc_net_3084 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3086 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3532 ( .LO ( optlc_net_3085 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3087 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3533 ( .LO ( optlc_net_3086 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3088 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3534 ( .LO ( optlc_net_3087 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3089 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3535 ( .LO ( optlc_net_3088 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3090 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3537 ( .LO ( optlc_net_3089 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3091 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3538 ( .LO ( optlc_net_3090 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3092 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3539 ( .LO ( optlc_net_3091 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3093 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3541 ( .LO ( optlc_net_3092 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3094 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3543 ( .LO ( optlc_net_3093 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3095 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3544 ( .LO ( optlc_net_3094 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3096 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3545 ( .LO ( optlc_net_3095 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3097 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3546 ( .LO ( optlc_net_3096 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3098 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3547 ( .LO ( optlc_net_3097 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3099 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3549 ( .LO ( optlc_net_3098 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3100 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3550 ( .LO ( optlc_net_3099 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3101 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3551 ( .LO ( optlc_net_3100 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3102 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3552 ( .LO ( optlc_net_3101 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3103 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3554 ( .LO ( optlc_net_3102 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3104 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3555 ( .LO ( optlc_net_3103 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3105 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3556 ( .LO ( optlc_net_3104 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3106 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3557 ( .LO ( optlc_net_3105 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3107 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3558 ( .LO ( optlc_net_3106 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3108 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3559 ( .LO ( optlc_net_3107 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3109 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3560 ( .LO ( optlc_net_3108 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3110 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3561 ( .LO ( optlc_net_3109 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3111 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3562 ( .LO ( optlc_net_3110 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3112 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3563 ( .LO ( optlc_net_3111 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3113 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3564 ( .LO ( optlc_net_3112 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3114 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3565 ( .LO ( optlc_net_3113 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3115 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3567 ( .LO ( optlc_net_3114 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3116 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3568 ( .LO ( optlc_net_3115 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3117 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3569 ( .LO ( optlc_net_3116 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3118 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3570 ( .LO ( optlc_net_3117 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3119 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3571 ( .LO ( optlc_net_3118 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3120 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3573 ( .LO ( optlc_net_3119 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3121 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3574 ( .LO ( optlc_net_3120 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3122 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3575 ( .LO ( optlc_net_3121 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3123 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3576 ( .LO ( optlc_net_3122 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3124 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3577 ( .LO ( optlc_net_3123 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3125 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3578 ( .LO ( optlc_net_3124 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3126 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3579 ( .LO ( optlc_net_3125 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3127 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3580 ( .LO ( optlc_net_3126 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3128 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3581 ( .LO ( optlc_net_3127 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3129 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3582 ( .LO ( optlc_net_3128 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3130 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3583 ( .LO ( optlc_net_3129 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3131 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3584 ( .LO ( optlc_net_3130 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3132 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3585 ( .LO ( optlc_net_3131 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3133 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3586 ( .LO ( optlc_net_3132 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3134 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3587 ( .LO ( optlc_net_3133 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3135 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3588 ( .LO ( optlc_net_3134 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3136 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3589 ( .LO ( optlc_net_3135 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3137 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3590 ( .LO ( optlc_net_3136 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3138 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3591 ( .LO ( optlc_net_3137 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3139 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3592 ( .LO ( optlc_net_3138 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3140 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3593 ( .LO ( optlc_net_3139 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3141 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3594 ( .LO ( optlc_net_3140 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3142 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3595 ( .LO ( optlc_net_3141 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3143 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3596 ( .LO ( optlc_net_3142 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3144 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3597 ( .LO ( optlc_net_3143 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3145 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3598 ( .LO ( optlc_net_3144 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3146 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3599 ( .LO ( optlc_net_3145 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3147 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3600 ( .LO ( optlc_net_3146 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3148 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3601 ( .LO ( optlc_net_3147 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3149 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3602 ( .LO ( optlc_net_3148 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3150 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3603 ( .LO ( optlc_net_3149 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3151 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3604 ( .LO ( optlc_net_3150 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3152 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3605 ( .LO ( optlc_net_3151 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3153 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3606 ( .LO ( optlc_net_3152 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3154 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3607 ( .LO ( optlc_net_3153 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3155 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3608 ( .LO ( optlc_net_3154 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3156 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3609 ( .LO ( optlc_net_3155 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3157 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3610 ( .LO ( optlc_net_3156 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3158 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3611 ( .LO ( optlc_net_3157 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3159 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3612 ( .LO ( optlc_net_3158 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3160 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3613 ( .LO ( optlc_net_3159 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3161 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3614 ( .LO ( optlc_net_3160 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3162 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3615 ( .LO ( optlc_net_3161 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3163 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3616 ( .LO ( optlc_net_3162 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3164 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3617 ( .LO ( optlc_net_3163 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3165 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3618 ( .LO ( optlc_net_3164 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3166 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3619 ( .LO ( optlc_net_3165 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3167 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3620 ( .LO ( optlc_net_3166 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3168 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3621 ( .LO ( optlc_net_3167 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3169 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3622 ( .LO ( optlc_net_3168 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3170 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3623 ( .LO ( optlc_net_3169 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3171 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3624 ( .LO ( optlc_net_3170 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3172 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3625 ( .LO ( optlc_net_3171 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3173 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3626 ( .LO ( optlc_net_3172 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3174 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3627 ( .LO ( optlc_net_3173 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3175 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3628 ( .LO ( optlc_net_3174 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3176 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3629 ( .LO ( optlc_net_3175 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3177 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3630 ( .LO ( optlc_net_3176 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3178 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3631 ( .LO ( optlc_net_3177 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3179 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3632 ( .LO ( optlc_net_3178 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3180 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3633 ( .LO ( optlc_net_3179 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3181 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3635 ( .LO ( optlc_net_3180 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3182 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3636 ( .LO ( optlc_net_3181 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3183 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3638 ( .LO ( optlc_net_3182 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3184 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3639 ( .LO ( optlc_net_3183 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3185 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3641 ( .LO ( optlc_net_3184 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3186 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3642 ( .LO ( optlc_net_3185 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3187 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3643 ( .LO ( optlc_net_3186 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3188 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3644 ( .LO ( optlc_net_3187 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3189 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3645 ( .LO ( optlc_net_3188 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3190 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3646 ( .LO ( optlc_net_3189 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3191 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3647 ( .LO ( optlc_net_3190 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3192 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3648 ( .LO ( optlc_net_3191 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3193 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3649 ( .LO ( optlc_net_3192 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3194 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3650 ( .LO ( optlc_net_3193 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3195 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3651 ( .LO ( optlc_net_3194 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3196 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3652 ( .LO ( optlc_net_3195 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3197 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3653 ( .LO ( optlc_net_3196 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3198 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3654 ( .LO ( optlc_net_3197 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3199 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3655 ( .LO ( optlc_net_3198 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3200 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3656 ( .LO ( optlc_net_3199 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3201 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3657 ( .LO ( optlc_net_3200 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3202 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3658 ( .LO ( optlc_net_3201 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3203 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3659 ( .LO ( optlc_net_3202 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3204 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3660 ( .LO ( optlc_net_3203 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3205 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3661 ( .LO ( optlc_net_3204 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3206 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3662 ( .LO ( optlc_net_3205 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3207 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3664 ( .LO ( optlc_net_3206 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3208 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3665 ( .LO ( optlc_net_3207 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3209 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3666 ( .LO ( optlc_net_3208 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3210 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3667 ( .LO ( optlc_net_3209 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3211 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3668 ( .LO ( optlc_net_3210 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3212 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3669 ( .LO ( optlc_net_3211 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3213 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3670 ( .LO ( optlc_net_3212 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3214 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3671 ( .LO ( optlc_net_3213 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3215 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3672 ( .LO ( optlc_net_3214 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3216 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3673 ( .LO ( optlc_net_3215 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3217 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3674 ( .LO ( optlc_net_3216 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3218 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3675 ( .LO ( optlc_net_3217 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3219 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3676 ( .LO ( optlc_net_3218 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3220 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3677 ( .LO ( optlc_net_3219 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3221 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3678 ( .LO ( optlc_net_3220 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3222 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3679 ( .LO ( optlc_net_3221 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3223 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3680 ( .LO ( optlc_net_3222 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3224 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3681 ( .LO ( optlc_net_3223 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3225 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3682 ( .LO ( optlc_net_3224 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3226 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3683 ( .LO ( optlc_net_3225 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3227 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3684 ( .LO ( optlc_net_3226 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3228 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3685 ( .LO ( optlc_net_3227 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3229 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3686 ( .LO ( optlc_net_3228 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3230 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3687 ( .LO ( optlc_net_3229 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3231 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3688 ( .LO ( optlc_net_3230 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3232 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3689 ( .LO ( optlc_net_3231 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3233 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3690 ( .LO ( optlc_net_3232 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3234 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3691 ( .LO ( optlc_net_3233 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3235 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3692 ( .LO ( optlc_net_3234 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3236 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3693 ( .LO ( optlc_net_3235 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3237 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3694 ( .LO ( optlc_net_3236 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3238 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3695 ( .LO ( optlc_net_3237 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3239 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3696 ( .LO ( optlc_net_3238 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3240 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3697 ( .LO ( optlc_net_3239 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3241 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3698 ( .LO ( optlc_net_3240 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3242 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3699 ( .LO ( optlc_net_3241 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3243 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3700 ( .LO ( optlc_net_3242 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3244 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3701 ( .LO ( optlc_net_3243 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3245 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3702 ( .LO ( optlc_net_3244 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3246 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3703 ( .LO ( optlc_net_3245 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3247 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3704 ( .LO ( optlc_net_3246 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3248 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3705 ( .LO ( optlc_net_3247 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3249 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3706 ( .LO ( optlc_net_3248 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3250 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3707 ( .LO ( optlc_net_3249 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3251 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3708 ( .LO ( optlc_net_3250 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3252 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3709 ( .LO ( optlc_net_3251 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3253 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3710 ( .LO ( optlc_net_3252 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3254 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3711 ( .LO ( optlc_net_3253 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3255 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3712 ( .LO ( optlc_net_3254 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3256 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3713 ( .LO ( optlc_net_3255 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3257 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3714 ( .LO ( optlc_net_3256 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3258 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3715 ( .LO ( optlc_net_3257 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3259 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3716 ( .LO ( optlc_net_3258 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3260 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3717 ( .LO ( optlc_net_3259 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3261 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3719 ( .LO ( optlc_net_3260 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3262 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3721 ( .LO ( optlc_net_3261 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3263 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3722 ( .LO ( optlc_net_3262 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3264 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3723 ( .LO ( optlc_net_3263 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3265 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3724 ( .LO ( optlc_net_3264 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3266 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3725 ( .LO ( optlc_net_3265 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3267 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3726 ( .LO ( optlc_net_3266 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3268 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3727 ( .LO ( optlc_net_3267 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3269 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3728 ( .LO ( optlc_net_3268 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3270 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3729 ( .LO ( optlc_net_3269 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3271 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3730 ( .LO ( optlc_net_3270 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3272 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3731 ( .LO ( optlc_net_3271 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3273 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3732 ( .LO ( optlc_net_3272 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3274 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3733 ( .LO ( optlc_net_3273 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3275 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3734 ( .LO ( optlc_net_3274 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3276 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3735 ( .LO ( optlc_net_3275 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3277 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3736 ( .LO ( optlc_net_3276 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3278 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3737 ( .LO ( optlc_net_3277 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3279 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3738 ( .LO ( optlc_net_3278 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3280 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3739 ( .LO ( optlc_net_3279 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3281 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3740 ( .LO ( optlc_net_3280 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3282 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3741 ( .LO ( optlc_net_3281 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3283 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3742 ( .LO ( optlc_net_3282 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3284 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3743 ( .LO ( optlc_net_3283 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3285 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3744 ( .LO ( optlc_net_3284 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3286 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3745 ( .LO ( optlc_net_3285 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3287 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3746 ( .LO ( optlc_net_3286 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3288 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3747 ( .LO ( optlc_net_3287 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3289 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3748 ( .LO ( optlc_net_3288 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3290 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3749 ( .LO ( optlc_net_3289 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3291 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3750 ( .LO ( optlc_net_3290 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3292 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3751 ( .LO ( optlc_net_3291 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3293 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3752 ( .LO ( optlc_net_3292 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3294 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3753 ( .LO ( optlc_net_3293 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3295 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3754 ( .LO ( optlc_net_3294 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3296 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3755 ( .LO ( optlc_net_3295 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3297 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3756 ( .LO ( optlc_net_3296 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3298 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3757 ( .LO ( optlc_net_3297 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3299 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3758 ( .LO ( optlc_net_3298 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3300 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3759 ( .LO ( optlc_net_3299 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3301 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3760 ( .LO ( optlc_net_3300 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3302 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3761 ( .LO ( optlc_net_3301 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3303 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3762 ( .LO ( optlc_net_3302 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3304 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3763 ( .LO ( optlc_net_3303 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3305 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3764 ( .LO ( optlc_net_3304 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3306 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3765 ( .LO ( optlc_net_3305 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3307 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3766 ( .LO ( optlc_net_3306 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3308 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3767 ( .LO ( optlc_net_3307 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3309 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3768 ( .LO ( optlc_net_3308 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3310 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3769 ( .LO ( optlc_net_3309 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3311 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3770 ( .LO ( optlc_net_3310 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3312 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3771 ( .LO ( optlc_net_3311 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3313 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3772 ( .LO ( optlc_net_3312 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3314 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3773 ( .LO ( optlc_net_3313 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3315 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3774 ( .LO ( optlc_net_3314 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3316 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3775 ( .LO ( optlc_net_3315 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3317 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3776 ( .LO ( optlc_net_3316 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3318 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3777 ( .LO ( optlc_net_3317 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3319 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3778 ( .LO ( optlc_net_3318 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3320 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3779 ( .LO ( optlc_net_3319 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3321 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3780 ( .LO ( optlc_net_3320 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3322 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3781 ( .LO ( optlc_net_3321 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3323 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3782 ( .LO ( optlc_net_3322 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3324 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3783 ( .LO ( optlc_net_3323 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3325 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3784 ( .LO ( optlc_net_3324 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3326 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3785 ( .LO ( optlc_net_3325 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3327 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3786 ( .LO ( optlc_net_3326 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3328 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3787 ( .LO ( optlc_net_3327 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3329 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3788 ( .LO ( optlc_net_3328 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3330 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3789 ( .LO ( optlc_net_3329 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3331 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3790 ( .LO ( optlc_net_3330 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3332 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3791 ( .LO ( optlc_net_3331 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3333 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3792 ( .LO ( optlc_net_3332 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3334 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3793 ( .LO ( optlc_net_3333 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3335 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3794 ( .LO ( optlc_net_3334 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3336 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3795 ( .LO ( optlc_net_3335 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3337 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3796 ( .LO ( optlc_net_3336 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3338 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3797 ( .LO ( optlc_net_3337 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3339 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3798 ( .LO ( optlc_net_3338 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3340 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3799 ( .LO ( optlc_net_3339 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3341 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3800 ( .LO ( optlc_net_3340 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3342 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3801 ( .LO ( optlc_net_3341 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3343 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3802 ( .LO ( optlc_net_3342 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3344 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3803 ( .LO ( optlc_net_3343 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3345 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3804 ( .LO ( optlc_net_3344 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3346 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3805 ( .LO ( optlc_net_3345 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3347 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3806 ( .LO ( optlc_net_3346 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3348 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3807 ( .LO ( optlc_net_3347 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3349 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3808 ( .LO ( optlc_net_3348 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3350 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3809 ( .LO ( optlc_net_3349 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3351 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3810 ( .LO ( optlc_net_3350 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3352 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3811 ( .LO ( optlc_net_3351 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3353 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3812 ( .LO ( optlc_net_3352 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3354 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3813 ( .LO ( optlc_net_3353 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3355 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3814 ( .LO ( optlc_net_3354 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3356 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3815 ( .LO ( optlc_net_3355 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3357 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3816 ( .LO ( optlc_net_3356 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3358 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3817 ( .LO ( optlc_net_3357 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3359 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3818 ( .LO ( optlc_net_3358 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3360 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3819 ( .LO ( optlc_net_3359 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3361 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3820 ( .LO ( optlc_net_3360 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3362 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3821 ( .LO ( optlc_net_3361 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3363 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3822 ( .LO ( optlc_net_3362 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3364 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3823 ( .LO ( optlc_net_3363 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3365 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3824 ( .LO ( optlc_net_3364 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3366 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3825 ( .LO ( optlc_net_3365 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3367 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3826 ( .LO ( optlc_net_3366 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3368 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3827 ( .LO ( optlc_net_3367 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3369 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3828 ( .LO ( optlc_net_3368 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3370 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3829 ( .LO ( optlc_net_3369 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3371 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3830 ( .LO ( optlc_net_3370 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3372 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3831 ( .LO ( optlc_net_3371 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3373 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3832 ( .LO ( optlc_net_3372 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3374 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3833 ( .LO ( optlc_net_3373 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3375 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3834 ( .LO ( optlc_net_3374 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3376 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3835 ( .LO ( optlc_net_3375 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3377 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3836 ( .LO ( optlc_net_3376 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3378 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3837 ( .LO ( optlc_net_3377 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3379 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3838 ( .LO ( optlc_net_3378 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3380 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3839 ( .LO ( optlc_net_3379 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3381 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3840 ( .LO ( optlc_net_3380 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3382 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3841 ( .LO ( optlc_net_3381 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3383 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3842 ( .LO ( optlc_net_3382 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3384 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3843 ( .LO ( optlc_net_3383 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3385 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3844 ( .LO ( optlc_net_3384 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3386 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3845 ( .LO ( optlc_net_3385 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3387 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3846 ( .LO ( optlc_net_3386 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3388 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3847 ( .LO ( optlc_net_3387 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3389 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3848 ( .LO ( optlc_net_3388 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3390 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3849 ( .LO ( optlc_net_3389 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3391 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3850 ( .LO ( optlc_net_3390 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3392 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3851 ( .LO ( optlc_net_3391 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3393 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3852 ( .LO ( optlc_net_3392 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3394 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3853 ( .LO ( optlc_net_3393 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3395 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3854 ( .LO ( optlc_net_3394 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3396 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3855 ( .LO ( optlc_net_3395 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3397 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3856 ( .LO ( optlc_net_3396 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3398 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3857 ( .LO ( optlc_net_3397 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3399 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3858 ( .LO ( optlc_net_3398 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3400 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3859 ( .LO ( optlc_net_3399 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3401 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3860 ( .LO ( optlc_net_3400 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3402 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3861 ( .LO ( optlc_net_3401 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3403 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3862 ( .LO ( optlc_net_3402 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3404 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3863 ( .LO ( optlc_net_3403 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3405 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3864 ( .LO ( optlc_net_3404 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3406 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3865 ( .LO ( optlc_net_3405 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3407 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3866 ( .LO ( optlc_net_3406 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3408 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3867 ( .LO ( optlc_net_3407 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3409 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3868 ( .LO ( optlc_net_3408 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3410 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3869 ( .LO ( optlc_net_3409 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3411 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3870 ( .LO ( optlc_net_3410 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3412 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3871 ( .LO ( optlc_net_3411 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3413 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3872 ( .LO ( optlc_net_3412 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3414 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3873 ( .LO ( optlc_net_3413 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3415 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3874 ( .LO ( optlc_net_3414 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3416 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3875 ( .LO ( optlc_net_3415 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3417 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3876 ( .LO ( optlc_net_3416 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3418 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3877 ( .LO ( optlc_net_3417 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3419 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3878 ( .LO ( optlc_net_3418 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3420 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3879 ( .LO ( optlc_net_3419 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3421 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3880 ( .LO ( optlc_net_3420 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3422 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3881 ( .LO ( optlc_net_3421 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3423 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3882 ( .LO ( optlc_net_3422 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3424 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3883 ( .LO ( optlc_net_3423 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3425 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3884 ( .LO ( optlc_net_3424 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3426 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3885 ( .LO ( optlc_net_3425 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3427 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3886 ( .LO ( optlc_net_3426 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3428 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3887 ( .LO ( optlc_net_3427 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3429 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3888 ( .LO ( optlc_net_3428 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3430 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3889 ( .LO ( optlc_net_3429 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3431 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3890 ( .LO ( optlc_net_3430 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3432 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3891 ( .LO ( optlc_net_3431 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3433 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3892 ( .LO ( optlc_net_3432 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3434 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3893 ( .LO ( optlc_net_3433 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3435 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3894 ( .LO ( optlc_net_3434 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3436 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3895 ( .LO ( optlc_net_3435 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3437 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3896 ( .LO ( optlc_net_3436 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3438 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3897 ( .LO ( optlc_net_3437 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3439 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3898 ( .LO ( optlc_net_3438 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3440 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3899 ( .LO ( optlc_net_3439 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3441 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3900 ( .LO ( optlc_net_3440 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3442 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3901 ( .LO ( optlc_net_3441 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3443 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3902 ( .LO ( optlc_net_3442 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3444 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3903 ( .LO ( optlc_net_3443 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3445 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3904 ( .LO ( optlc_net_3444 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3446 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3905 ( .LO ( optlc_net_3445 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3447 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3906 ( .LO ( optlc_net_3446 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3448 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3907 ( .LO ( optlc_net_3447 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3449 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3908 ( .LO ( optlc_net_3448 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3450 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3909 ( .LO ( optlc_net_3449 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3451 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3910 ( .LO ( optlc_net_3450 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3452 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3911 ( .LO ( optlc_net_3451 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3453 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3912 ( .LO ( optlc_net_3452 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3454 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3913 ( .LO ( optlc_net_3453 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3455 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3914 ( .LO ( optlc_net_3454 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3456 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3915 ( .LO ( optlc_net_3455 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3457 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3916 ( .LO ( optlc_net_3456 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3458 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3917 ( .LO ( optlc_net_3457 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3459 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3918 ( .LO ( optlc_net_3458 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3460 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3919 ( .LO ( optlc_net_3459 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3461 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3920 ( .LO ( optlc_net_3460 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3462 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3921 ( .LO ( optlc_net_3461 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3463 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3922 ( .LO ( optlc_net_3462 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3464 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3923 ( .LO ( optlc_net_3463 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3465 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3924 ( .LO ( optlc_net_3464 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3466 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3925 ( .LO ( optlc_net_3465 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3467 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3926 ( .LO ( optlc_net_3466 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3468 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3927 ( .LO ( optlc_net_3467 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3469 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3928 ( .LO ( optlc_net_3468 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3470 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3929 ( .LO ( optlc_net_3469 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3471 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3930 ( .LO ( optlc_net_3470 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3472 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3931 ( .LO ( optlc_net_3471 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3473 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3932 ( .LO ( optlc_net_3472 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3474 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3933 ( .LO ( optlc_net_3473 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3475 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3934 ( .LO ( optlc_net_3474 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3476 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3935 ( .LO ( optlc_net_3475 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3477 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3936 ( .LO ( optlc_net_3476 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3478 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3937 ( .LO ( optlc_net_3477 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3479 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3938 ( .LO ( optlc_net_3478 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3480 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3939 ( .LO ( optlc_net_3479 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3481 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3940 ( .LO ( optlc_net_3480 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3482 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3941 ( .LO ( optlc_net_3481 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3483 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3942 ( .LO ( optlc_net_3482 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3484 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3943 ( .LO ( optlc_net_3483 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3485 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3944 ( .LO ( optlc_net_3484 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3486 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3945 ( .LO ( optlc_net_3485 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3487 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3946 ( .LO ( optlc_net_3486 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3488 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3947 ( .LO ( optlc_net_3487 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3489 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3948 ( .LO ( optlc_net_3488 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3490 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3949 ( .LO ( optlc_net_3489 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3491 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3950 ( .LO ( optlc_net_3490 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3492 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3951 ( .LO ( optlc_net_3491 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3493 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3952 ( .LO ( optlc_net_3492 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3494 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3953 ( .LO ( optlc_net_3493 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3495 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3954 ( .LO ( optlc_net_3494 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3496 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3955 ( .LO ( optlc_net_3495 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3497 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3956 ( .LO ( optlc_net_3496 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3498 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3957 ( .LO ( optlc_net_3497 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3499 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3958 ( .LO ( optlc_net_3498 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3500 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3959 ( .LO ( optlc_net_3499 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3501 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3960 ( .LO ( optlc_net_3500 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3502 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3961 ( .LO ( optlc_net_3501 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3503 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3962 ( .LO ( optlc_net_3502 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3504 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3963 ( .LO ( optlc_net_3503 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3505 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3964 ( .LO ( optlc_net_3504 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3506 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3965 ( .LO ( optlc_net_3505 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3507 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3966 ( .LO ( optlc_net_3506 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3508 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3967 ( .LO ( optlc_net_3507 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3509 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3968 ( .LO ( optlc_net_3508 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3510 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3969 ( .LO ( optlc_net_3509 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3511 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3970 ( .LO ( optlc_net_3510 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3512 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3971 ( .LO ( optlc_net_3511 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3513 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3972 ( .LO ( optlc_net_3512 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3514 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3973 ( .LO ( optlc_net_3513 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3515 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3974 ( .LO ( optlc_net_3514 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3516 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3975 ( .LO ( optlc_net_3515 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3517 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3976 ( .LO ( optlc_net_3516 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3518 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3977 ( .LO ( optlc_net_3517 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3519 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3978 ( .LO ( optlc_net_3518 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3520 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3979 ( .LO ( optlc_net_3519 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3521 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3980 ( .LO ( optlc_net_3520 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3522 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3981 ( .LO ( optlc_net_3521 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3523 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3982 ( .LO ( optlc_net_3522 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3524 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3983 ( .LO ( optlc_net_3523 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3525 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3984 ( .LO ( optlc_net_3524 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3526 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3985 ( .LO ( optlc_net_3525 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3527 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3986 ( .LO ( optlc_net_3526 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3528 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3987 ( .LO ( optlc_net_3527 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3529 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3988 ( .LO ( optlc_net_3528 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3530 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_3989 ( .LO ( optlc_net_3529 ) , 
    .HI ( SYNOPSYS_UNCONNECTED_3531 ) ) ;
endmodule


