VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER fieldpoly
  TYPE MASTERSLICE ;
END fieldpoly

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER diff
  TYPE MASTERSLICE ;
END diff

LAYER licon1
  TYPE MASTERSLICE ;
END licon1

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_1__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 141.68 BY 130.56 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 2.23 27.2 2.37 28.56 ;
    END
  END prog_clk[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.43 129.2 80.57 130.56 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 129.2 57.57 130.56 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.27 129.2 82.41 130.56 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.99 129.2 74.13 130.56 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 129.2 52.05 130.56 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.19 129.2 60.33 130.56 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.91 129.2 75.05 130.56 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.63 129.2 66.77 130.56 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.15 129.2 72.29 130.56 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.55 129.2 67.69 130.56 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.07 129.2 73.21 130.56 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.83 129.2 75.97 130.56 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 129.2 52.97 130.56 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.41 129.2 63.55 130.56 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.67 129.2 54.81 130.56 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.75 129.2 53.89 130.56 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.39 129.2 69.53 130.56 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.35 129.2 81.49 130.56 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.57 129.2 84.71 130.56 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.27 129.2 59.41 130.56 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.67 129.2 31.81 130.56 ;
    END
  END top_left_grid_pin_34_[0]
  PIN top_left_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.59 129.2 32.73 130.56 ;
    END
  END top_left_grid_pin_35_[0]
  PIN top_left_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 127.01 29.9 127.31 ;
    END
  END top_left_grid_pin_36_[0]
  PIN top_left_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.75 129.2 30.89 130.56 ;
    END
  END top_left_grid_pin_37_[0]
  PIN top_left_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 124.97 29.9 125.27 ;
    END
  END top_left_grid_pin_38_[0]
  PIN top_left_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 123.61 29.9 123.91 ;
    END
  END top_left_grid_pin_39_[0]
  PIN top_left_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 122.25 29.9 122.55 ;
    END
  END top_left_grid_pin_40_[0]
  PIN top_left_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 117.49 29.9 117.79 ;
    END
  END top_left_grid_pin_41_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 48.81 141.68 49.11 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 99.13 141.68 99.43 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 55.61 141.68 55.91 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 37.93 141.68 38.23 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 93.69 141.68 93.99 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 95.05 141.68 95.35 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 77.37 141.68 77.67 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 69.21 141.68 69.51 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 44.73 141.68 45.03 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 50.85 141.68 51.15 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 36.57 141.68 36.87 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 43.37 141.68 43.67 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 96.41 141.68 96.71 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 32.49 141.68 32.79 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 90.97 141.68 91.27 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 56.97 141.68 57.27 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 39.29 141.68 39.59 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 33.85 141.68 34.15 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 65.13 141.68 65.43 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 31.13 141.68 31.43 ;
    END
  END chanx_right_in[19]
  PIN right_top_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.39 102 138.53 103.36 ;
    END
  END right_top_grid_pin_42_[0]
  PIN right_top_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 126.33 113.16 126.63 ;
    END
  END right_top_grid_pin_43_[0]
  PIN right_top_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.31 102 139.45 103.36 ;
    END
  END right_top_grid_pin_44_[0]
  PIN right_top_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.47 102 137.61 103.36 ;
    END
  END right_top_grid_pin_45_[0]
  PIN right_top_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 118.85 113.16 119.15 ;
    END
  END right_top_grid_pin_46_[0]
  PIN right_top_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 117.49 113.16 117.79 ;
    END
  END right_top_grid_pin_47_[0]
  PIN right_top_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.63 102 135.77 103.36 ;
    END
  END right_top_grid_pin_48_[0]
  PIN right_top_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.55 102 136.69 103.36 ;
    END
  END right_top_grid_pin_49_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.27 0 82.41 1.36 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.09 0 67.23 1.36 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.35 0 81.49 1.36 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.25 0 88.39 1.36 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.25 0 65.39 1.36 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.83 0 75.97 1.36 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.23 0 94.37 1.36 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.33 0 87.47 1.36 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.67 0 77.81 1.36 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.11 0 84.25 1.36 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.49 0 62.63 1.36 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.41 0 86.55 1.36 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.51 0 79.65 1.36 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.01 0 68.15 1.36 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.17 0 66.31 1.36 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.29 0 53.43 1.36 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.75 0 76.89 1.36 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.85 0 69.99 1.36 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 0 57.57 1.36 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.59 0 78.73 1.36 ;
    END
  END chany_bottom_in[19]
  PIN bottom_left_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 10.05 29.9 10.35 ;
    END
  END bottom_left_grid_pin_34_[0]
  PIN bottom_left_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 8.01 29.9 8.31 ;
    END
  END bottom_left_grid_pin_35_[0]
  PIN bottom_left_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 6.65 29.9 6.95 ;
    END
  END bottom_left_grid_pin_36_[0]
  PIN bottom_left_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 3.25 29.9 3.55 ;
    END
  END bottom_left_grid_pin_37_[0]
  PIN bottom_left_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 4.61 29.9 4.91 ;
    END
  END bottom_left_grid_pin_38_[0]
  PIN bottom_left_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 11.41 29.9 11.71 ;
    END
  END bottom_left_grid_pin_39_[0]
  PIN bottom_left_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 12.77 29.9 13.07 ;
    END
  END bottom_left_grid_pin_40_[0]
  PIN bottom_left_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 14.13 29.9 14.43 ;
    END
  END bottom_left_grid_pin_41_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 76.01 1.38 76.31 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.93 1.38 38.23 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 35.21 1.38 35.51 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.29 1.38 39.59 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 85.53 1.38 85.83 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 86.89 1.38 87.19 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.85 1.38 34.15 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.01 1.38 42.31 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.37 1.38 43.67 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 71.93 1.38 72.23 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.01 1.38 59.31 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.57 1.38 36.87 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 97.77 1.38 98.07 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 93.69 1.38 93.99 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 92.33 1.38 92.63 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 77.37 1.38 77.67 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 51.53 1.38 51.83 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 55.61 1.38 55.91 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 67.85 1.38 68.15 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 46.09 1.38 46.39 ;
    END
  END chanx_left_in[19]
  PIN left_top_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.29 102 7.43 103.36 ;
    END
  END left_top_grid_pin_42_[0]
  PIN left_top_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 118.85 29.9 119.15 ;
    END
  END left_top_grid_pin_43_[0]
  PIN left_top_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.07 102 4.21 103.36 ;
    END
  END left_top_grid_pin_44_[0]
  PIN left_top_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.99 102 5.13 103.36 ;
    END
  END left_top_grid_pin_45_[0]
  PIN left_top_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.23 102 2.37 103.36 ;
    END
  END left_top_grid_pin_46_[0]
  PIN left_top_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.15 102 3.29 103.36 ;
    END
  END left_top_grid_pin_47_[0]
  PIN left_top_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.43 102 11.57 103.36 ;
    END
  END left_top_grid_pin_48_[0]
  PIN left_top_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.51 102 10.65 103.36 ;
    END
  END left_top_grid_pin_49_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 88.25 141.68 88.55 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.75 129.2 76.89 130.56 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.11 129.2 61.25 130.56 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.67 129.2 77.81 130.56 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.23 129.2 71.37 130.56 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.83 129.2 98.97 130.56 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.65 129.2 83.79 130.56 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.31 129.2 70.45 130.56 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 129.2 50.21 130.56 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.47 129.2 68.61 130.56 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.35 129.2 58.49 130.56 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.53 129.2 96.67 130.56 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.77 129.2 93.91 130.56 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.51 129.2 79.65 130.56 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.33 129.2 64.47 130.56 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.45 129.2 97.59 130.56 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 129.2 51.13 130.56 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.87 129.2 87.01 130.56 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.03 129.2 62.17 130.56 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.61 129.2 95.75 130.56 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.59 129.2 78.73 130.56 ;
    END
  END chany_top_out[19]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 84.17 141.68 84.47 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 82.81 141.68 83.11 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 62.41 141.68 62.71 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 73.97 141.68 74.27 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 80.09 141.68 80.39 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 71.93 141.68 72.23 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 58.33 141.68 58.63 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 35.21 141.68 35.51 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 46.09 141.68 46.39 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 63.77 141.68 64.07 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 61.05 141.68 61.35 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 78.73 141.68 79.03 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 42.01 141.68 42.31 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 85.53 141.68 85.83 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 47.45 141.68 47.75 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 67.85 141.68 68.15 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 40.65 141.68 40.95 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 66.49 141.68 66.79 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 52.21 141.68 52.51 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 89.61 141.68 89.91 ;
    END
  END chanx_right_out[19]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.19 0 83.33 1.36 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.73 0 59.87 1.36 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.37 0 52.51 1.36 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.93 0 69.07 1.36 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.53 0 96.67 1.36 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.69 0 71.83 1.36 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.91 0 75.05 1.36 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.65 0 60.79 1.36 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.41 0 63.55 1.36 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.21 0 54.35 1.36 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.31 0 93.45 1.36 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.99 0 74.13 1.36 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.43 0 80.57 1.36 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.57 0 61.71 1.36 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.45 0 97.59 1.36 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.13 0 55.27 1.36 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.33 0 64.47 1.36 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.81 0 58.95 1.36 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.07 0 73.21 1.36 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.77 0 70.91 1.36 ;
    END
  END chany_bottom_out[19]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 61.05 1.38 61.35 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 81.45 1.38 81.75 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 82.81 1.38 83.11 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 74.65 1.38 74.95 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 80.09 1.38 80.39 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 47.45 1.38 47.75 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.17 1.38 50.47 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 65.81 1.38 66.11 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.81 1.38 49.11 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.21 1.38 69.51 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.89 1.38 53.19 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 96.41 1.38 96.71 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.73 1.38 45.03 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 99.13 1.38 99.43 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 54.25 1.38 54.55 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 40.65 1.38 40.95 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.81 1.38 32.11 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 88.25 1.38 88.55 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 70.57 1.38 70.87 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 90.97 1.38 91.27 ;
    END
  END chanx_left_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 64.45 1.38 64.75 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 28.52 2.48 29 2.96 ;
        RECT 112.68 2.48 113.16 2.96 ;
        RECT 28.52 7.92 29 8.4 ;
        RECT 112.68 7.92 113.16 8.4 ;
        RECT 28.52 13.36 29 13.84 ;
        RECT 112.68 13.36 113.16 13.84 ;
        RECT 28.52 18.8 29 19.28 ;
        RECT 112.68 18.8 113.16 19.28 ;
        RECT 28.52 24.24 29 24.72 ;
        RECT 112.68 24.24 113.16 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 141.2 29.68 141.68 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 141.2 35.12 141.68 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 141.2 40.56 141.68 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 141.2 46 141.68 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 141.2 51.44 141.68 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 141.2 56.88 141.68 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 141.2 62.32 141.68 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 141.2 67.76 141.68 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 141.2 73.2 141.68 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 141.2 78.64 141.68 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 141.2 84.08 141.68 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 141.2 89.52 141.68 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 141.2 94.96 141.68 95.44 ;
        RECT 0 100.4 0.48 100.88 ;
        RECT 141.2 100.4 141.68 100.88 ;
        RECT 28.52 105.84 29 106.32 ;
        RECT 112.68 105.84 113.16 106.32 ;
        RECT 28.52 111.28 29 111.76 ;
        RECT 112.68 111.28 113.16 111.76 ;
        RECT 28.52 116.72 29 117.2 ;
        RECT 112.68 116.72 113.16 117.2 ;
        RECT 28.52 122.16 29 122.64 ;
        RECT 112.68 122.16 113.16 122.64 ;
        RECT 28.52 127.6 29 128.08 ;
        RECT 112.68 127.6 113.16 128.08 ;
      LAYER met5 ;
        RECT 0 43.28 3.2 46.48 ;
        RECT 138.48 43.28 141.68 46.48 ;
        RECT 0 84.08 3.2 87.28 ;
        RECT 138.48 84.08 141.68 87.28 ;
        RECT 28.52 122.84 31.72 126.04 ;
        RECT 109.96 122.84 113.16 126.04 ;
      LAYER met4 ;
        RECT 41.1 0 41.7 0.6 ;
        RECT 70.54 0 71.14 0.6 ;
        RECT 99.98 0 100.58 0.6 ;
        RECT 134.94 27.2 135.54 27.8 ;
        RECT 134.94 102.76 135.54 103.36 ;
        RECT 41.1 129.96 41.7 130.56 ;
        RECT 70.54 129.96 71.14 130.56 ;
        RECT 99.98 129.96 100.58 130.56 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 28.52 0 113.16 0.24 ;
        RECT 28.52 5.2 29 5.68 ;
        RECT 112.68 5.2 113.16 5.68 ;
        RECT 28.52 10.64 29 11.12 ;
        RECT 112.68 10.64 113.16 11.12 ;
        RECT 28.52 16.08 29 16.56 ;
        RECT 112.68 16.08 113.16 16.56 ;
        RECT 28.52 21.52 29 22 ;
        RECT 112.68 21.52 113.16 22 ;
        RECT 0 26.96 141.68 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 141.2 32.4 141.68 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 141.2 37.84 141.68 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 141.2 43.28 141.68 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 141.2 48.72 141.68 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 141.2 54.16 141.68 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 141.2 59.6 141.68 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 141.2 65.04 141.68 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 141.2 70.48 141.68 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 141.2 75.92 141.68 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 141.2 81.36 141.68 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 141.2 86.8 141.68 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 141.2 92.24 141.68 92.72 ;
        RECT 0 97.68 0.48 98.16 ;
        RECT 141.2 97.68 141.68 98.16 ;
        RECT 0 103.12 141.68 103.6 ;
        RECT 28.52 108.56 29 109.04 ;
        RECT 112.68 108.56 113.16 109.04 ;
        RECT 28.52 114 29 114.48 ;
        RECT 112.68 114 113.16 114.48 ;
        RECT 28.52 119.44 29 119.92 ;
        RECT 112.68 119.44 113.16 119.92 ;
        RECT 28.52 124.88 29 125.36 ;
        RECT 112.68 124.88 113.16 125.36 ;
        RECT 28.52 130.32 113.16 130.56 ;
      LAYER met5 ;
        RECT 28.52 4.52 31.72 7.72 ;
        RECT 109.96 4.52 113.16 7.72 ;
        RECT 0 63.68 3.2 66.88 ;
        RECT 138.48 63.68 141.68 66.88 ;
      LAYER met4 ;
        RECT 55.82 0 56.42 0.6 ;
        RECT 85.26 0 85.86 0.6 ;
        RECT 6.14 27.2 6.74 27.8 ;
        RECT 6.14 102.76 6.74 103.36 ;
        RECT 55.82 129.96 56.42 130.56 ;
        RECT 85.26 129.96 85.86 130.56 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 28.52 130.475 113.16 130.645 ;
      RECT 109.48 127.755 113.16 127.925 ;
      RECT 28.52 127.755 32.2 127.925 ;
      RECT 112.24 125.035 113.16 125.205 ;
      RECT 28.52 125.035 32.2 125.205 ;
      RECT 112.24 122.315 113.16 122.485 ;
      RECT 28.52 122.315 32.2 122.485 ;
      RECT 112.24 119.595 113.16 119.765 ;
      RECT 28.52 119.595 32.2 119.765 ;
      RECT 112.24 116.875 113.16 117.045 ;
      RECT 28.52 116.875 32.2 117.045 ;
      RECT 112.7 114.155 113.16 114.325 ;
      RECT 28.52 114.155 30.36 114.325 ;
      RECT 112.24 111.435 113.16 111.605 ;
      RECT 28.52 111.435 32.2 111.605 ;
      RECT 112.24 108.715 113.16 108.885 ;
      RECT 28.52 108.715 32.2 108.885 ;
      RECT 112.24 105.995 113.16 106.165 ;
      RECT 28.52 105.995 32.2 106.165 ;
      RECT 110.4 103.275 141.68 103.445 ;
      RECT 0 103.275 30.36 103.445 ;
      RECT 139.84 100.555 141.68 100.725 ;
      RECT 0 100.555 3.68 100.725 ;
      RECT 141.22 97.835 141.68 98.005 ;
      RECT 0 97.835 1.84 98.005 ;
      RECT 140.76 95.115 141.68 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 140.76 92.395 141.68 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 140.76 89.675 141.68 89.845 ;
      RECT 0 89.675 1.84 89.845 ;
      RECT 140.76 86.955 141.68 87.125 ;
      RECT 0 86.955 1.84 87.125 ;
      RECT 140.76 84.235 141.68 84.405 ;
      RECT 0 84.235 1.84 84.405 ;
      RECT 140.76 81.515 141.68 81.685 ;
      RECT 0 81.515 1.84 81.685 ;
      RECT 140.76 78.795 141.68 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 140.76 76.075 141.68 76.245 ;
      RECT 0 76.075 1.84 76.245 ;
      RECT 140.76 73.355 141.68 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 140.76 70.635 141.68 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 140.76 67.915 141.68 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 140.76 65.195 141.68 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 140.76 62.475 141.68 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 140.76 59.755 141.68 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 140.76 57.035 141.68 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 140.76 54.315 141.68 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 140.76 51.595 141.68 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 140.76 48.875 141.68 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 140.76 46.155 141.68 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 140.76 43.435 141.68 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 141.22 40.715 141.68 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 140.76 37.995 141.68 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 140.76 35.275 141.68 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 140.76 32.555 141.68 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 141.22 29.835 141.68 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 110.86 27.115 141.68 27.285 ;
      RECT 0 27.115 32.2 27.285 ;
      RECT 112.7 24.395 113.16 24.565 ;
      RECT 28.52 24.395 32.2 24.565 ;
      RECT 112.24 21.675 113.16 21.845 ;
      RECT 28.52 21.675 32.2 21.845 ;
      RECT 112.24 18.955 113.16 19.125 ;
      RECT 28.52 18.955 32.2 19.125 ;
      RECT 109.48 16.235 113.16 16.405 ;
      RECT 28.52 16.235 32.2 16.405 ;
      RECT 109.48 13.515 113.16 13.685 ;
      RECT 28.52 13.515 32.2 13.685 ;
      RECT 109.48 10.795 113.16 10.965 ;
      RECT 28.52 10.795 32.2 10.965 ;
      RECT 109.48 8.075 113.16 8.245 ;
      RECT 28.52 8.075 32.2 8.245 ;
      RECT 112.24 5.355 113.16 5.525 ;
      RECT 28.52 5.355 32.2 5.525 ;
      RECT 109.48 2.635 113.16 2.805 ;
      RECT 28.52 2.635 32.2 2.805 ;
      RECT 28.52 -0.085 113.16 0.085 ;
    LAYER met2 ;
      RECT 85.42 130.375 85.7 130.745 ;
      RECT 55.98 130.375 56.26 130.745 ;
      RECT 84.97 128.7 85.23 129.02 ;
      RECT 75.31 128.7 75.57 129.02 ;
      RECT 6.3 103.175 6.58 103.545 ;
      RECT 6.3 27.015 6.58 27.385 ;
      RECT 63.81 1.54 64.07 1.86 ;
      RECT 69.3 1.57 69.62 1.83 ;
      RECT 85.42 -0.185 85.7 0.185 ;
      RECT 55.98 -0.185 56.26 0.185 ;
      POLYGON 112.88 130.28 112.88 103.08 135.35 103.08 135.35 101.72 136.05 101.72 136.05 103.08 136.27 103.08 136.27 101.72 136.97 101.72 136.97 103.08 137.19 103.08 137.19 101.72 137.89 101.72 137.89 103.08 138.11 103.08 138.11 101.72 138.81 101.72 138.81 103.08 139.03 103.08 139.03 101.72 139.73 101.72 139.73 103.08 141.4 103.08 141.4 27.48 112.88 27.48 112.88 0.28 97.87 0.28 97.87 1.64 97.17 1.64 97.17 0.28 96.95 0.28 96.95 1.64 96.25 1.64 96.25 0.28 94.65 0.28 94.65 1.64 93.95 1.64 93.95 0.28 93.73 0.28 93.73 1.64 93.03 1.64 93.03 0.28 88.67 0.28 88.67 1.64 87.97 1.64 87.97 0.28 87.75 0.28 87.75 1.64 87.05 1.64 87.05 0.28 86.83 0.28 86.83 1.64 86.13 1.64 86.13 0.28 84.53 0.28 84.53 1.64 83.83 1.64 83.83 0.28 83.61 0.28 83.61 1.64 82.91 1.64 82.91 0.28 82.69 0.28 82.69 1.64 81.99 1.64 81.99 0.28 81.77 0.28 81.77 1.64 81.07 1.64 81.07 0.28 80.85 0.28 80.85 1.64 80.15 1.64 80.15 0.28 79.93 0.28 79.93 1.64 79.23 1.64 79.23 0.28 79.01 0.28 79.01 1.64 78.31 1.64 78.31 0.28 78.09 0.28 78.09 1.64 77.39 1.64 77.39 0.28 77.17 0.28 77.17 1.64 76.47 1.64 76.47 0.28 76.25 0.28 76.25 1.64 75.55 1.64 75.55 0.28 75.33 0.28 75.33 1.64 74.63 1.64 74.63 0.28 74.41 0.28 74.41 1.64 73.71 1.64 73.71 0.28 73.49 0.28 73.49 1.64 72.79 1.64 72.79 0.28 72.11 0.28 72.11 1.64 71.41 1.64 71.41 0.28 71.19 0.28 71.19 1.64 70.49 1.64 70.49 0.28 70.27 0.28 70.27 1.64 69.57 1.64 69.57 0.28 69.35 0.28 69.35 1.64 68.65 1.64 68.65 0.28 68.43 0.28 68.43 1.64 67.73 1.64 67.73 0.28 67.51 0.28 67.51 1.64 66.81 1.64 66.81 0.28 66.59 0.28 66.59 1.64 65.89 1.64 65.89 0.28 65.67 0.28 65.67 1.64 64.97 1.64 64.97 0.28 64.75 0.28 64.75 1.64 64.05 1.64 64.05 0.28 63.83 0.28 63.83 1.64 63.13 1.64 63.13 0.28 62.91 0.28 62.91 1.64 62.21 1.64 62.21 0.28 61.99 0.28 61.99 1.64 61.29 1.64 61.29 0.28 61.07 0.28 61.07 1.64 60.37 1.64 60.37 0.28 60.15 0.28 60.15 1.64 59.45 1.64 59.45 0.28 59.23 0.28 59.23 1.64 58.53 1.64 58.53 0.28 57.85 0.28 57.85 1.64 57.15 1.64 57.15 0.28 55.55 0.28 55.55 1.64 54.85 1.64 54.85 0.28 54.63 0.28 54.63 1.64 53.93 1.64 53.93 0.28 53.71 0.28 53.71 1.64 53.01 1.64 53.01 0.28 52.79 0.28 52.79 1.64 52.09 1.64 52.09 0.28 28.8 0.28 28.8 27.48 2.65 27.48 2.65 28.84 1.95 28.84 1.95 27.48 0.28 27.48 0.28 103.08 1.95 103.08 1.95 101.72 2.65 101.72 2.65 103.08 2.87 103.08 2.87 101.72 3.57 101.72 3.57 103.08 3.79 103.08 3.79 101.72 4.49 101.72 4.49 103.08 4.71 103.08 4.71 101.72 5.41 101.72 5.41 103.08 7.01 103.08 7.01 101.72 7.71 101.72 7.71 103.08 10.23 103.08 10.23 101.72 10.93 101.72 10.93 103.08 11.15 103.08 11.15 101.72 11.85 101.72 11.85 103.08 28.8 103.08 28.8 130.28 30.47 130.28 30.47 128.92 31.17 128.92 31.17 130.28 31.39 130.28 31.39 128.92 32.09 128.92 32.09 130.28 32.31 130.28 32.31 128.92 33.01 128.92 33.01 130.28 49.79 130.28 49.79 128.92 50.49 128.92 50.49 130.28 50.71 130.28 50.71 128.92 51.41 128.92 51.41 130.28 51.63 130.28 51.63 128.92 52.33 128.92 52.33 130.28 52.55 130.28 52.55 128.92 53.25 128.92 53.25 130.28 53.47 130.28 53.47 128.92 54.17 128.92 54.17 130.28 54.39 130.28 54.39 128.92 55.09 128.92 55.09 130.28 57.15 130.28 57.15 128.92 57.85 128.92 57.85 130.28 58.07 130.28 58.07 128.92 58.77 128.92 58.77 130.28 58.99 130.28 58.99 128.92 59.69 128.92 59.69 130.28 59.91 130.28 59.91 128.92 60.61 128.92 60.61 130.28 60.83 130.28 60.83 128.92 61.53 128.92 61.53 130.28 61.75 130.28 61.75 128.92 62.45 128.92 62.45 130.28 63.13 130.28 63.13 128.92 63.83 128.92 63.83 130.28 64.05 130.28 64.05 128.92 64.75 128.92 64.75 130.28 66.35 130.28 66.35 128.92 67.05 128.92 67.05 130.28 67.27 130.28 67.27 128.92 67.97 128.92 67.97 130.28 68.19 130.28 68.19 128.92 68.89 128.92 68.89 130.28 69.11 130.28 69.11 128.92 69.81 128.92 69.81 130.28 70.03 130.28 70.03 128.92 70.73 128.92 70.73 130.28 70.95 130.28 70.95 128.92 71.65 128.92 71.65 130.28 71.87 130.28 71.87 128.92 72.57 128.92 72.57 130.28 72.79 130.28 72.79 128.92 73.49 128.92 73.49 130.28 73.71 130.28 73.71 128.92 74.41 128.92 74.41 130.28 74.63 130.28 74.63 128.92 75.33 128.92 75.33 130.28 75.55 130.28 75.55 128.92 76.25 128.92 76.25 130.28 76.47 130.28 76.47 128.92 77.17 128.92 77.17 130.28 77.39 130.28 77.39 128.92 78.09 128.92 78.09 130.28 78.31 130.28 78.31 128.92 79.01 128.92 79.01 130.28 79.23 130.28 79.23 128.92 79.93 128.92 79.93 130.28 80.15 130.28 80.15 128.92 80.85 128.92 80.85 130.28 81.07 130.28 81.07 128.92 81.77 128.92 81.77 130.28 81.99 130.28 81.99 128.92 82.69 128.92 82.69 130.28 83.37 130.28 83.37 128.92 84.07 128.92 84.07 130.28 84.29 130.28 84.29 128.92 84.99 128.92 84.99 130.28 86.59 130.28 86.59 128.92 87.29 128.92 87.29 130.28 93.49 130.28 93.49 128.92 94.19 128.92 94.19 130.28 95.33 130.28 95.33 128.92 96.03 128.92 96.03 130.28 96.25 130.28 96.25 128.92 96.95 128.92 96.95 130.28 97.17 130.28 97.17 128.92 97.87 128.92 97.87 130.28 98.55 130.28 98.55 128.92 99.25 128.92 99.25 130.28 ;
    LAYER met3 ;
      POLYGON 85.725 130.725 85.725 130.72 85.94 130.72 85.94 130.4 85.725 130.4 85.725 130.395 85.395 130.395 85.395 130.4 85.18 130.4 85.18 130.72 85.395 130.72 85.395 130.725 ;
      POLYGON 56.285 130.725 56.285 130.72 56.5 130.72 56.5 130.4 56.285 130.4 56.285 130.395 55.955 130.395 55.955 130.4 55.74 130.4 55.74 130.72 55.955 130.72 55.955 130.725 ;
      POLYGON 6.605 103.525 6.605 103.52 6.82 103.52 6.82 103.2 6.605 103.2 6.605 103.195 6.275 103.195 6.275 103.2 6.06 103.2 6.06 103.52 6.275 103.52 6.275 103.525 ;
      POLYGON 140.45 96.03 140.45 95.75 139.9 95.75 139.9 95.73 121.75 95.73 121.75 96.03 ;
      POLYGON 8.43 93.31 8.43 93.01 1.78 93.01 1.78 93.03 1.23 93.03 1.23 93.31 ;
      POLYGON 10.27 76.99 10.27 76.69 1.78 76.69 1.78 76.71 1.23 76.71 1.23 76.99 ;
      POLYGON 2.005 68.845 2.005 68.84 2.03 68.84 2.03 68.52 2.005 68.52 2.005 68.515 1.275 68.515 1.275 68.845 ;
      POLYGON 2.03 56.6 2.03 56.59 10.73 56.59 10.73 56.29 2.03 56.29 2.03 56.28 1.65 56.28 1.65 56.6 ;
      POLYGON 140.45 41.63 140.45 41.35 139.9 41.35 139.9 41.33 126.81 41.33 126.81 41.63 ;
      POLYGON 140.45 40.27 140.45 39.99 139.9 39.99 139.9 39.97 94.61 39.97 94.61 40.27 ;
      POLYGON 99.97 36.19 99.97 35.89 1.23 35.89 1.23 36.17 1.78 36.17 1.78 36.19 ;
      POLYGON 6.605 27.365 6.605 27.36 6.82 27.36 6.82 27.04 6.605 27.04 6.605 27.035 6.275 27.035 6.275 27.04 6.06 27.04 6.06 27.36 6.275 27.36 6.275 27.365 ;
      POLYGON 85.725 0.165 85.725 0.16 85.94 0.16 85.94 -0.16 85.725 -0.16 85.725 -0.165 85.395 -0.165 85.395 -0.16 85.18 -0.16 85.18 0.16 85.395 0.16 85.395 0.165 ;
      POLYGON 56.285 0.165 56.285 0.16 56.5 0.16 56.5 -0.16 56.285 -0.16 56.285 -0.165 55.955 -0.165 55.955 -0.16 55.74 -0.16 55.74 0.16 55.955 0.16 55.955 0.165 ;
      POLYGON 112.76 130.16 112.76 127.03 111.38 127.03 111.38 125.93 112.76 125.93 112.76 119.55 111.38 119.55 111.38 118.45 112.76 118.45 112.76 118.19 111.38 118.19 111.38 117.09 112.76 117.09 112.76 102.96 141.28 102.96 141.28 99.83 139.9 99.83 139.9 98.73 141.28 98.73 141.28 97.11 139.9 97.11 139.9 96.01 141.28 96.01 141.28 95.75 139.9 95.75 139.9 94.65 141.28 94.65 141.28 94.39 139.9 94.39 139.9 93.29 141.28 93.29 141.28 91.67 139.9 91.67 139.9 90.57 141.28 90.57 141.28 90.31 139.9 90.31 139.9 89.21 141.28 89.21 141.28 88.95 139.9 88.95 139.9 87.85 141.28 87.85 141.28 86.23 139.9 86.23 139.9 85.13 141.28 85.13 141.28 84.87 139.9 84.87 139.9 83.77 141.28 83.77 141.28 83.51 139.9 83.51 139.9 82.41 141.28 82.41 141.28 80.79 139.9 80.79 139.9 79.69 141.28 79.69 141.28 79.43 139.9 79.43 139.9 78.33 141.28 78.33 141.28 78.07 139.9 78.07 139.9 76.97 141.28 76.97 141.28 74.67 139.9 74.67 139.9 73.57 141.28 73.57 141.28 72.63 139.9 72.63 139.9 71.53 141.28 71.53 141.28 69.91 139.9 69.91 139.9 68.81 141.28 68.81 141.28 68.55 139.9 68.55 139.9 67.45 141.28 67.45 141.28 67.19 139.9 67.19 139.9 66.09 141.28 66.09 141.28 65.83 139.9 65.83 139.9 64.73 141.28 64.73 141.28 64.47 139.9 64.47 139.9 63.37 141.28 63.37 141.28 63.11 139.9 63.11 139.9 62.01 141.28 62.01 141.28 61.75 139.9 61.75 139.9 60.65 141.28 60.65 141.28 59.03 139.9 59.03 139.9 57.93 141.28 57.93 141.28 57.67 139.9 57.67 139.9 56.57 141.28 56.57 141.28 56.31 139.9 56.31 139.9 55.21 141.28 55.21 141.28 52.91 139.9 52.91 139.9 51.81 141.28 51.81 141.28 51.55 139.9 51.55 139.9 50.45 141.28 50.45 141.28 49.51 139.9 49.51 139.9 48.41 141.28 48.41 141.28 48.15 139.9 48.15 139.9 47.05 141.28 47.05 141.28 46.79 139.9 46.79 139.9 45.69 141.28 45.69 141.28 45.43 139.9 45.43 139.9 44.33 141.28 44.33 141.28 44.07 139.9 44.07 139.9 42.97 141.28 42.97 141.28 42.71 139.9 42.71 139.9 41.61 141.28 41.61 141.28 41.35 139.9 41.35 139.9 40.25 141.28 40.25 141.28 39.99 139.9 39.99 139.9 38.89 141.28 38.89 141.28 38.63 139.9 38.63 139.9 37.53 141.28 37.53 141.28 37.27 139.9 37.27 139.9 36.17 141.28 36.17 141.28 35.91 139.9 35.91 139.9 34.81 141.28 34.81 141.28 34.55 139.9 34.55 139.9 33.45 141.28 33.45 141.28 33.19 139.9 33.19 139.9 32.09 141.28 32.09 141.28 31.83 139.9 31.83 139.9 30.73 141.28 30.73 141.28 27.6 112.76 27.6 112.76 0.4 28.92 0.4 28.92 2.85 30.3 2.85 30.3 3.95 28.92 3.95 28.92 4.21 30.3 4.21 30.3 5.31 28.92 5.31 28.92 6.25 30.3 6.25 30.3 7.35 28.92 7.35 28.92 7.61 30.3 7.61 30.3 8.71 28.92 8.71 28.92 9.65 30.3 9.65 30.3 10.75 28.92 10.75 28.92 11.01 30.3 11.01 30.3 12.11 28.92 12.11 28.92 12.37 30.3 12.37 30.3 13.47 28.92 13.47 28.92 13.73 30.3 13.73 30.3 14.83 28.92 14.83 28.92 27.6 0.4 27.6 0.4 31.41 1.78 31.41 1.78 32.51 0.4 32.51 0.4 33.45 1.78 33.45 1.78 34.55 0.4 34.55 0.4 34.81 1.78 34.81 1.78 35.91 0.4 35.91 0.4 36.17 1.78 36.17 1.78 37.27 0.4 37.27 0.4 37.53 1.78 37.53 1.78 38.63 0.4 38.63 0.4 38.89 1.78 38.89 1.78 39.99 0.4 39.99 0.4 40.25 1.78 40.25 1.78 41.35 0.4 41.35 0.4 41.61 1.78 41.61 1.78 42.71 0.4 42.71 0.4 42.97 1.78 42.97 1.78 44.07 0.4 44.07 0.4 44.33 1.78 44.33 1.78 45.43 0.4 45.43 0.4 45.69 1.78 45.69 1.78 46.79 0.4 46.79 0.4 47.05 1.78 47.05 1.78 48.15 0.4 48.15 0.4 48.41 1.78 48.41 1.78 49.51 0.4 49.51 0.4 49.77 1.78 49.77 1.78 50.87 0.4 50.87 0.4 51.13 1.78 51.13 1.78 52.23 0.4 52.23 0.4 52.49 1.78 52.49 1.78 53.59 0.4 53.59 0.4 53.85 1.78 53.85 1.78 54.95 0.4 54.95 0.4 55.21 1.78 55.21 1.78 56.31 0.4 56.31 0.4 58.61 1.78 58.61 1.78 59.71 0.4 59.71 0.4 60.65 1.78 60.65 1.78 61.75 0.4 61.75 0.4 64.05 1.78 64.05 1.78 65.15 0.4 65.15 0.4 65.41 1.78 65.41 1.78 66.51 0.4 66.51 0.4 67.45 1.78 67.45 1.78 68.55 0.4 68.55 0.4 68.81 1.78 68.81 1.78 69.91 0.4 69.91 0.4 70.17 1.78 70.17 1.78 71.27 0.4 71.27 0.4 71.53 1.78 71.53 1.78 72.63 0.4 72.63 0.4 74.25 1.78 74.25 1.78 75.35 0.4 75.35 0.4 75.61 1.78 75.61 1.78 76.71 0.4 76.71 0.4 76.97 1.78 76.97 1.78 78.07 0.4 78.07 0.4 79.69 1.78 79.69 1.78 80.79 0.4 80.79 0.4 81.05 1.78 81.05 1.78 82.15 0.4 82.15 0.4 82.41 1.78 82.41 1.78 83.51 0.4 83.51 0.4 85.13 1.78 85.13 1.78 86.23 0.4 86.23 0.4 86.49 1.78 86.49 1.78 87.59 0.4 87.59 0.4 87.85 1.78 87.85 1.78 88.95 0.4 88.95 0.4 90.57 1.78 90.57 1.78 91.67 0.4 91.67 0.4 91.93 1.78 91.93 1.78 93.03 0.4 93.03 0.4 93.29 1.78 93.29 1.78 94.39 0.4 94.39 0.4 96.01 1.78 96.01 1.78 97.11 0.4 97.11 0.4 97.37 1.78 97.37 1.78 98.47 0.4 98.47 0.4 98.73 1.78 98.73 1.78 99.83 0.4 99.83 0.4 102.96 28.92 102.96 28.92 117.09 30.3 117.09 30.3 118.19 28.92 118.19 28.92 118.45 30.3 118.45 30.3 119.55 28.92 119.55 28.92 121.85 30.3 121.85 30.3 122.95 28.92 122.95 28.92 123.21 30.3 123.21 30.3 124.31 28.92 124.31 28.92 124.57 30.3 124.57 30.3 125.67 28.92 125.67 28.92 126.61 30.3 126.61 30.3 127.71 28.92 127.71 28.92 130.16 ;
    LAYER met4 ;
      POLYGON 112.76 130.16 112.76 102.96 134.54 102.96 134.54 102.36 135.94 102.36 135.94 102.96 141.28 102.96 141.28 27.6 135.94 27.6 135.94 28.2 134.54 28.2 134.54 27.6 112.76 27.6 112.76 0.4 100.98 0.4 100.98 1 99.58 1 99.58 0.4 86.26 0.4 86.26 1 84.86 1 84.86 0.4 71.54 0.4 71.54 1 70.14 1 70.14 0.4 56.82 0.4 56.82 1 55.42 1 55.42 0.4 42.1 0.4 42.1 1 40.7 1 40.7 0.4 28.92 0.4 28.92 27.6 7.14 27.6 7.14 28.2 5.74 28.2 5.74 27.6 0.4 27.6 0.4 102.96 5.74 102.96 5.74 102.36 7.14 102.36 7.14 102.96 28.92 102.96 28.92 130.16 40.7 130.16 40.7 129.56 42.1 129.56 42.1 130.16 55.42 130.16 55.42 129.56 56.82 129.56 56.82 130.16 70.14 130.16 70.14 129.56 71.54 129.56 71.54 130.16 84.86 130.16 84.86 129.56 86.26 129.56 86.26 130.16 99.58 130.16 99.58 129.56 100.98 129.56 100.98 130.16 ;
    LAYER met5 ;
      POLYGON 106.76 127.36 106.76 119.64 109.96 119.64 109.96 100.16 138.48 100.16 138.48 90.48 135.28 90.48 135.28 80.88 138.48 80.88 138.48 70.08 135.28 70.08 135.28 60.48 138.48 60.48 138.48 49.68 135.28 49.68 135.28 40.08 138.48 40.08 138.48 30.4 109.96 30.4 109.96 10.92 106.76 10.92 106.76 3.2 34.92 3.2 34.92 10.92 31.72 10.92 31.72 30.4 3.2 30.4 3.2 40.08 6.4 40.08 6.4 49.68 3.2 49.68 3.2 60.48 6.4 60.48 6.4 70.08 3.2 70.08 3.2 80.88 6.4 80.88 6.4 90.48 3.2 90.48 3.2 100.16 31.72 100.16 31.72 119.64 34.92 119.64 34.92 127.36 ;
    LAYER met1 ;
      POLYGON 112.88 130.04 112.88 128.36 112.4 128.36 112.4 127.32 112.88 127.32 112.88 125.64 112.4 125.64 112.4 124.6 112.88 124.6 112.88 122.92 112.4 122.92 112.4 121.88 112.88 121.88 112.88 120.2 112.4 120.2 112.4 119.16 112.88 119.16 112.88 117.48 112.4 117.48 112.4 116.44 112.88 116.44 112.88 114.76 112.4 114.76 112.4 113.72 112.88 113.72 112.88 112.04 112.4 112.04 112.4 111 112.88 111 112.88 109.32 112.4 109.32 112.4 108.28 112.88 108.28 112.88 106.6 112.4 106.6 112.4 105.56 112.88 105.56 112.88 103.88 28.8 103.88 28.8 105.56 29.28 105.56 29.28 106.6 28.8 106.6 28.8 108.28 29.28 108.28 29.28 109.32 28.8 109.32 28.8 111 29.28 111 29.28 112.04 28.8 112.04 28.8 113.72 29.28 113.72 29.28 114.76 28.8 114.76 28.8 116.44 29.28 116.44 29.28 117.48 28.8 117.48 28.8 119.16 29.28 119.16 29.28 120.2 28.8 120.2 28.8 121.88 29.28 121.88 29.28 122.92 28.8 122.92 28.8 124.6 29.28 124.6 29.28 125.64 28.8 125.64 28.8 127.32 29.28 127.32 29.28 128.36 28.8 128.36 28.8 130.04 ;
      POLYGON 141.4 102.84 141.4 101.16 140.92 101.16 140.92 100.12 141.4 100.12 141.4 98.44 140.92 98.44 140.92 97.4 141.4 97.4 141.4 95.72 140.92 95.72 140.92 94.68 141.4 94.68 141.4 93 140.92 93 140.92 91.96 141.4 91.96 141.4 90.28 140.92 90.28 140.92 89.24 141.4 89.24 141.4 87.56 140.92 87.56 140.92 86.52 141.4 86.52 141.4 84.84 140.92 84.84 140.92 83.8 141.4 83.8 141.4 82.12 140.92 82.12 140.92 81.08 141.4 81.08 141.4 79.4 140.92 79.4 140.92 78.36 141.4 78.36 141.4 76.68 140.92 76.68 140.92 75.64 141.4 75.64 141.4 73.96 140.92 73.96 140.92 72.92 141.4 72.92 141.4 71.24 140.92 71.24 140.92 70.2 141.4 70.2 141.4 68.52 140.92 68.52 140.92 67.48 141.4 67.48 141.4 65.8 140.92 65.8 140.92 64.76 141.4 64.76 141.4 63.08 140.92 63.08 140.92 62.04 141.4 62.04 141.4 60.36 140.92 60.36 140.92 59.32 141.4 59.32 141.4 57.64 140.92 57.64 140.92 56.6 141.4 56.6 141.4 54.92 140.92 54.92 140.92 53.88 141.4 53.88 141.4 52.2 140.92 52.2 140.92 51.16 141.4 51.16 141.4 49.48 140.92 49.48 140.92 48.44 141.4 48.44 141.4 46.76 140.92 46.76 140.92 45.72 141.4 45.72 141.4 44.04 140.92 44.04 140.92 43 141.4 43 141.4 41.32 140.92 41.32 140.92 40.28 141.4 40.28 141.4 38.6 140.92 38.6 140.92 37.56 141.4 37.56 141.4 35.88 140.92 35.88 140.92 34.84 141.4 34.84 141.4 33.16 140.92 33.16 140.92 32.12 141.4 32.12 141.4 30.44 140.92 30.44 140.92 29.4 141.4 29.4 141.4 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 0.76 97.4 0.76 98.44 0.28 98.44 0.28 100.12 0.76 100.12 0.76 101.16 0.28 101.16 0.28 102.84 ;
      POLYGON 112.88 26.68 112.88 25 112.4 25 112.4 23.96 112.88 23.96 112.88 22.28 112.4 22.28 112.4 21.24 112.88 21.24 112.88 19.56 112.4 19.56 112.4 18.52 112.88 18.52 112.88 16.84 112.4 16.84 112.4 15.8 112.88 15.8 112.88 14.12 112.4 14.12 112.4 13.08 112.88 13.08 112.88 11.4 112.4 11.4 112.4 10.36 112.88 10.36 112.88 8.68 112.4 8.68 112.4 7.64 112.88 7.64 112.88 5.96 112.4 5.96 112.4 4.92 112.88 4.92 112.88 3.24 112.4 3.24 112.4 2.2 112.88 2.2 112.88 0.52 28.8 0.52 28.8 2.2 29.28 2.2 29.28 3.24 28.8 3.24 28.8 4.92 29.28 4.92 29.28 5.96 28.8 5.96 28.8 7.64 29.28 7.64 29.28 8.68 28.8 8.68 28.8 10.36 29.28 10.36 29.28 11.4 28.8 11.4 28.8 13.08 29.28 13.08 29.28 14.12 28.8 14.12 28.8 15.8 29.28 15.8 29.28 16.84 28.8 16.84 28.8 18.52 29.28 18.52 29.28 19.56 28.8 19.56 28.8 21.24 29.28 21.24 29.28 22.28 28.8 22.28 28.8 23.96 29.28 23.96 29.28 25 28.8 25 28.8 26.68 ;
    LAYER li1 ;
      POLYGON 112.82 130.22 112.82 103.02 141.34 103.02 141.34 27.54 112.82 27.54 112.82 0.34 28.86 0.34 28.86 27.54 0.34 27.54 0.34 103.02 28.86 103.02 28.86 130.22 ;
    LAYER mcon ;
      RECT 112.845 130.475 113.015 130.645 ;
      RECT 112.385 130.475 112.555 130.645 ;
      RECT 111.925 130.475 112.095 130.645 ;
      RECT 111.465 130.475 111.635 130.645 ;
      RECT 111.005 130.475 111.175 130.645 ;
      RECT 110.545 130.475 110.715 130.645 ;
      RECT 110.085 130.475 110.255 130.645 ;
      RECT 109.625 130.475 109.795 130.645 ;
      RECT 109.165 130.475 109.335 130.645 ;
      RECT 108.705 130.475 108.875 130.645 ;
      RECT 108.245 130.475 108.415 130.645 ;
      RECT 107.785 130.475 107.955 130.645 ;
      RECT 107.325 130.475 107.495 130.645 ;
      RECT 106.865 130.475 107.035 130.645 ;
      RECT 106.405 130.475 106.575 130.645 ;
      RECT 105.945 130.475 106.115 130.645 ;
      RECT 105.485 130.475 105.655 130.645 ;
      RECT 105.025 130.475 105.195 130.645 ;
      RECT 104.565 130.475 104.735 130.645 ;
      RECT 104.105 130.475 104.275 130.645 ;
      RECT 103.645 130.475 103.815 130.645 ;
      RECT 103.185 130.475 103.355 130.645 ;
      RECT 102.725 130.475 102.895 130.645 ;
      RECT 102.265 130.475 102.435 130.645 ;
      RECT 101.805 130.475 101.975 130.645 ;
      RECT 101.345 130.475 101.515 130.645 ;
      RECT 100.885 130.475 101.055 130.645 ;
      RECT 100.425 130.475 100.595 130.645 ;
      RECT 99.965 130.475 100.135 130.645 ;
      RECT 99.505 130.475 99.675 130.645 ;
      RECT 99.045 130.475 99.215 130.645 ;
      RECT 98.585 130.475 98.755 130.645 ;
      RECT 98.125 130.475 98.295 130.645 ;
      RECT 97.665 130.475 97.835 130.645 ;
      RECT 97.205 130.475 97.375 130.645 ;
      RECT 96.745 130.475 96.915 130.645 ;
      RECT 96.285 130.475 96.455 130.645 ;
      RECT 95.825 130.475 95.995 130.645 ;
      RECT 95.365 130.475 95.535 130.645 ;
      RECT 94.905 130.475 95.075 130.645 ;
      RECT 94.445 130.475 94.615 130.645 ;
      RECT 93.985 130.475 94.155 130.645 ;
      RECT 93.525 130.475 93.695 130.645 ;
      RECT 93.065 130.475 93.235 130.645 ;
      RECT 92.605 130.475 92.775 130.645 ;
      RECT 92.145 130.475 92.315 130.645 ;
      RECT 91.685 130.475 91.855 130.645 ;
      RECT 91.225 130.475 91.395 130.645 ;
      RECT 90.765 130.475 90.935 130.645 ;
      RECT 90.305 130.475 90.475 130.645 ;
      RECT 89.845 130.475 90.015 130.645 ;
      RECT 89.385 130.475 89.555 130.645 ;
      RECT 88.925 130.475 89.095 130.645 ;
      RECT 88.465 130.475 88.635 130.645 ;
      RECT 88.005 130.475 88.175 130.645 ;
      RECT 87.545 130.475 87.715 130.645 ;
      RECT 87.085 130.475 87.255 130.645 ;
      RECT 86.625 130.475 86.795 130.645 ;
      RECT 86.165 130.475 86.335 130.645 ;
      RECT 85.705 130.475 85.875 130.645 ;
      RECT 85.245 130.475 85.415 130.645 ;
      RECT 84.785 130.475 84.955 130.645 ;
      RECT 84.325 130.475 84.495 130.645 ;
      RECT 83.865 130.475 84.035 130.645 ;
      RECT 83.405 130.475 83.575 130.645 ;
      RECT 82.945 130.475 83.115 130.645 ;
      RECT 82.485 130.475 82.655 130.645 ;
      RECT 82.025 130.475 82.195 130.645 ;
      RECT 81.565 130.475 81.735 130.645 ;
      RECT 81.105 130.475 81.275 130.645 ;
      RECT 80.645 130.475 80.815 130.645 ;
      RECT 80.185 130.475 80.355 130.645 ;
      RECT 79.725 130.475 79.895 130.645 ;
      RECT 79.265 130.475 79.435 130.645 ;
      RECT 78.805 130.475 78.975 130.645 ;
      RECT 78.345 130.475 78.515 130.645 ;
      RECT 77.885 130.475 78.055 130.645 ;
      RECT 77.425 130.475 77.595 130.645 ;
      RECT 76.965 130.475 77.135 130.645 ;
      RECT 76.505 130.475 76.675 130.645 ;
      RECT 76.045 130.475 76.215 130.645 ;
      RECT 75.585 130.475 75.755 130.645 ;
      RECT 75.125 130.475 75.295 130.645 ;
      RECT 74.665 130.475 74.835 130.645 ;
      RECT 74.205 130.475 74.375 130.645 ;
      RECT 73.745 130.475 73.915 130.645 ;
      RECT 73.285 130.475 73.455 130.645 ;
      RECT 72.825 130.475 72.995 130.645 ;
      RECT 72.365 130.475 72.535 130.645 ;
      RECT 71.905 130.475 72.075 130.645 ;
      RECT 71.445 130.475 71.615 130.645 ;
      RECT 70.985 130.475 71.155 130.645 ;
      RECT 70.525 130.475 70.695 130.645 ;
      RECT 70.065 130.475 70.235 130.645 ;
      RECT 69.605 130.475 69.775 130.645 ;
      RECT 69.145 130.475 69.315 130.645 ;
      RECT 68.685 130.475 68.855 130.645 ;
      RECT 68.225 130.475 68.395 130.645 ;
      RECT 67.765 130.475 67.935 130.645 ;
      RECT 67.305 130.475 67.475 130.645 ;
      RECT 66.845 130.475 67.015 130.645 ;
      RECT 66.385 130.475 66.555 130.645 ;
      RECT 65.925 130.475 66.095 130.645 ;
      RECT 65.465 130.475 65.635 130.645 ;
      RECT 65.005 130.475 65.175 130.645 ;
      RECT 64.545 130.475 64.715 130.645 ;
      RECT 64.085 130.475 64.255 130.645 ;
      RECT 63.625 130.475 63.795 130.645 ;
      RECT 63.165 130.475 63.335 130.645 ;
      RECT 62.705 130.475 62.875 130.645 ;
      RECT 62.245 130.475 62.415 130.645 ;
      RECT 61.785 130.475 61.955 130.645 ;
      RECT 61.325 130.475 61.495 130.645 ;
      RECT 60.865 130.475 61.035 130.645 ;
      RECT 60.405 130.475 60.575 130.645 ;
      RECT 59.945 130.475 60.115 130.645 ;
      RECT 59.485 130.475 59.655 130.645 ;
      RECT 59.025 130.475 59.195 130.645 ;
      RECT 58.565 130.475 58.735 130.645 ;
      RECT 58.105 130.475 58.275 130.645 ;
      RECT 57.645 130.475 57.815 130.645 ;
      RECT 57.185 130.475 57.355 130.645 ;
      RECT 56.725 130.475 56.895 130.645 ;
      RECT 56.265 130.475 56.435 130.645 ;
      RECT 55.805 130.475 55.975 130.645 ;
      RECT 55.345 130.475 55.515 130.645 ;
      RECT 54.885 130.475 55.055 130.645 ;
      RECT 54.425 130.475 54.595 130.645 ;
      RECT 53.965 130.475 54.135 130.645 ;
      RECT 53.505 130.475 53.675 130.645 ;
      RECT 53.045 130.475 53.215 130.645 ;
      RECT 52.585 130.475 52.755 130.645 ;
      RECT 52.125 130.475 52.295 130.645 ;
      RECT 51.665 130.475 51.835 130.645 ;
      RECT 51.205 130.475 51.375 130.645 ;
      RECT 50.745 130.475 50.915 130.645 ;
      RECT 50.285 130.475 50.455 130.645 ;
      RECT 49.825 130.475 49.995 130.645 ;
      RECT 49.365 130.475 49.535 130.645 ;
      RECT 48.905 130.475 49.075 130.645 ;
      RECT 48.445 130.475 48.615 130.645 ;
      RECT 47.985 130.475 48.155 130.645 ;
      RECT 47.525 130.475 47.695 130.645 ;
      RECT 47.065 130.475 47.235 130.645 ;
      RECT 46.605 130.475 46.775 130.645 ;
      RECT 46.145 130.475 46.315 130.645 ;
      RECT 45.685 130.475 45.855 130.645 ;
      RECT 45.225 130.475 45.395 130.645 ;
      RECT 44.765 130.475 44.935 130.645 ;
      RECT 44.305 130.475 44.475 130.645 ;
      RECT 43.845 130.475 44.015 130.645 ;
      RECT 43.385 130.475 43.555 130.645 ;
      RECT 42.925 130.475 43.095 130.645 ;
      RECT 42.465 130.475 42.635 130.645 ;
      RECT 42.005 130.475 42.175 130.645 ;
      RECT 41.545 130.475 41.715 130.645 ;
      RECT 41.085 130.475 41.255 130.645 ;
      RECT 40.625 130.475 40.795 130.645 ;
      RECT 40.165 130.475 40.335 130.645 ;
      RECT 39.705 130.475 39.875 130.645 ;
      RECT 39.245 130.475 39.415 130.645 ;
      RECT 38.785 130.475 38.955 130.645 ;
      RECT 38.325 130.475 38.495 130.645 ;
      RECT 37.865 130.475 38.035 130.645 ;
      RECT 37.405 130.475 37.575 130.645 ;
      RECT 36.945 130.475 37.115 130.645 ;
      RECT 36.485 130.475 36.655 130.645 ;
      RECT 36.025 130.475 36.195 130.645 ;
      RECT 35.565 130.475 35.735 130.645 ;
      RECT 35.105 130.475 35.275 130.645 ;
      RECT 34.645 130.475 34.815 130.645 ;
      RECT 34.185 130.475 34.355 130.645 ;
      RECT 33.725 130.475 33.895 130.645 ;
      RECT 33.265 130.475 33.435 130.645 ;
      RECT 32.805 130.475 32.975 130.645 ;
      RECT 32.345 130.475 32.515 130.645 ;
      RECT 31.885 130.475 32.055 130.645 ;
      RECT 31.425 130.475 31.595 130.645 ;
      RECT 30.965 130.475 31.135 130.645 ;
      RECT 30.505 130.475 30.675 130.645 ;
      RECT 30.045 130.475 30.215 130.645 ;
      RECT 29.585 130.475 29.755 130.645 ;
      RECT 29.125 130.475 29.295 130.645 ;
      RECT 28.665 130.475 28.835 130.645 ;
      RECT 112.845 127.755 113.015 127.925 ;
      RECT 112.385 127.755 112.555 127.925 ;
      RECT 29.125 127.755 29.295 127.925 ;
      RECT 28.665 127.755 28.835 127.925 ;
      RECT 112.845 125.035 113.015 125.205 ;
      RECT 112.385 125.035 112.555 125.205 ;
      RECT 29.125 125.035 29.295 125.205 ;
      RECT 28.665 125.035 28.835 125.205 ;
      RECT 112.845 122.315 113.015 122.485 ;
      RECT 112.385 122.315 112.555 122.485 ;
      RECT 29.125 122.315 29.295 122.485 ;
      RECT 28.665 122.315 28.835 122.485 ;
      RECT 112.845 119.595 113.015 119.765 ;
      RECT 112.385 119.595 112.555 119.765 ;
      RECT 29.125 119.595 29.295 119.765 ;
      RECT 28.665 119.595 28.835 119.765 ;
      RECT 112.845 116.875 113.015 117.045 ;
      RECT 112.385 116.875 112.555 117.045 ;
      RECT 29.125 116.875 29.295 117.045 ;
      RECT 28.665 116.875 28.835 117.045 ;
      RECT 112.845 114.155 113.015 114.325 ;
      RECT 112.385 114.155 112.555 114.325 ;
      RECT 29.125 114.155 29.295 114.325 ;
      RECT 28.665 114.155 28.835 114.325 ;
      RECT 112.845 111.435 113.015 111.605 ;
      RECT 112.385 111.435 112.555 111.605 ;
      RECT 29.125 111.435 29.295 111.605 ;
      RECT 28.665 111.435 28.835 111.605 ;
      RECT 112.845 108.715 113.015 108.885 ;
      RECT 112.385 108.715 112.555 108.885 ;
      RECT 29.125 108.715 29.295 108.885 ;
      RECT 28.665 108.715 28.835 108.885 ;
      RECT 112.845 105.995 113.015 106.165 ;
      RECT 112.385 105.995 112.555 106.165 ;
      RECT 29.125 105.995 29.295 106.165 ;
      RECT 28.665 105.995 28.835 106.165 ;
      RECT 141.365 103.275 141.535 103.445 ;
      RECT 140.905 103.275 141.075 103.445 ;
      RECT 140.445 103.275 140.615 103.445 ;
      RECT 139.985 103.275 140.155 103.445 ;
      RECT 139.525 103.275 139.695 103.445 ;
      RECT 139.065 103.275 139.235 103.445 ;
      RECT 138.605 103.275 138.775 103.445 ;
      RECT 138.145 103.275 138.315 103.445 ;
      RECT 137.685 103.275 137.855 103.445 ;
      RECT 137.225 103.275 137.395 103.445 ;
      RECT 136.765 103.275 136.935 103.445 ;
      RECT 136.305 103.275 136.475 103.445 ;
      RECT 135.845 103.275 136.015 103.445 ;
      RECT 135.385 103.275 135.555 103.445 ;
      RECT 134.925 103.275 135.095 103.445 ;
      RECT 134.465 103.275 134.635 103.445 ;
      RECT 134.005 103.275 134.175 103.445 ;
      RECT 133.545 103.275 133.715 103.445 ;
      RECT 133.085 103.275 133.255 103.445 ;
      RECT 132.625 103.275 132.795 103.445 ;
      RECT 132.165 103.275 132.335 103.445 ;
      RECT 131.705 103.275 131.875 103.445 ;
      RECT 131.245 103.275 131.415 103.445 ;
      RECT 130.785 103.275 130.955 103.445 ;
      RECT 130.325 103.275 130.495 103.445 ;
      RECT 129.865 103.275 130.035 103.445 ;
      RECT 129.405 103.275 129.575 103.445 ;
      RECT 128.945 103.275 129.115 103.445 ;
      RECT 128.485 103.275 128.655 103.445 ;
      RECT 128.025 103.275 128.195 103.445 ;
      RECT 127.565 103.275 127.735 103.445 ;
      RECT 127.105 103.275 127.275 103.445 ;
      RECT 126.645 103.275 126.815 103.445 ;
      RECT 126.185 103.275 126.355 103.445 ;
      RECT 125.725 103.275 125.895 103.445 ;
      RECT 125.265 103.275 125.435 103.445 ;
      RECT 124.805 103.275 124.975 103.445 ;
      RECT 124.345 103.275 124.515 103.445 ;
      RECT 123.885 103.275 124.055 103.445 ;
      RECT 123.425 103.275 123.595 103.445 ;
      RECT 122.965 103.275 123.135 103.445 ;
      RECT 122.505 103.275 122.675 103.445 ;
      RECT 122.045 103.275 122.215 103.445 ;
      RECT 121.585 103.275 121.755 103.445 ;
      RECT 121.125 103.275 121.295 103.445 ;
      RECT 120.665 103.275 120.835 103.445 ;
      RECT 120.205 103.275 120.375 103.445 ;
      RECT 119.745 103.275 119.915 103.445 ;
      RECT 119.285 103.275 119.455 103.445 ;
      RECT 118.825 103.275 118.995 103.445 ;
      RECT 118.365 103.275 118.535 103.445 ;
      RECT 117.905 103.275 118.075 103.445 ;
      RECT 117.445 103.275 117.615 103.445 ;
      RECT 116.985 103.275 117.155 103.445 ;
      RECT 116.525 103.275 116.695 103.445 ;
      RECT 116.065 103.275 116.235 103.445 ;
      RECT 115.605 103.275 115.775 103.445 ;
      RECT 115.145 103.275 115.315 103.445 ;
      RECT 114.685 103.275 114.855 103.445 ;
      RECT 114.225 103.275 114.395 103.445 ;
      RECT 113.765 103.275 113.935 103.445 ;
      RECT 113.305 103.275 113.475 103.445 ;
      RECT 112.845 103.275 113.015 103.445 ;
      RECT 112.385 103.275 112.555 103.445 ;
      RECT 111.925 103.275 112.095 103.445 ;
      RECT 111.465 103.275 111.635 103.445 ;
      RECT 111.005 103.275 111.175 103.445 ;
      RECT 110.545 103.275 110.715 103.445 ;
      RECT 110.085 103.275 110.255 103.445 ;
      RECT 109.625 103.275 109.795 103.445 ;
      RECT 109.165 103.275 109.335 103.445 ;
      RECT 108.705 103.275 108.875 103.445 ;
      RECT 108.245 103.275 108.415 103.445 ;
      RECT 107.785 103.275 107.955 103.445 ;
      RECT 107.325 103.275 107.495 103.445 ;
      RECT 106.865 103.275 107.035 103.445 ;
      RECT 106.405 103.275 106.575 103.445 ;
      RECT 105.945 103.275 106.115 103.445 ;
      RECT 105.485 103.275 105.655 103.445 ;
      RECT 105.025 103.275 105.195 103.445 ;
      RECT 104.565 103.275 104.735 103.445 ;
      RECT 104.105 103.275 104.275 103.445 ;
      RECT 103.645 103.275 103.815 103.445 ;
      RECT 103.185 103.275 103.355 103.445 ;
      RECT 102.725 103.275 102.895 103.445 ;
      RECT 102.265 103.275 102.435 103.445 ;
      RECT 101.805 103.275 101.975 103.445 ;
      RECT 101.345 103.275 101.515 103.445 ;
      RECT 100.885 103.275 101.055 103.445 ;
      RECT 100.425 103.275 100.595 103.445 ;
      RECT 99.965 103.275 100.135 103.445 ;
      RECT 99.505 103.275 99.675 103.445 ;
      RECT 99.045 103.275 99.215 103.445 ;
      RECT 98.585 103.275 98.755 103.445 ;
      RECT 98.125 103.275 98.295 103.445 ;
      RECT 97.665 103.275 97.835 103.445 ;
      RECT 97.205 103.275 97.375 103.445 ;
      RECT 96.745 103.275 96.915 103.445 ;
      RECT 96.285 103.275 96.455 103.445 ;
      RECT 95.825 103.275 95.995 103.445 ;
      RECT 95.365 103.275 95.535 103.445 ;
      RECT 94.905 103.275 95.075 103.445 ;
      RECT 94.445 103.275 94.615 103.445 ;
      RECT 93.985 103.275 94.155 103.445 ;
      RECT 93.525 103.275 93.695 103.445 ;
      RECT 93.065 103.275 93.235 103.445 ;
      RECT 92.605 103.275 92.775 103.445 ;
      RECT 92.145 103.275 92.315 103.445 ;
      RECT 91.685 103.275 91.855 103.445 ;
      RECT 91.225 103.275 91.395 103.445 ;
      RECT 90.765 103.275 90.935 103.445 ;
      RECT 90.305 103.275 90.475 103.445 ;
      RECT 89.845 103.275 90.015 103.445 ;
      RECT 89.385 103.275 89.555 103.445 ;
      RECT 88.925 103.275 89.095 103.445 ;
      RECT 88.465 103.275 88.635 103.445 ;
      RECT 88.005 103.275 88.175 103.445 ;
      RECT 87.545 103.275 87.715 103.445 ;
      RECT 87.085 103.275 87.255 103.445 ;
      RECT 86.625 103.275 86.795 103.445 ;
      RECT 86.165 103.275 86.335 103.445 ;
      RECT 85.705 103.275 85.875 103.445 ;
      RECT 85.245 103.275 85.415 103.445 ;
      RECT 84.785 103.275 84.955 103.445 ;
      RECT 84.325 103.275 84.495 103.445 ;
      RECT 83.865 103.275 84.035 103.445 ;
      RECT 83.405 103.275 83.575 103.445 ;
      RECT 82.945 103.275 83.115 103.445 ;
      RECT 82.485 103.275 82.655 103.445 ;
      RECT 82.025 103.275 82.195 103.445 ;
      RECT 81.565 103.275 81.735 103.445 ;
      RECT 81.105 103.275 81.275 103.445 ;
      RECT 80.645 103.275 80.815 103.445 ;
      RECT 80.185 103.275 80.355 103.445 ;
      RECT 79.725 103.275 79.895 103.445 ;
      RECT 79.265 103.275 79.435 103.445 ;
      RECT 78.805 103.275 78.975 103.445 ;
      RECT 78.345 103.275 78.515 103.445 ;
      RECT 77.885 103.275 78.055 103.445 ;
      RECT 77.425 103.275 77.595 103.445 ;
      RECT 76.965 103.275 77.135 103.445 ;
      RECT 76.505 103.275 76.675 103.445 ;
      RECT 76.045 103.275 76.215 103.445 ;
      RECT 75.585 103.275 75.755 103.445 ;
      RECT 75.125 103.275 75.295 103.445 ;
      RECT 74.665 103.275 74.835 103.445 ;
      RECT 74.205 103.275 74.375 103.445 ;
      RECT 73.745 103.275 73.915 103.445 ;
      RECT 73.285 103.275 73.455 103.445 ;
      RECT 72.825 103.275 72.995 103.445 ;
      RECT 72.365 103.275 72.535 103.445 ;
      RECT 71.905 103.275 72.075 103.445 ;
      RECT 71.445 103.275 71.615 103.445 ;
      RECT 70.985 103.275 71.155 103.445 ;
      RECT 70.525 103.275 70.695 103.445 ;
      RECT 70.065 103.275 70.235 103.445 ;
      RECT 69.605 103.275 69.775 103.445 ;
      RECT 69.145 103.275 69.315 103.445 ;
      RECT 68.685 103.275 68.855 103.445 ;
      RECT 68.225 103.275 68.395 103.445 ;
      RECT 67.765 103.275 67.935 103.445 ;
      RECT 67.305 103.275 67.475 103.445 ;
      RECT 66.845 103.275 67.015 103.445 ;
      RECT 66.385 103.275 66.555 103.445 ;
      RECT 65.925 103.275 66.095 103.445 ;
      RECT 65.465 103.275 65.635 103.445 ;
      RECT 65.005 103.275 65.175 103.445 ;
      RECT 64.545 103.275 64.715 103.445 ;
      RECT 64.085 103.275 64.255 103.445 ;
      RECT 63.625 103.275 63.795 103.445 ;
      RECT 63.165 103.275 63.335 103.445 ;
      RECT 62.705 103.275 62.875 103.445 ;
      RECT 62.245 103.275 62.415 103.445 ;
      RECT 61.785 103.275 61.955 103.445 ;
      RECT 61.325 103.275 61.495 103.445 ;
      RECT 60.865 103.275 61.035 103.445 ;
      RECT 60.405 103.275 60.575 103.445 ;
      RECT 59.945 103.275 60.115 103.445 ;
      RECT 59.485 103.275 59.655 103.445 ;
      RECT 59.025 103.275 59.195 103.445 ;
      RECT 58.565 103.275 58.735 103.445 ;
      RECT 58.105 103.275 58.275 103.445 ;
      RECT 57.645 103.275 57.815 103.445 ;
      RECT 57.185 103.275 57.355 103.445 ;
      RECT 56.725 103.275 56.895 103.445 ;
      RECT 56.265 103.275 56.435 103.445 ;
      RECT 55.805 103.275 55.975 103.445 ;
      RECT 55.345 103.275 55.515 103.445 ;
      RECT 54.885 103.275 55.055 103.445 ;
      RECT 54.425 103.275 54.595 103.445 ;
      RECT 53.965 103.275 54.135 103.445 ;
      RECT 53.505 103.275 53.675 103.445 ;
      RECT 53.045 103.275 53.215 103.445 ;
      RECT 52.585 103.275 52.755 103.445 ;
      RECT 52.125 103.275 52.295 103.445 ;
      RECT 51.665 103.275 51.835 103.445 ;
      RECT 51.205 103.275 51.375 103.445 ;
      RECT 50.745 103.275 50.915 103.445 ;
      RECT 50.285 103.275 50.455 103.445 ;
      RECT 49.825 103.275 49.995 103.445 ;
      RECT 49.365 103.275 49.535 103.445 ;
      RECT 48.905 103.275 49.075 103.445 ;
      RECT 48.445 103.275 48.615 103.445 ;
      RECT 47.985 103.275 48.155 103.445 ;
      RECT 47.525 103.275 47.695 103.445 ;
      RECT 47.065 103.275 47.235 103.445 ;
      RECT 46.605 103.275 46.775 103.445 ;
      RECT 46.145 103.275 46.315 103.445 ;
      RECT 45.685 103.275 45.855 103.445 ;
      RECT 45.225 103.275 45.395 103.445 ;
      RECT 44.765 103.275 44.935 103.445 ;
      RECT 44.305 103.275 44.475 103.445 ;
      RECT 43.845 103.275 44.015 103.445 ;
      RECT 43.385 103.275 43.555 103.445 ;
      RECT 42.925 103.275 43.095 103.445 ;
      RECT 42.465 103.275 42.635 103.445 ;
      RECT 42.005 103.275 42.175 103.445 ;
      RECT 41.545 103.275 41.715 103.445 ;
      RECT 41.085 103.275 41.255 103.445 ;
      RECT 40.625 103.275 40.795 103.445 ;
      RECT 40.165 103.275 40.335 103.445 ;
      RECT 39.705 103.275 39.875 103.445 ;
      RECT 39.245 103.275 39.415 103.445 ;
      RECT 38.785 103.275 38.955 103.445 ;
      RECT 38.325 103.275 38.495 103.445 ;
      RECT 37.865 103.275 38.035 103.445 ;
      RECT 37.405 103.275 37.575 103.445 ;
      RECT 36.945 103.275 37.115 103.445 ;
      RECT 36.485 103.275 36.655 103.445 ;
      RECT 36.025 103.275 36.195 103.445 ;
      RECT 35.565 103.275 35.735 103.445 ;
      RECT 35.105 103.275 35.275 103.445 ;
      RECT 34.645 103.275 34.815 103.445 ;
      RECT 34.185 103.275 34.355 103.445 ;
      RECT 33.725 103.275 33.895 103.445 ;
      RECT 33.265 103.275 33.435 103.445 ;
      RECT 32.805 103.275 32.975 103.445 ;
      RECT 32.345 103.275 32.515 103.445 ;
      RECT 31.885 103.275 32.055 103.445 ;
      RECT 31.425 103.275 31.595 103.445 ;
      RECT 30.965 103.275 31.135 103.445 ;
      RECT 30.505 103.275 30.675 103.445 ;
      RECT 30.045 103.275 30.215 103.445 ;
      RECT 29.585 103.275 29.755 103.445 ;
      RECT 29.125 103.275 29.295 103.445 ;
      RECT 28.665 103.275 28.835 103.445 ;
      RECT 28.205 103.275 28.375 103.445 ;
      RECT 27.745 103.275 27.915 103.445 ;
      RECT 27.285 103.275 27.455 103.445 ;
      RECT 26.825 103.275 26.995 103.445 ;
      RECT 26.365 103.275 26.535 103.445 ;
      RECT 25.905 103.275 26.075 103.445 ;
      RECT 25.445 103.275 25.615 103.445 ;
      RECT 24.985 103.275 25.155 103.445 ;
      RECT 24.525 103.275 24.695 103.445 ;
      RECT 24.065 103.275 24.235 103.445 ;
      RECT 23.605 103.275 23.775 103.445 ;
      RECT 23.145 103.275 23.315 103.445 ;
      RECT 22.685 103.275 22.855 103.445 ;
      RECT 22.225 103.275 22.395 103.445 ;
      RECT 21.765 103.275 21.935 103.445 ;
      RECT 21.305 103.275 21.475 103.445 ;
      RECT 20.845 103.275 21.015 103.445 ;
      RECT 20.385 103.275 20.555 103.445 ;
      RECT 19.925 103.275 20.095 103.445 ;
      RECT 19.465 103.275 19.635 103.445 ;
      RECT 19.005 103.275 19.175 103.445 ;
      RECT 18.545 103.275 18.715 103.445 ;
      RECT 18.085 103.275 18.255 103.445 ;
      RECT 17.625 103.275 17.795 103.445 ;
      RECT 17.165 103.275 17.335 103.445 ;
      RECT 16.705 103.275 16.875 103.445 ;
      RECT 16.245 103.275 16.415 103.445 ;
      RECT 15.785 103.275 15.955 103.445 ;
      RECT 15.325 103.275 15.495 103.445 ;
      RECT 14.865 103.275 15.035 103.445 ;
      RECT 14.405 103.275 14.575 103.445 ;
      RECT 13.945 103.275 14.115 103.445 ;
      RECT 13.485 103.275 13.655 103.445 ;
      RECT 13.025 103.275 13.195 103.445 ;
      RECT 12.565 103.275 12.735 103.445 ;
      RECT 12.105 103.275 12.275 103.445 ;
      RECT 11.645 103.275 11.815 103.445 ;
      RECT 11.185 103.275 11.355 103.445 ;
      RECT 10.725 103.275 10.895 103.445 ;
      RECT 10.265 103.275 10.435 103.445 ;
      RECT 9.805 103.275 9.975 103.445 ;
      RECT 9.345 103.275 9.515 103.445 ;
      RECT 8.885 103.275 9.055 103.445 ;
      RECT 8.425 103.275 8.595 103.445 ;
      RECT 7.965 103.275 8.135 103.445 ;
      RECT 7.505 103.275 7.675 103.445 ;
      RECT 7.045 103.275 7.215 103.445 ;
      RECT 6.585 103.275 6.755 103.445 ;
      RECT 6.125 103.275 6.295 103.445 ;
      RECT 5.665 103.275 5.835 103.445 ;
      RECT 5.205 103.275 5.375 103.445 ;
      RECT 4.745 103.275 4.915 103.445 ;
      RECT 4.285 103.275 4.455 103.445 ;
      RECT 3.825 103.275 3.995 103.445 ;
      RECT 3.365 103.275 3.535 103.445 ;
      RECT 2.905 103.275 3.075 103.445 ;
      RECT 2.445 103.275 2.615 103.445 ;
      RECT 1.985 103.275 2.155 103.445 ;
      RECT 1.525 103.275 1.695 103.445 ;
      RECT 1.065 103.275 1.235 103.445 ;
      RECT 0.605 103.275 0.775 103.445 ;
      RECT 0.145 103.275 0.315 103.445 ;
      RECT 141.365 100.555 141.535 100.725 ;
      RECT 140.905 100.555 141.075 100.725 ;
      RECT 0.605 100.555 0.775 100.725 ;
      RECT 0.145 100.555 0.315 100.725 ;
      RECT 141.365 97.835 141.535 98.005 ;
      RECT 140.905 97.835 141.075 98.005 ;
      RECT 0.605 97.835 0.775 98.005 ;
      RECT 0.145 97.835 0.315 98.005 ;
      RECT 141.365 95.115 141.535 95.285 ;
      RECT 140.905 95.115 141.075 95.285 ;
      RECT 0.605 95.115 0.775 95.285 ;
      RECT 0.145 95.115 0.315 95.285 ;
      RECT 141.365 92.395 141.535 92.565 ;
      RECT 140.905 92.395 141.075 92.565 ;
      RECT 0.605 92.395 0.775 92.565 ;
      RECT 0.145 92.395 0.315 92.565 ;
      RECT 141.365 89.675 141.535 89.845 ;
      RECT 140.905 89.675 141.075 89.845 ;
      RECT 0.605 89.675 0.775 89.845 ;
      RECT 0.145 89.675 0.315 89.845 ;
      RECT 141.365 86.955 141.535 87.125 ;
      RECT 140.905 86.955 141.075 87.125 ;
      RECT 0.605 86.955 0.775 87.125 ;
      RECT 0.145 86.955 0.315 87.125 ;
      RECT 141.365 84.235 141.535 84.405 ;
      RECT 140.905 84.235 141.075 84.405 ;
      RECT 0.605 84.235 0.775 84.405 ;
      RECT 0.145 84.235 0.315 84.405 ;
      RECT 141.365 81.515 141.535 81.685 ;
      RECT 140.905 81.515 141.075 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 141.365 78.795 141.535 78.965 ;
      RECT 140.905 78.795 141.075 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 141.365 76.075 141.535 76.245 ;
      RECT 140.905 76.075 141.075 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 141.365 73.355 141.535 73.525 ;
      RECT 140.905 73.355 141.075 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 141.365 70.635 141.535 70.805 ;
      RECT 140.905 70.635 141.075 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 141.365 67.915 141.535 68.085 ;
      RECT 140.905 67.915 141.075 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 141.365 65.195 141.535 65.365 ;
      RECT 140.905 65.195 141.075 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 141.365 62.475 141.535 62.645 ;
      RECT 140.905 62.475 141.075 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 141.365 59.755 141.535 59.925 ;
      RECT 140.905 59.755 141.075 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 141.365 57.035 141.535 57.205 ;
      RECT 140.905 57.035 141.075 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 141.365 54.315 141.535 54.485 ;
      RECT 140.905 54.315 141.075 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 141.365 51.595 141.535 51.765 ;
      RECT 140.905 51.595 141.075 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 141.365 48.875 141.535 49.045 ;
      RECT 140.905 48.875 141.075 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 141.365 46.155 141.535 46.325 ;
      RECT 140.905 46.155 141.075 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 141.365 43.435 141.535 43.605 ;
      RECT 140.905 43.435 141.075 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 141.365 40.715 141.535 40.885 ;
      RECT 140.905 40.715 141.075 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 141.365 37.995 141.535 38.165 ;
      RECT 140.905 37.995 141.075 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 141.365 35.275 141.535 35.445 ;
      RECT 140.905 35.275 141.075 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 141.365 32.555 141.535 32.725 ;
      RECT 140.905 32.555 141.075 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 141.365 29.835 141.535 30.005 ;
      RECT 140.905 29.835 141.075 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 141.365 27.115 141.535 27.285 ;
      RECT 140.905 27.115 141.075 27.285 ;
      RECT 140.445 27.115 140.615 27.285 ;
      RECT 139.985 27.115 140.155 27.285 ;
      RECT 139.525 27.115 139.695 27.285 ;
      RECT 139.065 27.115 139.235 27.285 ;
      RECT 138.605 27.115 138.775 27.285 ;
      RECT 138.145 27.115 138.315 27.285 ;
      RECT 137.685 27.115 137.855 27.285 ;
      RECT 137.225 27.115 137.395 27.285 ;
      RECT 136.765 27.115 136.935 27.285 ;
      RECT 136.305 27.115 136.475 27.285 ;
      RECT 135.845 27.115 136.015 27.285 ;
      RECT 135.385 27.115 135.555 27.285 ;
      RECT 134.925 27.115 135.095 27.285 ;
      RECT 134.465 27.115 134.635 27.285 ;
      RECT 134.005 27.115 134.175 27.285 ;
      RECT 133.545 27.115 133.715 27.285 ;
      RECT 133.085 27.115 133.255 27.285 ;
      RECT 132.625 27.115 132.795 27.285 ;
      RECT 132.165 27.115 132.335 27.285 ;
      RECT 131.705 27.115 131.875 27.285 ;
      RECT 131.245 27.115 131.415 27.285 ;
      RECT 130.785 27.115 130.955 27.285 ;
      RECT 130.325 27.115 130.495 27.285 ;
      RECT 129.865 27.115 130.035 27.285 ;
      RECT 129.405 27.115 129.575 27.285 ;
      RECT 128.945 27.115 129.115 27.285 ;
      RECT 128.485 27.115 128.655 27.285 ;
      RECT 128.025 27.115 128.195 27.285 ;
      RECT 127.565 27.115 127.735 27.285 ;
      RECT 127.105 27.115 127.275 27.285 ;
      RECT 126.645 27.115 126.815 27.285 ;
      RECT 126.185 27.115 126.355 27.285 ;
      RECT 125.725 27.115 125.895 27.285 ;
      RECT 125.265 27.115 125.435 27.285 ;
      RECT 124.805 27.115 124.975 27.285 ;
      RECT 124.345 27.115 124.515 27.285 ;
      RECT 123.885 27.115 124.055 27.285 ;
      RECT 123.425 27.115 123.595 27.285 ;
      RECT 122.965 27.115 123.135 27.285 ;
      RECT 122.505 27.115 122.675 27.285 ;
      RECT 122.045 27.115 122.215 27.285 ;
      RECT 121.585 27.115 121.755 27.285 ;
      RECT 121.125 27.115 121.295 27.285 ;
      RECT 120.665 27.115 120.835 27.285 ;
      RECT 120.205 27.115 120.375 27.285 ;
      RECT 119.745 27.115 119.915 27.285 ;
      RECT 119.285 27.115 119.455 27.285 ;
      RECT 118.825 27.115 118.995 27.285 ;
      RECT 118.365 27.115 118.535 27.285 ;
      RECT 117.905 27.115 118.075 27.285 ;
      RECT 117.445 27.115 117.615 27.285 ;
      RECT 116.985 27.115 117.155 27.285 ;
      RECT 116.525 27.115 116.695 27.285 ;
      RECT 116.065 27.115 116.235 27.285 ;
      RECT 115.605 27.115 115.775 27.285 ;
      RECT 115.145 27.115 115.315 27.285 ;
      RECT 114.685 27.115 114.855 27.285 ;
      RECT 114.225 27.115 114.395 27.285 ;
      RECT 113.765 27.115 113.935 27.285 ;
      RECT 113.305 27.115 113.475 27.285 ;
      RECT 112.845 27.115 113.015 27.285 ;
      RECT 112.385 27.115 112.555 27.285 ;
      RECT 111.925 27.115 112.095 27.285 ;
      RECT 111.465 27.115 111.635 27.285 ;
      RECT 111.005 27.115 111.175 27.285 ;
      RECT 110.545 27.115 110.715 27.285 ;
      RECT 110.085 27.115 110.255 27.285 ;
      RECT 109.625 27.115 109.795 27.285 ;
      RECT 109.165 27.115 109.335 27.285 ;
      RECT 108.705 27.115 108.875 27.285 ;
      RECT 108.245 27.115 108.415 27.285 ;
      RECT 107.785 27.115 107.955 27.285 ;
      RECT 107.325 27.115 107.495 27.285 ;
      RECT 106.865 27.115 107.035 27.285 ;
      RECT 106.405 27.115 106.575 27.285 ;
      RECT 105.945 27.115 106.115 27.285 ;
      RECT 105.485 27.115 105.655 27.285 ;
      RECT 105.025 27.115 105.195 27.285 ;
      RECT 104.565 27.115 104.735 27.285 ;
      RECT 104.105 27.115 104.275 27.285 ;
      RECT 103.645 27.115 103.815 27.285 ;
      RECT 103.185 27.115 103.355 27.285 ;
      RECT 102.725 27.115 102.895 27.285 ;
      RECT 102.265 27.115 102.435 27.285 ;
      RECT 101.805 27.115 101.975 27.285 ;
      RECT 101.345 27.115 101.515 27.285 ;
      RECT 100.885 27.115 101.055 27.285 ;
      RECT 100.425 27.115 100.595 27.285 ;
      RECT 99.965 27.115 100.135 27.285 ;
      RECT 99.505 27.115 99.675 27.285 ;
      RECT 99.045 27.115 99.215 27.285 ;
      RECT 98.585 27.115 98.755 27.285 ;
      RECT 98.125 27.115 98.295 27.285 ;
      RECT 97.665 27.115 97.835 27.285 ;
      RECT 97.205 27.115 97.375 27.285 ;
      RECT 96.745 27.115 96.915 27.285 ;
      RECT 96.285 27.115 96.455 27.285 ;
      RECT 95.825 27.115 95.995 27.285 ;
      RECT 95.365 27.115 95.535 27.285 ;
      RECT 94.905 27.115 95.075 27.285 ;
      RECT 94.445 27.115 94.615 27.285 ;
      RECT 93.985 27.115 94.155 27.285 ;
      RECT 93.525 27.115 93.695 27.285 ;
      RECT 93.065 27.115 93.235 27.285 ;
      RECT 92.605 27.115 92.775 27.285 ;
      RECT 92.145 27.115 92.315 27.285 ;
      RECT 91.685 27.115 91.855 27.285 ;
      RECT 91.225 27.115 91.395 27.285 ;
      RECT 90.765 27.115 90.935 27.285 ;
      RECT 90.305 27.115 90.475 27.285 ;
      RECT 89.845 27.115 90.015 27.285 ;
      RECT 89.385 27.115 89.555 27.285 ;
      RECT 88.925 27.115 89.095 27.285 ;
      RECT 88.465 27.115 88.635 27.285 ;
      RECT 88.005 27.115 88.175 27.285 ;
      RECT 87.545 27.115 87.715 27.285 ;
      RECT 87.085 27.115 87.255 27.285 ;
      RECT 86.625 27.115 86.795 27.285 ;
      RECT 86.165 27.115 86.335 27.285 ;
      RECT 85.705 27.115 85.875 27.285 ;
      RECT 85.245 27.115 85.415 27.285 ;
      RECT 84.785 27.115 84.955 27.285 ;
      RECT 84.325 27.115 84.495 27.285 ;
      RECT 83.865 27.115 84.035 27.285 ;
      RECT 83.405 27.115 83.575 27.285 ;
      RECT 82.945 27.115 83.115 27.285 ;
      RECT 82.485 27.115 82.655 27.285 ;
      RECT 82.025 27.115 82.195 27.285 ;
      RECT 81.565 27.115 81.735 27.285 ;
      RECT 81.105 27.115 81.275 27.285 ;
      RECT 80.645 27.115 80.815 27.285 ;
      RECT 80.185 27.115 80.355 27.285 ;
      RECT 79.725 27.115 79.895 27.285 ;
      RECT 79.265 27.115 79.435 27.285 ;
      RECT 78.805 27.115 78.975 27.285 ;
      RECT 78.345 27.115 78.515 27.285 ;
      RECT 77.885 27.115 78.055 27.285 ;
      RECT 77.425 27.115 77.595 27.285 ;
      RECT 76.965 27.115 77.135 27.285 ;
      RECT 76.505 27.115 76.675 27.285 ;
      RECT 76.045 27.115 76.215 27.285 ;
      RECT 75.585 27.115 75.755 27.285 ;
      RECT 75.125 27.115 75.295 27.285 ;
      RECT 74.665 27.115 74.835 27.285 ;
      RECT 74.205 27.115 74.375 27.285 ;
      RECT 73.745 27.115 73.915 27.285 ;
      RECT 73.285 27.115 73.455 27.285 ;
      RECT 72.825 27.115 72.995 27.285 ;
      RECT 72.365 27.115 72.535 27.285 ;
      RECT 71.905 27.115 72.075 27.285 ;
      RECT 71.445 27.115 71.615 27.285 ;
      RECT 70.985 27.115 71.155 27.285 ;
      RECT 70.525 27.115 70.695 27.285 ;
      RECT 70.065 27.115 70.235 27.285 ;
      RECT 69.605 27.115 69.775 27.285 ;
      RECT 69.145 27.115 69.315 27.285 ;
      RECT 68.685 27.115 68.855 27.285 ;
      RECT 68.225 27.115 68.395 27.285 ;
      RECT 67.765 27.115 67.935 27.285 ;
      RECT 67.305 27.115 67.475 27.285 ;
      RECT 66.845 27.115 67.015 27.285 ;
      RECT 66.385 27.115 66.555 27.285 ;
      RECT 65.925 27.115 66.095 27.285 ;
      RECT 65.465 27.115 65.635 27.285 ;
      RECT 65.005 27.115 65.175 27.285 ;
      RECT 64.545 27.115 64.715 27.285 ;
      RECT 64.085 27.115 64.255 27.285 ;
      RECT 63.625 27.115 63.795 27.285 ;
      RECT 63.165 27.115 63.335 27.285 ;
      RECT 62.705 27.115 62.875 27.285 ;
      RECT 62.245 27.115 62.415 27.285 ;
      RECT 61.785 27.115 61.955 27.285 ;
      RECT 61.325 27.115 61.495 27.285 ;
      RECT 60.865 27.115 61.035 27.285 ;
      RECT 60.405 27.115 60.575 27.285 ;
      RECT 59.945 27.115 60.115 27.285 ;
      RECT 59.485 27.115 59.655 27.285 ;
      RECT 59.025 27.115 59.195 27.285 ;
      RECT 58.565 27.115 58.735 27.285 ;
      RECT 58.105 27.115 58.275 27.285 ;
      RECT 57.645 27.115 57.815 27.285 ;
      RECT 57.185 27.115 57.355 27.285 ;
      RECT 56.725 27.115 56.895 27.285 ;
      RECT 56.265 27.115 56.435 27.285 ;
      RECT 55.805 27.115 55.975 27.285 ;
      RECT 55.345 27.115 55.515 27.285 ;
      RECT 54.885 27.115 55.055 27.285 ;
      RECT 54.425 27.115 54.595 27.285 ;
      RECT 53.965 27.115 54.135 27.285 ;
      RECT 53.505 27.115 53.675 27.285 ;
      RECT 53.045 27.115 53.215 27.285 ;
      RECT 52.585 27.115 52.755 27.285 ;
      RECT 52.125 27.115 52.295 27.285 ;
      RECT 51.665 27.115 51.835 27.285 ;
      RECT 51.205 27.115 51.375 27.285 ;
      RECT 50.745 27.115 50.915 27.285 ;
      RECT 50.285 27.115 50.455 27.285 ;
      RECT 49.825 27.115 49.995 27.285 ;
      RECT 49.365 27.115 49.535 27.285 ;
      RECT 48.905 27.115 49.075 27.285 ;
      RECT 48.445 27.115 48.615 27.285 ;
      RECT 47.985 27.115 48.155 27.285 ;
      RECT 47.525 27.115 47.695 27.285 ;
      RECT 47.065 27.115 47.235 27.285 ;
      RECT 46.605 27.115 46.775 27.285 ;
      RECT 46.145 27.115 46.315 27.285 ;
      RECT 45.685 27.115 45.855 27.285 ;
      RECT 45.225 27.115 45.395 27.285 ;
      RECT 44.765 27.115 44.935 27.285 ;
      RECT 44.305 27.115 44.475 27.285 ;
      RECT 43.845 27.115 44.015 27.285 ;
      RECT 43.385 27.115 43.555 27.285 ;
      RECT 42.925 27.115 43.095 27.285 ;
      RECT 42.465 27.115 42.635 27.285 ;
      RECT 42.005 27.115 42.175 27.285 ;
      RECT 41.545 27.115 41.715 27.285 ;
      RECT 41.085 27.115 41.255 27.285 ;
      RECT 40.625 27.115 40.795 27.285 ;
      RECT 40.165 27.115 40.335 27.285 ;
      RECT 39.705 27.115 39.875 27.285 ;
      RECT 39.245 27.115 39.415 27.285 ;
      RECT 38.785 27.115 38.955 27.285 ;
      RECT 38.325 27.115 38.495 27.285 ;
      RECT 37.865 27.115 38.035 27.285 ;
      RECT 37.405 27.115 37.575 27.285 ;
      RECT 36.945 27.115 37.115 27.285 ;
      RECT 36.485 27.115 36.655 27.285 ;
      RECT 36.025 27.115 36.195 27.285 ;
      RECT 35.565 27.115 35.735 27.285 ;
      RECT 35.105 27.115 35.275 27.285 ;
      RECT 34.645 27.115 34.815 27.285 ;
      RECT 34.185 27.115 34.355 27.285 ;
      RECT 33.725 27.115 33.895 27.285 ;
      RECT 33.265 27.115 33.435 27.285 ;
      RECT 32.805 27.115 32.975 27.285 ;
      RECT 32.345 27.115 32.515 27.285 ;
      RECT 31.885 27.115 32.055 27.285 ;
      RECT 31.425 27.115 31.595 27.285 ;
      RECT 30.965 27.115 31.135 27.285 ;
      RECT 30.505 27.115 30.675 27.285 ;
      RECT 30.045 27.115 30.215 27.285 ;
      RECT 29.585 27.115 29.755 27.285 ;
      RECT 29.125 27.115 29.295 27.285 ;
      RECT 28.665 27.115 28.835 27.285 ;
      RECT 28.205 27.115 28.375 27.285 ;
      RECT 27.745 27.115 27.915 27.285 ;
      RECT 27.285 27.115 27.455 27.285 ;
      RECT 26.825 27.115 26.995 27.285 ;
      RECT 26.365 27.115 26.535 27.285 ;
      RECT 25.905 27.115 26.075 27.285 ;
      RECT 25.445 27.115 25.615 27.285 ;
      RECT 24.985 27.115 25.155 27.285 ;
      RECT 24.525 27.115 24.695 27.285 ;
      RECT 24.065 27.115 24.235 27.285 ;
      RECT 23.605 27.115 23.775 27.285 ;
      RECT 23.145 27.115 23.315 27.285 ;
      RECT 22.685 27.115 22.855 27.285 ;
      RECT 22.225 27.115 22.395 27.285 ;
      RECT 21.765 27.115 21.935 27.285 ;
      RECT 21.305 27.115 21.475 27.285 ;
      RECT 20.845 27.115 21.015 27.285 ;
      RECT 20.385 27.115 20.555 27.285 ;
      RECT 19.925 27.115 20.095 27.285 ;
      RECT 19.465 27.115 19.635 27.285 ;
      RECT 19.005 27.115 19.175 27.285 ;
      RECT 18.545 27.115 18.715 27.285 ;
      RECT 18.085 27.115 18.255 27.285 ;
      RECT 17.625 27.115 17.795 27.285 ;
      RECT 17.165 27.115 17.335 27.285 ;
      RECT 16.705 27.115 16.875 27.285 ;
      RECT 16.245 27.115 16.415 27.285 ;
      RECT 15.785 27.115 15.955 27.285 ;
      RECT 15.325 27.115 15.495 27.285 ;
      RECT 14.865 27.115 15.035 27.285 ;
      RECT 14.405 27.115 14.575 27.285 ;
      RECT 13.945 27.115 14.115 27.285 ;
      RECT 13.485 27.115 13.655 27.285 ;
      RECT 13.025 27.115 13.195 27.285 ;
      RECT 12.565 27.115 12.735 27.285 ;
      RECT 12.105 27.115 12.275 27.285 ;
      RECT 11.645 27.115 11.815 27.285 ;
      RECT 11.185 27.115 11.355 27.285 ;
      RECT 10.725 27.115 10.895 27.285 ;
      RECT 10.265 27.115 10.435 27.285 ;
      RECT 9.805 27.115 9.975 27.285 ;
      RECT 9.345 27.115 9.515 27.285 ;
      RECT 8.885 27.115 9.055 27.285 ;
      RECT 8.425 27.115 8.595 27.285 ;
      RECT 7.965 27.115 8.135 27.285 ;
      RECT 7.505 27.115 7.675 27.285 ;
      RECT 7.045 27.115 7.215 27.285 ;
      RECT 6.585 27.115 6.755 27.285 ;
      RECT 6.125 27.115 6.295 27.285 ;
      RECT 5.665 27.115 5.835 27.285 ;
      RECT 5.205 27.115 5.375 27.285 ;
      RECT 4.745 27.115 4.915 27.285 ;
      RECT 4.285 27.115 4.455 27.285 ;
      RECT 3.825 27.115 3.995 27.285 ;
      RECT 3.365 27.115 3.535 27.285 ;
      RECT 2.905 27.115 3.075 27.285 ;
      RECT 2.445 27.115 2.615 27.285 ;
      RECT 1.985 27.115 2.155 27.285 ;
      RECT 1.525 27.115 1.695 27.285 ;
      RECT 1.065 27.115 1.235 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 112.845 24.395 113.015 24.565 ;
      RECT 112.385 24.395 112.555 24.565 ;
      RECT 29.125 24.395 29.295 24.565 ;
      RECT 28.665 24.395 28.835 24.565 ;
      RECT 112.845 21.675 113.015 21.845 ;
      RECT 112.385 21.675 112.555 21.845 ;
      RECT 29.125 21.675 29.295 21.845 ;
      RECT 28.665 21.675 28.835 21.845 ;
      RECT 112.845 18.955 113.015 19.125 ;
      RECT 112.385 18.955 112.555 19.125 ;
      RECT 29.125 18.955 29.295 19.125 ;
      RECT 28.665 18.955 28.835 19.125 ;
      RECT 112.845 16.235 113.015 16.405 ;
      RECT 112.385 16.235 112.555 16.405 ;
      RECT 29.125 16.235 29.295 16.405 ;
      RECT 28.665 16.235 28.835 16.405 ;
      RECT 112.845 13.515 113.015 13.685 ;
      RECT 112.385 13.515 112.555 13.685 ;
      RECT 29.125 13.515 29.295 13.685 ;
      RECT 28.665 13.515 28.835 13.685 ;
      RECT 112.845 10.795 113.015 10.965 ;
      RECT 112.385 10.795 112.555 10.965 ;
      RECT 29.125 10.795 29.295 10.965 ;
      RECT 28.665 10.795 28.835 10.965 ;
      RECT 112.845 8.075 113.015 8.245 ;
      RECT 112.385 8.075 112.555 8.245 ;
      RECT 29.125 8.075 29.295 8.245 ;
      RECT 28.665 8.075 28.835 8.245 ;
      RECT 112.845 5.355 113.015 5.525 ;
      RECT 112.385 5.355 112.555 5.525 ;
      RECT 29.125 5.355 29.295 5.525 ;
      RECT 28.665 5.355 28.835 5.525 ;
      RECT 112.845 2.635 113.015 2.805 ;
      RECT 112.385 2.635 112.555 2.805 ;
      RECT 29.125 2.635 29.295 2.805 ;
      RECT 28.665 2.635 28.835 2.805 ;
      RECT 112.845 -0.085 113.015 0.085 ;
      RECT 112.385 -0.085 112.555 0.085 ;
      RECT 111.925 -0.085 112.095 0.085 ;
      RECT 111.465 -0.085 111.635 0.085 ;
      RECT 111.005 -0.085 111.175 0.085 ;
      RECT 110.545 -0.085 110.715 0.085 ;
      RECT 110.085 -0.085 110.255 0.085 ;
      RECT 109.625 -0.085 109.795 0.085 ;
      RECT 109.165 -0.085 109.335 0.085 ;
      RECT 108.705 -0.085 108.875 0.085 ;
      RECT 108.245 -0.085 108.415 0.085 ;
      RECT 107.785 -0.085 107.955 0.085 ;
      RECT 107.325 -0.085 107.495 0.085 ;
      RECT 106.865 -0.085 107.035 0.085 ;
      RECT 106.405 -0.085 106.575 0.085 ;
      RECT 105.945 -0.085 106.115 0.085 ;
      RECT 105.485 -0.085 105.655 0.085 ;
      RECT 105.025 -0.085 105.195 0.085 ;
      RECT 104.565 -0.085 104.735 0.085 ;
      RECT 104.105 -0.085 104.275 0.085 ;
      RECT 103.645 -0.085 103.815 0.085 ;
      RECT 103.185 -0.085 103.355 0.085 ;
      RECT 102.725 -0.085 102.895 0.085 ;
      RECT 102.265 -0.085 102.435 0.085 ;
      RECT 101.805 -0.085 101.975 0.085 ;
      RECT 101.345 -0.085 101.515 0.085 ;
      RECT 100.885 -0.085 101.055 0.085 ;
      RECT 100.425 -0.085 100.595 0.085 ;
      RECT 99.965 -0.085 100.135 0.085 ;
      RECT 99.505 -0.085 99.675 0.085 ;
      RECT 99.045 -0.085 99.215 0.085 ;
      RECT 98.585 -0.085 98.755 0.085 ;
      RECT 98.125 -0.085 98.295 0.085 ;
      RECT 97.665 -0.085 97.835 0.085 ;
      RECT 97.205 -0.085 97.375 0.085 ;
      RECT 96.745 -0.085 96.915 0.085 ;
      RECT 96.285 -0.085 96.455 0.085 ;
      RECT 95.825 -0.085 95.995 0.085 ;
      RECT 95.365 -0.085 95.535 0.085 ;
      RECT 94.905 -0.085 95.075 0.085 ;
      RECT 94.445 -0.085 94.615 0.085 ;
      RECT 93.985 -0.085 94.155 0.085 ;
      RECT 93.525 -0.085 93.695 0.085 ;
      RECT 93.065 -0.085 93.235 0.085 ;
      RECT 92.605 -0.085 92.775 0.085 ;
      RECT 92.145 -0.085 92.315 0.085 ;
      RECT 91.685 -0.085 91.855 0.085 ;
      RECT 91.225 -0.085 91.395 0.085 ;
      RECT 90.765 -0.085 90.935 0.085 ;
      RECT 90.305 -0.085 90.475 0.085 ;
      RECT 89.845 -0.085 90.015 0.085 ;
      RECT 89.385 -0.085 89.555 0.085 ;
      RECT 88.925 -0.085 89.095 0.085 ;
      RECT 88.465 -0.085 88.635 0.085 ;
      RECT 88.005 -0.085 88.175 0.085 ;
      RECT 87.545 -0.085 87.715 0.085 ;
      RECT 87.085 -0.085 87.255 0.085 ;
      RECT 86.625 -0.085 86.795 0.085 ;
      RECT 86.165 -0.085 86.335 0.085 ;
      RECT 85.705 -0.085 85.875 0.085 ;
      RECT 85.245 -0.085 85.415 0.085 ;
      RECT 84.785 -0.085 84.955 0.085 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
    LAYER via ;
      RECT 85.485 130.485 85.635 130.635 ;
      RECT 56.045 130.485 56.195 130.635 ;
      RECT 62.025 128.785 62.175 128.935 ;
      RECT 85.485 103.285 85.635 103.435 ;
      RECT 56.045 103.285 56.195 103.435 ;
      RECT 6.365 103.285 6.515 103.435 ;
      RECT 139.305 101.585 139.455 101.735 ;
      RECT 4.985 101.585 5.135 101.735 ;
      RECT 4.065 101.585 4.215 101.735 ;
      RECT 85.485 27.125 85.635 27.275 ;
      RECT 56.045 27.125 56.195 27.275 ;
      RECT 6.365 27.125 6.515 27.275 ;
      RECT 80.425 1.625 80.575 1.775 ;
      RECT 85.485 -0.075 85.635 0.075 ;
      RECT 56.045 -0.075 56.195 0.075 ;
    LAYER via2 ;
      RECT 85.46 130.46 85.66 130.66 ;
      RECT 56.02 130.46 56.22 130.66 ;
      RECT 29.8 125.02 30 125.22 ;
      RECT 29.8 118.9 30 119.1 ;
      RECT 111.68 117.54 111.88 117.74 ;
      RECT 6.34 103.26 6.54 103.46 ;
      RECT 1.28 99.18 1.48 99.38 ;
      RECT 1.28 91.02 1.48 91.22 ;
      RECT 1.74 64.5 1.94 64.7 ;
      RECT 139.74 63.82 139.94 64.02 ;
      RECT 1.74 52.94 1.94 53.14 ;
      RECT 140.2 48.86 140.4 49.06 ;
      RECT 1.74 47.5 1.94 47.7 ;
      RECT 6.34 27.1 6.54 27.3 ;
      RECT 29.8 3.3 30 3.5 ;
      RECT 85.46 -0.1 85.66 0.1 ;
      RECT 56.02 -0.1 56.22 0.1 ;
    LAYER via3 ;
      RECT 85.46 130.46 85.66 130.66 ;
      RECT 56.02 130.46 56.22 130.66 ;
      RECT 6.34 103.26 6.54 103.46 ;
      RECT 1.74 65.86 1.94 66.06 ;
      RECT 1.74 54.3 1.94 54.5 ;
      RECT 6.34 27.1 6.54 27.3 ;
      RECT 85.46 -0.1 85.66 0.1 ;
      RECT 56.02 -0.1 56.22 0.1 ;
    LAYER via4 ;
      RECT 134.84 86.08 135.64 86.88 ;
      RECT 134.84 84.48 135.64 85.28 ;
      RECT 6.04 65.68 6.84 66.48 ;
      RECT 6.04 64.08 6.84 64.88 ;
      RECT 134.84 45.28 135.64 46.08 ;
      RECT 134.84 43.68 135.64 44.48 ;
    LAYER fieldpoly ;
      POLYGON 113.02 130.42 113.02 103.22 141.54 103.22 141.54 27.34 113.02 27.34 113.02 0.14 28.66 0.14 28.66 27.34 0.14 27.34 0.14 103.22 28.66 103.22 28.66 130.42 ;
    LAYER diff ;
      POLYGON 113.16 130.56 113.16 103.36 141.68 103.36 141.68 27.2 113.16 27.2 113.16 0 28.52 0 28.52 27.2 0 27.2 0 103.36 28.52 103.36 28.52 130.56 ;
    LAYER nwell ;
      POLYGON 113.35 129.255 113.35 126.425 112.51 126.425 112.51 127.65 109.29 127.65 109.29 129.255 ;
      RECT 28.33 126.425 32.39 129.255 ;
      POLYGON 113.35 123.815 113.35 120.985 112.51 120.985 112.51 122.21 112.05 122.21 112.05 123.815 ;
      POLYGON 30.55 123.815 30.55 122.59 32.39 122.59 32.39 120.985 28.33 120.985 28.33 123.815 ;
      POLYGON 113.35 118.375 113.35 115.545 112.51 115.545 112.51 116.77 112.05 116.77 112.05 118.375 ;
      POLYGON 32.39 118.375 32.39 116.77 30.55 116.77 30.55 115.545 28.33 115.545 28.33 118.375 ;
      POLYGON 113.35 112.935 113.35 110.105 112.05 110.105 112.05 111.71 112.51 111.71 112.51 112.935 ;
      POLYGON 30.55 112.935 30.55 111.71 32.39 111.71 32.39 110.105 28.33 110.105 28.33 112.935 ;
      RECT 112.05 104.665 113.35 107.495 ;
      POLYGON 32.39 107.495 32.39 105.89 30.55 105.89 30.55 104.665 28.33 104.665 28.33 107.495 ;
      POLYGON 141.87 102.055 141.87 99.225 141.03 99.225 141.03 100.45 139.65 100.45 139.65 102.055 ;
      POLYGON 3.87 102.055 3.87 100.45 2.03 100.45 2.03 99.225 -0.19 99.225 -0.19 102.055 ;
      POLYGON 141.87 96.615 141.87 93.785 140.57 93.785 140.57 95.39 141.03 95.39 141.03 96.615 ;
      POLYGON 2.03 96.615 2.03 95.39 3.87 95.39 3.87 93.785 -0.19 93.785 -0.19 96.615 ;
      POLYGON 141.87 91.175 141.87 88.345 141.03 88.345 141.03 89.57 140.57 89.57 140.57 91.175 ;
      RECT -0.19 88.345 2.03 91.175 ;
      RECT 140.57 82.905 141.87 85.735 ;
      RECT -0.19 82.905 2.03 85.735 ;
      RECT 140.57 77.465 141.87 80.295 ;
      RECT -0.19 77.465 2.03 80.295 ;
      RECT 140.57 72.025 141.87 74.855 ;
      RECT -0.19 72.025 2.03 74.855 ;
      RECT 140.57 66.585 141.87 69.415 ;
      RECT -0.19 66.585 2.03 69.415 ;
      RECT 140.57 61.145 141.87 63.975 ;
      POLYGON 2.03 63.975 2.03 62.75 3.87 62.75 3.87 61.145 -0.19 61.145 -0.19 63.975 ;
      RECT 140.57 55.705 141.87 58.535 ;
      RECT -0.19 55.705 2.03 58.535 ;
      RECT 140.57 50.265 141.87 53.095 ;
      RECT -0.19 50.265 2.03 53.095 ;
      RECT 140.57 44.825 141.87 47.655 ;
      RECT -0.19 44.825 2.03 47.655 ;
      RECT 141.03 39.385 141.87 42.215 ;
      RECT -0.19 39.385 2.03 42.215 ;
      RECT 140.57 33.945 141.87 36.775 ;
      RECT -0.19 33.945 3.87 36.775 ;
      RECT 141.03 28.505 141.87 31.335 ;
      RECT -0.19 28.505 3.87 31.335 ;
      RECT 112.51 23.065 113.35 25.895 ;
      RECT 28.33 23.065 32.39 25.895 ;
      POLYGON 113.35 20.455 113.35 17.625 112.51 17.625 112.51 18.85 112.05 18.85 112.05 20.455 ;
      RECT 28.33 17.625 32.39 20.455 ;
      POLYGON 113.35 15.015 113.35 12.185 112.51 12.185 112.51 13.41 109.29 13.41 109.29 15.015 ;
      POLYGON 30.55 15.015 30.55 13.79 32.39 13.79 32.39 12.185 28.33 12.185 28.33 15.015 ;
      POLYGON 113.35 9.575 113.35 6.745 112.05 6.745 112.05 7.97 109.29 7.97 109.29 9.575 ;
      RECT 28.33 6.745 32.39 9.575 ;
      POLYGON 113.35 4.135 113.35 1.305 109.29 1.305 109.29 2.91 112.51 2.91 112.51 4.135 ;
      RECT 28.33 1.305 32.39 4.135 ;
      POLYGON 113.16 130.56 113.16 103.36 141.68 103.36 141.68 27.2 113.16 27.2 113.16 0 28.52 0 28.52 27.2 0 27.2 0 103.36 28.52 103.36 28.52 130.56 ;
    LAYER pwell ;
      RECT 109.61 130.51 109.83 130.68 ;
      RECT 105.93 130.51 106.15 130.68 ;
      RECT 102.25 130.51 102.47 130.68 ;
      RECT 98.57 130.51 98.79 130.68 ;
      RECT 94.89 130.51 95.11 130.68 ;
      RECT 91.21 130.51 91.43 130.68 ;
      RECT 87.53 130.51 87.75 130.68 ;
      RECT 83.85 130.51 84.07 130.68 ;
      RECT 80.17 130.51 80.39 130.68 ;
      RECT 76.49 130.51 76.71 130.68 ;
      RECT 72.81 130.51 73.03 130.68 ;
      RECT 69.13 130.51 69.35 130.68 ;
      RECT 65.45 130.51 65.67 130.68 ;
      RECT 61.77 130.51 61.99 130.68 ;
      RECT 58.09 130.51 58.31 130.68 ;
      RECT 54.41 130.51 54.63 130.68 ;
      RECT 50.73 130.51 50.95 130.68 ;
      RECT 47.05 130.51 47.27 130.68 ;
      RECT 43.37 130.51 43.59 130.68 ;
      RECT 39.69 130.51 39.91 130.68 ;
      RECT 36.01 130.51 36.23 130.68 ;
      RECT 32.33 130.51 32.55 130.68 ;
      RECT 28.65 130.51 28.87 130.68 ;
      RECT 136.29 103.31 136.51 103.48 ;
      RECT 132.61 103.31 132.83 103.48 ;
      RECT 128.93 103.31 129.15 103.48 ;
      RECT 125.25 103.31 125.47 103.48 ;
      RECT 121.57 103.31 121.79 103.48 ;
      RECT 117.89 103.31 118.11 103.48 ;
      RECT 114.21 103.31 114.43 103.48 ;
      RECT 25.89 103.31 26.11 103.48 ;
      RECT 22.21 103.31 22.43 103.48 ;
      RECT 18.53 103.31 18.75 103.48 ;
      RECT 14.85 103.31 15.07 103.48 ;
      RECT 11.17 103.31 11.39 103.48 ;
      RECT 7.49 103.31 7.71 103.48 ;
      RECT 3.81 103.31 4.03 103.48 ;
      RECT 0.13 103.31 0.35 103.48 ;
      RECT 140.015 103.3 140.125 103.42 ;
      RECT 140.455 27.15 140.615 27.26 ;
      RECT 141.36 27.145 141.48 27.255 ;
      RECT 136.75 27.08 136.97 27.25 ;
      RECT 133.07 27.08 133.29 27.25 ;
      RECT 129.39 27.08 129.61 27.25 ;
      RECT 125.71 27.08 125.93 27.25 ;
      RECT 122.03 27.08 122.25 27.25 ;
      RECT 118.35 27.08 118.57 27.25 ;
      RECT 114.67 27.08 114.89 27.25 ;
      RECT 25.89 27.08 26.11 27.25 ;
      RECT 22.21 27.08 22.43 27.25 ;
      RECT 18.53 27.08 18.75 27.25 ;
      RECT 14.85 27.08 15.07 27.25 ;
      RECT 11.17 27.08 11.39 27.25 ;
      RECT 7.49 27.08 7.71 27.25 ;
      RECT 3.81 27.08 4.03 27.25 ;
      RECT 0.13 27.08 0.35 27.25 ;
      RECT 109.61 -0.12 109.83 0.05 ;
      RECT 105.93 -0.12 106.15 0.05 ;
      RECT 102.25 -0.12 102.47 0.05 ;
      RECT 98.57 -0.12 98.79 0.05 ;
      RECT 94.89 -0.12 95.11 0.05 ;
      RECT 91.21 -0.12 91.43 0.05 ;
      RECT 87.53 -0.12 87.75 0.05 ;
      RECT 83.85 -0.12 84.07 0.05 ;
      RECT 80.17 -0.12 80.39 0.05 ;
      RECT 76.49 -0.12 76.71 0.05 ;
      RECT 72.81 -0.12 73.03 0.05 ;
      RECT 69.13 -0.12 69.35 0.05 ;
      RECT 65.45 -0.12 65.67 0.05 ;
      RECT 61.77 -0.12 61.99 0.05 ;
      RECT 58.09 -0.12 58.31 0.05 ;
      RECT 54.41 -0.12 54.63 0.05 ;
      RECT 50.73 -0.12 50.95 0.05 ;
      RECT 47.05 -0.12 47.27 0.05 ;
      RECT 43.37 -0.12 43.59 0.05 ;
      RECT 39.69 -0.12 39.91 0.05 ;
      RECT 36.01 -0.12 36.23 0.05 ;
      RECT 32.33 -0.12 32.55 0.05 ;
      RECT 28.65 -0.12 28.87 0.05 ;
      POLYGON 113.16 130.56 113.16 103.36 141.68 103.36 141.68 27.2 113.16 27.2 113.16 0 28.52 0 28.52 27.2 0 27.2 0 103.36 28.52 103.36 28.52 130.56 ;
    LAYER OVERLAP ;
      POLYGON 28.52 0 28.52 27.2 0 27.2 0 103.36 28.52 103.36 28.52 130.56 113.16 130.56 113.16 103.36 141.68 103.36 141.68 27.2 113.16 27.2 113.16 0 ;
  END
END sb_1__1_

END LIBRARY
