VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_0__0_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 103.96 BY 125.12 ;
  SYMMETRY X Y ;
  PIN pReset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 63.34 0.595 63.48 ;
    END
  END pReset[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 19.63 124.32 19.93 125.12 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.7 124.635 68.84 125.12 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.36 124.635 55.5 125.12 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.74 124.635 10.88 125.12 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.98 124.635 8.12 125.12 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5 124.635 59.64 125.12 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.66 124.635 11.8 125.12 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.5 124.635 13.64 125.12 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.46 124.635 25.6 125.12 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.54 124.635 24.68 125.12 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.5 124.635 36.64 125.12 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 124.635 61.48 125.12 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.06 124.635 53.2 125.12 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.86 124.635 67 125.12 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.08 124.635 70.22 125.12 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.2 124.635 57.34 125.12 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.42 124.635 60.56 125.12 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.3 124.635 27.44 125.12 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 124.635 35.72 125.12 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 124.635 65.16 125.12 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.94 124.635 66.08 125.12 ;
    END
  END chany_top_in[20]
  PIN chany_top_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.12 124.635 58.26 125.12 ;
    END
  END chany_top_in[21]
  PIN chany_top_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.58 124.635 12.72 125.12 ;
    END
  END chany_top_in[22]
  PIN chany_top_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.42 124.635 14.56 125.12 ;
    END
  END chany_top_in[23]
  PIN chany_top_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.06 124.635 30.2 125.12 ;
    END
  END chany_top_in[24]
  PIN chany_top_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.82 124.635 9.96 125.12 ;
    END
  END chany_top_in[25]
  PIN chany_top_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 124.635 64.24 125.12 ;
    END
  END chany_top_in[26]
  PIN chany_top_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 124.635 56.42 125.12 ;
    END
  END chany_top_in[27]
  PIN chany_top_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71 124.635 71.14 125.12 ;
    END
  END chany_top_in[28]
  PIN chany_top_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.54 124.635 47.68 125.12 ;
    END
  END chany_top_in[29]
  PIN top_left_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.84 124.635 3.98 125.12 ;
    END
  END top_left_grid_pin_1_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 23.56 103.96 23.7 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 109.67 103.96 109.97 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 28.32 103.96 28.46 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 69.12 103.96 69.26 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 110.26 103.96 110.4 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 48.04 103.96 48.18 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 42.6 103.96 42.74 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 109.58 103.96 109.72 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 60.96 103.96 61.1 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 105.16 103.96 105.3 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 102.44 103.96 102.58 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 85.1 103.96 85.24 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 26.28 103.96 26.42 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 106.86 103.96 107 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 50.76 103.96 50.9 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 83.83 103.96 84.13 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 64.02 103.96 64.16 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 47.36 103.96 47.5 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 25.6 103.96 25.74 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 71.84 103.96 71.98 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 98.7 103.96 98.84 ;
    END
  END chanx_right_in[20]
  PIN chanx_right_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 93.6 103.96 93.74 ;
    END
  END chanx_right_in[21]
  PIN chanx_right_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 85.19 103.96 85.49 ;
    END
  END chanx_right_in[22]
  PIN chanx_right_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 82.72 103.96 82.86 ;
    END
  END chanx_right_in[23]
  PIN chanx_right_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 45.32 103.96 45.46 ;
    END
  END chanx_right_in[24]
  PIN chanx_right_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 107.54 103.96 107.68 ;
    END
  END chanx_right_in[25]
  PIN chanx_right_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 97.43 103.96 97.73 ;
    END
  END chanx_right_in[26]
  PIN chanx_right_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 50.08 103.96 50.22 ;
    END
  END chanx_right_in[27]
  PIN chanx_right_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 69.8 103.96 69.94 ;
    END
  END chanx_right_in[28]
  PIN chanx_right_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 83.4 103.96 83.54 ;
    END
  END chanx_right_in[29]
  PIN right_bottom_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 98.79 103.96 99.09 ;
    END
  END right_bottom_grid_pin_1_[0]
  PIN right_bottom_grid_pin_3_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 58.92 103.96 59.06 ;
    END
  END right_bottom_grid_pin_3_[0]
  PIN right_bottom_grid_pin_5_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 93.35 103.96 93.65 ;
    END
  END right_bottom_grid_pin_5_[0]
  PIN right_bottom_grid_pin_7_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 39.88 103.96 40.02 ;
    END
  END right_bottom_grid_pin_7_[0]
  PIN right_bottom_grid_pin_9_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 115.79 103.96 116.09 ;
    END
  END right_bottom_grid_pin_9_[0]
  PIN right_bottom_grid_pin_11_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 114.43 103.96 114.73 ;
    END
  END right_bottom_grid_pin_11_[0]
  PIN right_bottom_grid_pin_13_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 113.07 103.96 113.37 ;
    END
  END right_bottom_grid_pin_13_[0]
  PIN right_bottom_grid_pin_15_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 94.71 103.96 95.01 ;
    END
  END right_bottom_grid_pin_15_[0]
  PIN right_bottom_grid_pin_17_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 100.83 103.96 101.13 ;
    END
  END right_bottom_grid_pin_17_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 61.64 103.96 61.78 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.34 124.635 15.48 125.12 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 124.635 62.4 125.12 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.26 124.635 16.4 125.12 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.06 124.635 7.2 125.12 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.62 124.635 46.76 125.12 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.62 124.635 23.76 125.12 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.9 124.635 9.04 125.12 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.42 124.635 37.56 125.12 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.18 124.635 63.32 125.12 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.18 124.635 17.32 125.12 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.7 124.635 45.84 125.12 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.7 124.635 22.84 125.12 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.38 124.635 26.52 125.12 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.1 124.635 18.24 125.12 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.78 124.635 67.92 125.12 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 124.635 38.48 125.12 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.78 124.635 44.92 125.12 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.78 124.635 21.92 125.12 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.76 124.635 4.9 125.12 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 124.635 39.4 125.12 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.86 124.635 44 125.12 ;
    END
  END chany_top_out[20]
  PIN chany_top_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.02 124.635 19.16 125.12 ;
    END
  END chany_top_out[21]
  PIN chany_top_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.14 124.635 6.28 125.12 ;
    END
  END chany_top_out[22]
  PIN chany_top_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.18 124.635 40.32 125.12 ;
    END
  END chany_top_out[23]
  PIN chany_top_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.22 124.635 28.36 125.12 ;
    END
  END chany_top_out[24]
  PIN chany_top_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.94 124.635 43.08 125.12 ;
    END
  END chany_top_out[25]
  PIN chany_top_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 124.635 41.24 125.12 ;
    END
  END chany_top_out[26]
  PIN chany_top_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.86 124.635 21 125.12 ;
    END
  END chany_top_out[27]
  PIN chany_top_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.94 124.635 20.08 125.12 ;
    END
  END chany_top_out[28]
  PIN chany_top_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.02 124.635 42.16 125.12 ;
    END
  END chany_top_out[29]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 44.64 103.96 44.78 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 77.96 103.96 78.1 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 63.34 103.96 63.48 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 115.02 103.96 115.16 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 115.7 103.96 115.84 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 29 103.96 29.14 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 102.19 103.96 102.49 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 101.42 103.96 101.56 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 80 103.96 80.14 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 113.32 103.96 113.46 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 117.74 103.96 117.88 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 88.16 103.96 88.3 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 94.28 103.96 94.42 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 99.72 103.96 99.86 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 72.52 103.96 72.66 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 97 103.96 97.14 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 95.98 103.96 96.12 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 91.22 103.96 91.36 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 103.55 103.96 103.85 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 104.91 103.96 105.21 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 80.68 103.96 80.82 ;
    END
  END chanx_right_out[20]
  PIN chanx_right_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 104.14 103.96 104.28 ;
    END
  END chanx_right_out[21]
  PIN chanx_right_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 106.27 103.96 106.57 ;
    END
  END chanx_right_out[22]
  PIN chanx_right_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 90.54 103.96 90.68 ;
    END
  END chanx_right_out[23]
  PIN chanx_right_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 96.07 103.96 96.37 ;
    END
  END chanx_right_out[24]
  PIN chanx_right_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 108.31 103.96 108.61 ;
    END
  END chanx_right_out[25]
  PIN chanx_right_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 85.78 103.96 85.92 ;
    END
  END chanx_right_out[26]
  PIN chanx_right_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 112.3 103.96 112.44 ;
    END
  END chanx_right_out[27]
  PIN chanx_right_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 111.71 103.96 112.01 ;
    END
  END chanx_right_out[28]
  PIN chanx_right_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 88.84 103.96 88.98 ;
    END
  END chanx_right_out[29]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.44 0 100.58 0.485 ;
    END
  END ccff_tail[0]
  PIN pReset_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 36.14 103.96 36.28 ;
    END
  END pReset_E_in
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 103.365 7.24 103.96 7.38 ;
    END
  END prog_clk_0_E_in
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 17.44 3.2 20.64 ;
        RECT 100.76 17.44 103.96 20.64 ;
        RECT 0 58.24 3.2 61.44 ;
        RECT 100.76 58.24 103.96 61.44 ;
        RECT 0 99.04 3.2 102.24 ;
        RECT 100.76 99.04 103.96 102.24 ;
      LAYER met4 ;
        RECT 14.42 0 15.02 0.6 ;
        RECT 43.86 0 44.46 0.6 ;
        RECT 89.86 0 90.46 0.6 ;
        RECT 89.86 119.08 90.46 119.68 ;
        RECT 14.42 124.52 15.02 125.12 ;
        RECT 43.86 124.52 44.46 125.12 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 103.48 2.48 103.96 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 103.48 7.92 103.96 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 103.48 13.36 103.96 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 103.48 18.8 103.96 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 103.48 24.24 103.96 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 103.48 29.68 103.96 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 103.48 35.12 103.96 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 103.48 40.56 103.96 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 103.48 46 103.96 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 103.48 51.44 103.96 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 103.48 56.88 103.96 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 103.48 62.32 103.96 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 103.48 67.76 103.96 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 103.48 73.2 103.96 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 103.48 78.64 103.96 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 103.48 84.08 103.96 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 103.48 89.52 103.96 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 103.48 94.96 103.96 95.44 ;
        RECT 0 100.4 0.48 100.88 ;
        RECT 103.48 100.4 103.96 100.88 ;
        RECT 0 105.84 0.48 106.32 ;
        RECT 103.48 105.84 103.96 106.32 ;
        RECT 0 111.28 0.48 111.76 ;
        RECT 103.48 111.28 103.96 111.76 ;
        RECT 0 116.72 0.48 117.2 ;
        RECT 103.48 116.72 103.96 117.2 ;
        RECT 0 122.16 0.48 122.64 ;
        RECT 73.12 122.16 73.6 122.64 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 37.84 3.2 41.04 ;
        RECT 100.76 37.84 103.96 41.04 ;
        RECT 0 78.64 3.2 81.84 ;
        RECT 100.76 78.64 103.96 81.84 ;
      LAYER met4 ;
        RECT 29.14 0 29.74 0.6 ;
        RECT 58.58 0 59.18 0.6 ;
        RECT 29.14 124.52 29.74 125.12 ;
        RECT 58.58 124.52 59.18 125.12 ;
      LAYER met1 ;
        RECT 0 -0.24 0.48 0.24 ;
        RECT 103.48 -0.24 103.96 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 103.48 5.2 103.96 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 103.48 10.64 103.96 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 103.48 16.08 103.96 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 103.48 21.52 103.96 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 103.48 26.96 103.96 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 103.48 32.4 103.96 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 103.48 37.84 103.96 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 103.48 43.28 103.96 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 103.48 48.72 103.96 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 103.48 54.16 103.96 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 103.48 59.6 103.96 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 103.48 65.04 103.96 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 103.48 70.48 103.96 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 103.48 75.92 103.96 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 103.48 81.36 103.96 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 103.48 86.8 103.96 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 103.48 92.24 103.96 92.72 ;
        RECT 0 97.68 0.48 98.16 ;
        RECT 103.48 97.68 103.96 98.16 ;
        RECT 0 103.12 0.48 103.6 ;
        RECT 103.48 103.12 103.96 103.6 ;
        RECT 0 108.56 0.48 109.04 ;
        RECT 103.48 108.56 103.96 109.04 ;
        RECT 0 114 0.48 114.48 ;
        RECT 103.48 114 103.96 114.48 ;
        RECT 0 119.44 0.48 119.92 ;
        RECT 103.48 119.44 103.96 119.92 ;
        RECT 0 124.88 0.48 125.36 ;
        RECT 73.12 124.88 73.6 125.36 ;
    END
  END VSS
  OBS
    LAYER met1 ;
      POLYGON 72.84 125.36 72.84 124.88 59.04 124.88 59.04 124.87 58.72 124.87 58.72 124.88 29.6 124.88 29.6 124.87 29.28 124.87 29.28 124.88 0.76 124.88 0.76 125.36 ;
      RECT 53.96 119.44 103.2 119.92 ;
      POLYGON 59.04 0.25 59.04 0.24 103.2 0.24 103.2 -0.24 0.76 -0.24 0.76 0.24 29.28 0.24 29.28 0.25 29.6 0.25 29.6 0.24 58.72 0.24 58.72 0.25 ;
      POLYGON 72.84 124.84 72.84 124.6 73.32 124.6 73.32 122.92 72.84 122.92 72.84 121.88 73.32 121.88 73.32 119.4 103.2 119.4 103.2 119.16 103.68 119.16 103.68 118.16 103.085 118.16 103.085 117.46 103.2 117.46 103.2 116.44 103.68 116.44 103.68 116.12 103.085 116.12 103.085 114.74 103.2 114.74 103.2 113.74 103.085 113.74 103.085 113.04 103.68 113.04 103.68 112.72 103.085 112.72 103.085 112.02 103.2 112.02 103.2 111 103.68 111 103.68 110.68 103.085 110.68 103.085 109.3 103.2 109.3 103.2 108.28 103.68 108.28 103.68 107.96 103.085 107.96 103.085 106.58 103.2 106.58 103.2 105.58 103.085 105.58 103.085 104.88 103.68 104.88 103.68 104.56 103.085 104.56 103.085 103.86 103.2 103.86 103.2 102.86 103.085 102.86 103.085 102.16 103.68 102.16 103.68 101.84 103.085 101.84 103.085 101.14 103.2 101.14 103.2 100.14 103.085 100.14 103.085 99.44 103.68 99.44 103.68 99.12 103.085 99.12 103.085 98.42 103.2 98.42 103.2 97.42 103.085 97.42 103.085 96.72 103.68 96.72 103.68 96.4 103.085 96.4 103.085 95.7 103.2 95.7 103.2 94.7 103.085 94.7 103.085 93.32 103.68 93.32 103.68 93 103.2 93 103.2 91.96 103.68 91.96 103.68 91.64 103.085 91.64 103.085 90.26 103.2 90.26 103.2 89.26 103.085 89.26 103.085 87.88 103.68 87.88 103.68 87.56 103.2 87.56 103.2 86.52 103.68 86.52 103.68 86.2 103.085 86.2 103.085 84.82 103.2 84.82 103.2 83.82 103.085 83.82 103.085 82.44 103.68 82.44 103.68 82.12 103.2 82.12 103.2 81.1 103.085 81.1 103.085 79.72 103.68 79.72 103.68 79.4 103.2 79.4 103.2 78.38 103.085 78.38 103.085 77.68 103.68 77.68 103.68 76.68 103.2 76.68 103.2 75.64 103.68 75.64 103.68 73.96 103.2 73.96 103.2 72.94 103.085 72.94 103.085 71.56 103.68 71.56 103.68 71.24 103.2 71.24 103.2 70.22 103.085 70.22 103.085 68.84 103.68 68.84 103.68 68.52 103.2 68.52 103.2 67.48 103.68 67.48 103.68 65.8 103.2 65.8 103.2 64.76 103.68 64.76 103.68 64.44 103.085 64.44 103.085 63.06 103.2 63.06 103.2 62.06 103.085 62.06 103.085 60.68 103.68 60.68 103.68 60.36 103.2 60.36 103.2 59.34 103.085 59.34 103.085 58.64 103.68 58.64 103.68 57.64 103.2 57.64 103.2 56.6 103.68 56.6 103.68 54.92 103.2 54.92 103.2 53.88 103.68 53.88 103.68 52.2 103.2 52.2 103.2 51.18 103.085 51.18 103.085 49.8 103.68 49.8 103.68 49.48 103.2 49.48 103.2 48.46 103.085 48.46 103.085 47.08 103.68 47.08 103.68 46.76 103.2 46.76 103.2 45.74 103.085 45.74 103.085 44.36 103.68 44.36 103.68 44.04 103.2 44.04 103.2 43.02 103.085 43.02 103.085 42.32 103.68 42.32 103.68 41.32 103.2 41.32 103.2 40.3 103.085 40.3 103.085 39.6 103.68 39.6 103.68 38.6 103.2 38.6 103.2 37.56 103.68 37.56 103.68 36.56 103.085 36.56 103.085 35.86 103.2 35.86 103.2 34.84 103.68 34.84 103.68 33.16 103.2 33.16 103.2 32.12 103.68 32.12 103.68 30.44 103.2 30.44 103.2 29.42 103.085 29.42 103.085 28.04 103.68 28.04 103.68 27.72 103.2 27.72 103.2 26.7 103.085 26.7 103.085 25.32 103.68 25.32 103.68 25 103.2 25 103.2 23.98 103.085 23.98 103.085 23.28 103.68 23.28 103.68 22.28 103.2 22.28 103.2 21.24 103.68 21.24 103.68 19.56 103.2 19.56 103.2 18.52 103.68 18.52 103.68 16.84 103.2 16.84 103.2 15.8 103.68 15.8 103.68 14.12 103.2 14.12 103.2 13.08 103.68 13.08 103.68 11.4 103.2 11.4 103.2 10.36 103.68 10.36 103.68 8.68 103.2 8.68 103.2 7.66 103.085 7.66 103.085 6.96 103.68 6.96 103.68 5.96 103.2 5.96 103.2 4.92 103.68 4.92 103.68 3.24 103.2 3.24 103.2 2.2 103.68 2.2 103.68 0.52 103.2 0.52 103.2 0.28 0.76 0.28 0.76 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.06 0.875 63.06 0.875 63.76 0.28 63.76 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 0.76 97.4 0.76 98.44 0.28 98.44 0.28 100.12 0.76 100.12 0.76 101.16 0.28 101.16 0.28 102.84 0.76 102.84 0.76 103.88 0.28 103.88 0.28 105.56 0.76 105.56 0.76 106.6 0.28 106.6 0.28 108.28 0.76 108.28 0.76 109.32 0.28 109.32 0.28 111 0.76 111 0.76 112.04 0.28 112.04 0.28 113.72 0.76 113.72 0.76 114.76 0.28 114.76 0.28 116.44 0.76 116.44 0.76 117.48 0.28 117.48 0.28 119.16 0.76 119.16 0.76 120.2 0.28 120.2 0.28 121.88 0.76 121.88 0.76 122.92 0.28 122.92 0.28 124.6 0.76 124.6 0.76 124.84 ;
    LAYER met4 ;
      POLYGON 51.225 124.945 51.225 124.615 51.21 124.615 51.21 62.07 50.91 62.07 50.91 124.615 50.895 124.615 50.895 124.945 ;
      POLYGON 49.385 124.945 49.385 124.615 49.37 124.615 49.37 49.83 49.07 49.83 49.07 124.615 49.055 124.615 49.055 124.945 ;
      POLYGON 73.305 119.505 73.305 119.175 73.29 119.175 73.29 91.99 72.99 91.99 72.99 119.175 72.975 119.175 72.975 119.505 ;
      POLYGON 73.2 124.72 73.2 119.28 89.46 119.28 89.46 118.68 90.86 118.68 90.86 119.28 103.56 119.28 103.56 0.4 90.86 0.4 90.86 1 89.46 1 89.46 0.4 59.58 0.4 59.58 1 58.18 1 58.18 0.4 44.86 0.4 44.86 1 43.46 1 43.46 0.4 30.14 0.4 30.14 1 28.74 1 28.74 0.4 15.42 0.4 15.42 1 14.02 1 14.02 0.4 0.4 0.4 0.4 124.72 14.02 124.72 14.02 124.12 15.42 124.12 15.42 124.72 19.23 124.72 19.23 123.92 20.33 123.92 20.33 124.72 28.74 124.72 28.74 124.12 30.14 124.12 30.14 124.72 43.46 124.72 43.46 124.12 44.86 124.12 44.86 124.72 58.18 124.72 58.18 124.12 59.58 124.12 59.58 124.72 ;
    LAYER met2 ;
      RECT 58.74 124.815 59.02 125.185 ;
      RECT 29.3 124.815 29.58 125.185 ;
      POLYGON 22.38 125.02 22.38 119.95 22.24 119.95 22.24 124.88 22.2 124.88 22.2 125.02 ;
      POLYGON 14.14 125.02 14.14 124.88 14.1 124.88 14.1 121.31 13.96 121.31 13.96 125.02 ;
      POLYGON 13.22 125.02 13.22 124.88 13.18 124.88 13.18 110.6 13.04 110.6 13.04 125.02 ;
      RECT 37.82 124.45 38.08 124.77 ;
      RECT 69.1 124.11 69.36 124.43 ;
      RECT 62.66 124.11 62.92 124.43 ;
      RECT 59.9 124.11 60.16 124.43 ;
      RECT 35.98 124.11 36.24 124.43 ;
      RECT 24.94 124.11 25.2 124.43 ;
      POLYGON 73.44 120.26 73.44 112.98 73.3 112.98 73.3 120.12 72.38 120.12 72.38 120.26 ;
      RECT 58.74 -0.065 59.02 0.305 ;
      RECT 29.3 -0.065 29.58 0.305 ;
      POLYGON 73.32 124.84 73.32 119.4 103.68 119.4 103.68 0.28 100.86 0.28 100.86 0.765 100.16 0.765 100.16 0.28 0.28 0.28 0.28 124.84 3.56 124.84 3.56 124.355 4.26 124.355 4.26 124.84 4.48 124.84 4.48 124.355 5.18 124.355 5.18 124.84 5.86 124.84 5.86 124.355 6.56 124.355 6.56 124.84 6.78 124.84 6.78 124.355 7.48 124.355 7.48 124.84 7.7 124.84 7.7 124.355 8.4 124.355 8.4 124.84 8.62 124.84 8.62 124.355 9.32 124.355 9.32 124.84 9.54 124.84 9.54 124.355 10.24 124.355 10.24 124.84 10.46 124.84 10.46 124.355 11.16 124.355 11.16 124.84 11.38 124.84 11.38 124.355 12.08 124.355 12.08 124.84 12.3 124.84 12.3 124.355 13 124.355 13 124.84 13.22 124.84 13.22 124.355 13.92 124.355 13.92 124.84 14.14 124.84 14.14 124.355 14.84 124.355 14.84 124.84 15.06 124.84 15.06 124.355 15.76 124.355 15.76 124.84 15.98 124.84 15.98 124.355 16.68 124.355 16.68 124.84 16.9 124.84 16.9 124.355 17.6 124.355 17.6 124.84 17.82 124.84 17.82 124.355 18.52 124.355 18.52 124.84 18.74 124.84 18.74 124.355 19.44 124.355 19.44 124.84 19.66 124.84 19.66 124.355 20.36 124.355 20.36 124.84 20.58 124.84 20.58 124.355 21.28 124.355 21.28 124.84 21.5 124.84 21.5 124.355 22.2 124.355 22.2 124.84 22.42 124.84 22.42 124.355 23.12 124.355 23.12 124.84 23.34 124.84 23.34 124.355 24.04 124.355 24.04 124.84 24.26 124.84 24.26 124.355 24.96 124.355 24.96 124.84 25.18 124.84 25.18 124.355 25.88 124.355 25.88 124.84 26.1 124.84 26.1 124.355 26.8 124.355 26.8 124.84 27.02 124.84 27.02 124.355 27.72 124.355 27.72 124.84 27.94 124.84 27.94 124.355 28.64 124.355 28.64 124.84 29.78 124.84 29.78 124.355 30.48 124.355 30.48 124.84 35.3 124.84 35.3 124.355 36 124.355 36 124.84 36.22 124.84 36.22 124.355 36.92 124.355 36.92 124.84 37.14 124.84 37.14 124.355 37.84 124.355 37.84 124.84 38.06 124.84 38.06 124.355 38.76 124.355 38.76 124.84 38.98 124.84 38.98 124.355 39.68 124.355 39.68 124.84 39.9 124.84 39.9 124.355 40.6 124.355 40.6 124.84 40.82 124.84 40.82 124.355 41.52 124.355 41.52 124.84 41.74 124.84 41.74 124.355 42.44 124.355 42.44 124.84 42.66 124.84 42.66 124.355 43.36 124.355 43.36 124.84 43.58 124.84 43.58 124.355 44.28 124.355 44.28 124.84 44.5 124.84 44.5 124.355 45.2 124.355 45.2 124.84 45.42 124.84 45.42 124.355 46.12 124.355 46.12 124.84 46.34 124.84 46.34 124.355 47.04 124.355 47.04 124.84 47.26 124.84 47.26 124.355 47.96 124.355 47.96 124.84 52.78 124.84 52.78 124.355 53.48 124.355 53.48 124.84 55.08 124.84 55.08 124.355 55.78 124.355 55.78 124.84 56 124.84 56 124.355 56.7 124.355 56.7 124.84 56.92 124.84 56.92 124.355 57.62 124.355 57.62 124.84 57.84 124.84 57.84 124.355 58.54 124.355 58.54 124.84 59.22 124.84 59.22 124.355 59.92 124.355 59.92 124.84 60.14 124.84 60.14 124.355 60.84 124.355 60.84 124.84 61.06 124.84 61.06 124.355 61.76 124.355 61.76 124.84 61.98 124.84 61.98 124.355 62.68 124.355 62.68 124.84 62.9 124.84 62.9 124.355 63.6 124.355 63.6 124.84 63.82 124.84 63.82 124.355 64.52 124.355 64.52 124.84 64.74 124.84 64.74 124.355 65.44 124.355 65.44 124.84 65.66 124.84 65.66 124.355 66.36 124.355 66.36 124.84 66.58 124.84 66.58 124.355 67.28 124.355 67.28 124.84 67.5 124.84 67.5 124.355 68.2 124.355 68.2 124.84 68.42 124.84 68.42 124.355 69.12 124.355 69.12 124.84 69.8 124.84 69.8 124.355 70.5 124.355 70.5 124.84 70.72 124.84 70.72 124.355 71.42 124.355 71.42 124.84 ;
    LAYER met3 ;
      POLYGON 59.045 125.165 59.045 125.16 59.26 125.16 59.26 124.84 59.045 124.84 59.045 124.835 58.715 124.835 58.715 124.84 58.5 124.84 58.5 125.16 58.715 125.16 58.715 125.165 ;
      POLYGON 29.605 125.165 29.605 125.16 29.82 125.16 29.82 124.84 29.605 124.84 29.605 124.835 29.275 124.835 29.275 124.84 29.06 124.84 29.06 125.16 29.275 125.16 29.275 125.165 ;
      POLYGON 55.595 124.945 55.595 124.615 55.265 124.615 55.265 124.63 51.25 124.63 51.25 124.62 50.87 124.62 50.87 124.94 51.25 124.94 51.25 124.93 55.265 124.93 55.265 124.945 ;
      POLYGON 45.015 124.945 45.015 124.93 49.03 124.93 49.03 124.94 49.41 124.94 49.41 124.62 49.03 124.62 49.03 124.63 45.015 124.63 45.015 124.615 44.685 124.615 44.685 124.945 ;
      POLYGON 73.33 119.5 73.33 119.18 72.95 119.18 72.95 119.19 70.92 119.19 70.92 119.49 72.95 119.49 72.95 119.5 ;
      POLYGON 59.045 0.285 59.045 0.28 59.26 0.28 59.26 -0.04 59.045 -0.04 59.045 -0.045 58.715 -0.045 58.715 -0.04 58.5 -0.04 58.5 0.28 58.715 0.28 58.715 0.285 ;
      POLYGON 29.605 0.285 29.605 0.28 29.82 0.28 29.82 -0.04 29.605 -0.04 29.605 -0.045 29.275 -0.045 29.275 -0.04 29.06 -0.04 29.06 0.28 29.275 0.28 29.275 0.285 ;
      POLYGON 73.2 124.72 73.2 119.28 103.56 119.28 103.56 116.49 102.76 116.49 102.76 115.39 103.56 115.39 103.56 115.13 102.76 115.13 102.76 114.03 103.56 114.03 103.56 113.77 102.76 113.77 102.76 112.67 103.56 112.67 103.56 112.41 102.76 112.41 102.76 111.31 103.56 111.31 103.56 110.37 102.76 110.37 102.76 109.27 103.56 109.27 103.56 109.01 102.76 109.01 102.76 107.91 103.56 107.91 103.56 106.97 102.76 106.97 102.76 105.87 103.56 105.87 103.56 105.61 102.76 105.61 102.76 104.51 103.56 104.51 103.56 104.25 102.76 104.25 102.76 103.15 103.56 103.15 103.56 102.89 102.76 102.89 102.76 101.79 103.56 101.79 103.56 101.53 102.76 101.53 102.76 100.43 103.56 100.43 103.56 99.49 102.76 99.49 102.76 98.39 103.56 98.39 103.56 98.13 102.76 98.13 102.76 97.03 103.56 97.03 103.56 96.77 102.76 96.77 102.76 95.67 103.56 95.67 103.56 95.41 102.76 95.41 102.76 94.31 103.56 94.31 103.56 94.05 102.76 94.05 102.76 92.95 103.56 92.95 103.56 85.89 102.76 85.89 102.76 84.79 103.56 84.79 103.56 84.53 102.76 84.53 102.76 83.43 103.56 83.43 103.56 0.4 0.4 0.4 0.4 124.72 ;
    LAYER met5 ;
      POLYGON 72 123.52 72 118.08 102.36 118.08 102.36 103.84 99.16 103.84 99.16 97.44 102.36 97.44 102.36 83.44 99.16 83.44 99.16 77.04 102.36 77.04 102.36 63.04 99.16 63.04 99.16 56.64 102.36 56.64 102.36 42.64 99.16 42.64 99.16 36.24 102.36 36.24 102.36 22.24 99.16 22.24 99.16 15.84 102.36 15.84 102.36 1.6 1.6 1.6 1.6 15.84 4.8 15.84 4.8 22.24 1.6 22.24 1.6 36.24 4.8 36.24 4.8 42.64 1.6 42.64 1.6 56.64 4.8 56.64 4.8 63.04 1.6 63.04 1.6 77.04 4.8 77.04 4.8 83.44 1.6 83.44 1.6 97.44 4.8 97.44 4.8 103.84 1.6 103.84 1.6 123.52 ;
    LAYER li1 ;
      POLYGON 73.6 125.205 73.6 125.035 69.395 125.035 69.395 124.655 69.065 124.655 69.065 125.035 67.07 125.035 67.07 124.235 66.815 124.235 66.815 125.035 66.225 125.035 66.225 124.655 65.895 124.655 65.895 125.035 63.81 125.035 63.81 124.535 63.61 124.535 63.61 125.035 57.905 125.035 57.905 124.575 57.6 124.575 57.6 125.035 56.115 125.035 56.115 124.595 55.925 124.595 55.925 125.035 54.025 125.035 54.025 124.575 53.695 124.575 53.695 125.035 51.095 125.035 51.095 124.675 50.765 124.675 50.765 125.035 50.065 125.035 50.065 124.655 49.735 124.655 49.735 125.035 42.265 125.035 42.265 124.635 41.935 124.635 41.935 125.035 39.975 125.035 39.975 124.5 39.465 124.5 39.465 125.035 32.145 125.035 32.145 124.575 31.84 124.575 31.84 125.035 30.355 125.035 30.355 124.595 30.165 124.595 30.165 125.035 28.265 125.035 28.265 124.575 27.935 124.575 27.935 125.035 25.335 125.035 25.335 124.675 25.005 124.675 25.005 125.035 24.305 125.035 24.305 124.655 23.975 124.655 23.975 125.035 18.765 125.035 18.765 124.235 18.435 124.235 18.435 125.035 17.925 125.035 17.925 124.555 17.595 124.555 17.595 125.035 17.085 125.035 17.085 124.555 16.755 124.555 16.755 125.035 16.165 125.035 16.165 124.555 15.995 124.555 15.995 125.035 15.325 125.035 15.325 124.555 15.155 124.555 15.155 125.035 0 125.035 0 125.205 ;
      RECT 69.92 122.315 73.6 122.485 ;
      RECT 0 122.315 3.68 122.485 ;
      POLYGON 103.96 119.765 103.96 119.595 99.725 119.595 99.725 118.795 99.395 118.795 99.395 119.595 98.885 119.595 98.885 119.115 98.555 119.115 98.555 119.595 98.045 119.595 98.045 119.115 97.715 119.115 97.715 119.595 97.125 119.595 97.125 119.115 96.955 119.115 96.955 119.595 96.285 119.595 96.285 119.115 96.115 119.115 96.115 119.595 94.785 119.595 94.785 119.115 94.615 119.115 94.615 119.595 93.945 119.595 93.945 119.115 93.775 119.115 93.775 119.595 93.185 119.595 93.185 119.115 92.855 119.115 92.855 119.595 92.345 119.595 92.345 119.115 92.015 119.115 92.015 119.595 91.505 119.595 91.505 118.795 91.175 118.795 91.175 119.595 88.265 119.595 88.265 119.135 87.96 119.135 87.96 119.595 86.475 119.595 86.475 119.155 86.285 119.155 86.285 119.595 84.385 119.595 84.385 119.135 84.055 119.135 84.055 119.595 81.455 119.595 81.455 119.235 81.125 119.235 81.125 119.595 80.425 119.595 80.425 119.215 80.095 119.215 80.095 119.595 73.085 119.595 73.085 119.135 72.78 119.135 72.78 119.595 71.295 119.595 71.295 119.155 71.105 119.155 71.105 119.595 69.205 119.595 69.205 119.135 68.875 119.135 68.875 119.595 66.275 119.595 66.275 119.235 65.945 119.235 65.945 119.595 65.245 119.595 65.245 119.215 64.915 119.215 64.915 119.595 64.4 119.595 64.4 119.765 ;
      RECT 0 119.595 3.68 119.765 ;
      RECT 103.5 116.875 103.96 117.045 ;
      RECT 0 116.875 3.68 117.045 ;
      RECT 103.04 114.155 103.96 114.325 ;
      RECT 0 114.155 3.68 114.325 ;
      RECT 103.04 111.435 103.96 111.605 ;
      RECT 0 111.435 3.68 111.605 ;
      RECT 103.04 108.715 103.96 108.885 ;
      RECT 0 108.715 3.68 108.885 ;
      RECT 102.12 105.995 103.96 106.165 ;
      RECT 0 105.995 3.68 106.165 ;
      RECT 102.12 103.275 103.96 103.445 ;
      RECT 0 103.275 3.68 103.445 ;
      RECT 103.04 100.555 103.96 100.725 ;
      RECT 0 100.555 3.68 100.725 ;
      RECT 103.04 97.835 103.96 98.005 ;
      RECT 0 97.835 3.68 98.005 ;
      RECT 103.04 95.115 103.96 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 103.04 92.395 103.96 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 103.04 89.675 103.96 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 103.04 86.955 103.96 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 103.04 84.235 103.96 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 103.04 81.515 103.96 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 103.04 78.795 103.96 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 100.28 76.075 103.96 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 100.28 73.355 103.96 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 103.04 70.635 103.96 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 103.04 67.915 103.96 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 103.04 65.195 103.96 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 103.04 62.475 103.96 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 103.04 59.755 103.96 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 103.04 57.035 103.96 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 100.28 54.315 103.96 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 100.28 51.595 103.96 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 103.04 48.875 103.96 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 100.28 46.155 103.96 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 100.28 43.435 103.96 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 103.04 40.715 103.96 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 103.04 37.995 103.96 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 103.5 35.275 103.96 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 103.04 32.555 103.96 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 103.04 29.835 103.96 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 103.5 27.115 103.96 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 103.04 24.395 103.96 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 103.04 21.675 103.96 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 103.04 18.955 103.96 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 103.04 16.235 103.96 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 103.04 13.515 103.96 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 103.04 10.795 103.96 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 103.04 8.075 103.96 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 103.04 5.355 103.96 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 103.04 2.635 103.96 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 103.96 0.085 ;
      POLYGON 73.43 124.95 73.43 119.51 103.79 119.51 103.79 0.17 0.17 0.17 0.17 124.95 ;
    LAYER via ;
      RECT 58.805 124.925 58.955 125.075 ;
      RECT 29.365 124.925 29.515 125.075 ;
      RECT 15.335 124.535 15.485 124.685 ;
      RECT 58.805 0.045 58.955 0.195 ;
      RECT 29.365 0.045 29.515 0.195 ;
    LAYER via2 ;
      RECT 58.78 124.9 58.98 125.1 ;
      RECT 29.34 124.9 29.54 125.1 ;
      RECT 55.33 124.68 55.53 124.88 ;
      RECT 44.75 124.68 44.95 124.88 ;
      RECT 58.78 0.02 58.98 0.22 ;
      RECT 29.34 0.02 29.54 0.22 ;
    LAYER via3 ;
      RECT 58.78 124.9 58.98 125.1 ;
      RECT 29.34 124.9 29.54 125.1 ;
      RECT 50.96 124.68 51.16 124.88 ;
      RECT 49.12 124.68 49.32 124.88 ;
      RECT 73.04 119.24 73.24 119.44 ;
      RECT 58.78 0.02 58.98 0.22 ;
      RECT 29.34 0.02 29.54 0.22 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 125.12 73.6 125.12 73.6 119.68 103.96 119.68 103.96 0 ;
  END
END sb_0__0_

END LIBRARY
