//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module sky130_fd_sc_hd__inv_1
(
    A,
    Y
);

    input A;
    output Y;

    wire A;
    wire Y;

endmodule

module sky130_fd_sc_hd__buf_2
(
    A,
    X
);

    input A;
    output X;

    wire A;
    wire X;

endmodule

module sky130_fd_sc_hd__buf_4
(
    A,
    X
);

    input A;
    output X;

    wire A;
    wire X;

endmodule

module sky130_fd_sc_hd__inv_2
(
    A,
    Y
);

    input A;
    output Y;

    wire A;
    wire Y;

endmodule

module sky130_fd_sc_hd__or2_1
(
    A,
    B,
    X
);

    input A;
    input B;
    output X;

    wire A;
    wire B;
    wire X;

endmodule

module sky130_fd_sc_hd__mux2_1
(
    A1,
    A0,
    S,
    X
);

    input A1;
    input A0;
    input S;
    output X;

    wire A1;
    wire A0;
    wire S;
    wire X;

endmodule

module sky130_fd_sc_hd__sdfrtp_1
(
    SCE,
    D,
    SCD,
    RESET_B,
    CLK,
    Q
);

    input SCE;
    input D;
    input SCD;
    input RESET_B;
    input CLK;
    output Q;

    wire SCE;
    wire D;
    wire SCD;
    wire RESET_B;
    wire CLK;
    wire Q;

endmodule

module sky130_fd_sc_hd__dfrtp_1
(
    RESET_B,
    CLK,
    D,
    Q
);

    input RESET_B;
    input CLK;
    input D;
    output Q;

    wire RESET_B;
    wire CLK;
    wire D;
    wire Q;

endmodule

module io
(
    IO_ISOL_N,
    SOC_IN,
    SOC_OUT,
    SOC_DIR,
    FPGA_OUT,
    FPGA_DIR,
    FPGA_IN
);

    input IO_ISOL_N;
    input SOC_IN;
    output SOC_OUT;
    output SOC_DIR;
    input FPGA_OUT;
    input FPGA_DIR;
    output FPGA_IN;

    wire IO_ISOL_N;
    wire SOC_IN;
    wire SOC_OUT;
    wire SOC_DIR;
    wire FPGA_OUT;
    wire FPGA_DIR;
    wire FPGA_IN;

endmodule

module sky130_fd_sc_hd__mux2_1_wrapper
(
    A0,
    A1,
    S,
    X
);

    input A0;
    input A1;
    input S;
    output X;

    wire A0;
    wire A1;
    wire S;
    wire X;

endmodule

