VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_2__2_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 92 BY 97.92 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met3 ;
        RECT 0 35.21 1.38 35.51 ;
    END
  END prog_clk[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.59 0 55.73 1.36 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.53 0 50.67 1.36 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.89 0 57.19 1.36 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.85 0 46.99 1.36 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.21 0 54.35 1.36 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.29 0 53.43 1.36 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.39 0 69.53 1.36 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.95 0 63.09 1.36 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.61 0 72.75 1.36 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.79 0 64.93 1.36 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.95 0 40.09 1.36 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.03 0 62.17 1.36 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.71 0 42.85 1.36 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.09 0 44.23 1.36 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.51 0 56.65 1.36 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.19 0 60.33 1.36 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.47 0 68.61 1.36 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.53 0 73.67 1.36 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.45 0 74.59 1.36 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.11 0 61.25 1.36 ;
    END
  END chany_bottom_in[19]
  PIN bottom_right_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.03 0 39.17 1.36 ;
    END
  END bottom_right_grid_pin_1_[0]
  PIN bottom_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 12.73 10.88 13.03 12.24 ;
    END
  END bottom_left_grid_pin_42_[0]
  PIN bottom_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 9.05 10.88 9.35 12.24 ;
    END
  END bottom_left_grid_pin_43_[0]
  PIN bottom_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.33 10.88 18.47 12.24 ;
    END
  END bottom_left_grid_pin_44_[0]
  PIN bottom_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.29 10.88 7.43 12.24 ;
    END
  END bottom_left_grid_pin_45_[0]
  PIN bottom_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.13 10.88 9.27 12.24 ;
    END
  END bottom_left_grid_pin_46_[0]
  PIN bottom_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.11 10.88 15.25 12.24 ;
    END
  END bottom_left_grid_pin_47_[0]
  PIN bottom_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.21 10.88 8.35 12.24 ;
    END
  END bottom_left_grid_pin_48_[0]
  PIN bottom_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.05 10.88 10.19 12.24 ;
    END
  END bottom_left_grid_pin_49_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.69 1.38 42.99 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 54.93 1.38 55.23 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 49.49 1.38 49.79 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 21.61 1.38 21.91 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.97 1.38 23.27 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.17 1.38 33.47 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 26.37 1.38 26.67 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.09 1.38 29.39 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 41.33 1.38 41.63 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.29 1.38 56.59 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 57.65 1.38 57.95 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.01 1.38 59.31 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 18.89 1.38 19.19 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 20.25 1.38 20.55 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 17.53 1.38 17.83 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 30.45 1.38 30.75 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 64.45 1.38 64.75 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.85 1.38 51.15 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.21 1.38 69.51 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 38.61 1.38 38.91 ;
    END
  END chanx_left_in[19]
  PIN left_top_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 61.05 1.38 61.35 ;
    END
  END left_top_grid_pin_1_[0]
  PIN left_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.99 0 28.13 1.36 ;
    END
  END left_bottom_grid_pin_34_[0]
  PIN left_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.81 10.88 12.95 12.24 ;
    END
  END left_bottom_grid_pin_35_[0]
  PIN left_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.99 10.88 5.13 12.24 ;
    END
  END left_bottom_grid_pin_36_[0]
  PIN left_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.07 10.88 4.21 12.24 ;
    END
  END left_bottom_grid_pin_37_[0]
  PIN left_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.37 10.88 6.51 12.24 ;
    END
  END left_bottom_grid_pin_38_[0]
  PIN left_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 4.45 10.88 4.75 12.24 ;
    END
  END left_bottom_grid_pin_39_[0]
  PIN left_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.89 10.88 12.03 12.24 ;
    END
  END left_bottom_grid_pin_40_[0]
  PIN left_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.03 10.88 16.17 12.24 ;
    END
  END left_bottom_grid_pin_41_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.23 96.56 2.37 97.92 ;
    END
  END ccff_head[0]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.87 0 64.01 1.36 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.73 0 59.03 1.36 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.81 0 81.95 1.36 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.87 0 41.01 1.36 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.19 0 37.33 1.36 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.79 0 41.93 1.36 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.17 0 66.31 1.36 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.77 0 47.91 1.36 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 0 57.57 1.36 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.11 0 38.25 1.36 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.69 0 71.83 1.36 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.97 0 34.11 1.36 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.81 0 58.95 1.36 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.13 0 32.27 1.36 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.09 0 67.23 1.36 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.15 0 49.29 1.36 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.37 0 52.51 1.36 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 0 45.61 1.36 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.77 0 70.91 1.36 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.21 0 31.35 1.36 ;
    END
  END chany_bottom_out[19]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 71.93 1.38 72.23 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 89.61 1.38 89.91 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 73.29 1.38 73.59 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.21 1.38 52.51 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 70.57 1.38 70.87 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 67.85 1.38 68.15 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 46.77 1.38 47.07 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.13 1.38 48.43 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 77.37 1.38 77.67 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.05 1.38 44.35 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 53.57 1.38 53.87 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.25 1.38 37.55 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 74.65 1.38 74.95 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 27.73 1.38 28.03 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 63.09 1.38 63.39 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.97 1.38 40.27 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 24.33 1.38 24.63 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.81 1.38 32.11 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 45.41 1.38 45.71 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 65.81 1.38 66.11 ;
    END
  END chanx_left_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 14.81 1.38 15.11 ;
    END
  END ccff_tail[0]
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 16.17 1.38 16.47 ;
    END
  END SC_IN_TOP
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 78.73 1.38 79.03 ;
    END
  END SC_IN_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.21 96.56 31.35 97.92 ;
    END
  END SC_OUT_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 76.01 1.38 76.31 ;
    END
  END SC_OUT_BOT
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 25.76 2.48 26.24 2.96 ;
        RECT 91.52 2.48 92 2.96 ;
        RECT 25.76 7.92 26.24 8.4 ;
        RECT 91.52 7.92 92 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 91.52 13.36 92 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 91.52 18.8 92 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 91.52 24.24 92 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 91.52 29.68 92 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 91.52 35.12 92 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 91.52 40.56 92 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 91.52 46 92 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 91.52 51.44 92 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 91.52 56.88 92 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 91.52 62.32 92 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 91.52 67.76 92 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 91.52 73.2 92 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 91.52 78.64 92 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 91.52 84.08 92 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 91.52 89.52 92 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 91.52 94.96 92 95.44 ;
      LAYER met4 ;
        RECT 36.5 0 37.1 0.6 ;
        RECT 65.94 0 66.54 0.6 ;
        RECT 36.5 97.32 37.1 97.92 ;
        RECT 65.94 97.32 66.54 97.92 ;
      LAYER met5 ;
        RECT 0 22.2 3.2 25.4 ;
        RECT 88.8 22.2 92 25.4 ;
        RECT 0 63 3.2 66.2 ;
        RECT 88.8 63 92 66.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 25.76 0 92 0.24 ;
        RECT 25.76 5.2 26.24 5.68 ;
        RECT 91.52 5.2 92 5.68 ;
        RECT 0 10.64 92 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 91.52 16.08 92 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 91.52 21.52 92 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 91.52 26.96 92 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 91.52 32.4 92 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 91.52 37.84 92 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 91.52 43.28 92 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 91.52 48.72 92 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 91.52 54.16 92 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 91.52 59.6 92 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 91.52 65.04 92 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 91.52 70.48 92 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 91.52 75.92 92 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 91.52 81.36 92 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 91.52 86.8 92 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 91.52 92.24 92 92.72 ;
        RECT 0 97.68 92 97.92 ;
      LAYER met4 ;
        RECT 51.22 0 51.82 0.6 ;
        RECT 80.66 0 81.26 0.6 ;
        RECT 10.74 10.88 11.34 11.48 ;
        RECT 10.74 97.32 11.34 97.92 ;
        RECT 51.22 97.32 51.82 97.92 ;
        RECT 80.66 97.32 81.26 97.92 ;
      LAYER met5 ;
        RECT 0 42.6 3.2 45.8 ;
        RECT 88.8 42.6 92 45.8 ;
        RECT 0 83.4 3.2 86.6 ;
        RECT 88.8 83.4 92 86.6 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 0 97.835 92 98.005 ;
      RECT 91.54 95.115 92 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 91.54 92.395 92 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 91.54 89.675 92 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 91.54 86.955 92 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 91.54 84.235 92 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 91.54 81.515 92 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 91.54 78.795 92 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 88.32 76.075 92 76.245 ;
      RECT 0 76.075 1.84 76.245 ;
      RECT 88.32 73.355 92 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 88.32 70.635 92 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 88.32 67.915 92 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 91.54 65.195 92 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 91.54 62.475 92 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 91.08 59.755 92 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 91.08 57.035 92 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 90.16 54.315 92 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 90.16 51.595 92 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 90.16 48.875 92 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 90.16 46.155 92 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 91.54 43.435 92 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 91.54 40.715 92 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 91.08 37.995 92 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 91.08 35.275 92 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 91.54 32.555 92 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 91.54 29.835 92 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 91.54 27.115 92 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 91.54 24.395 92 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 91.08 21.675 92 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 91.08 18.955 92 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 91.54 16.235 92 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 91.54 13.515 92 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 91.08 10.795 92 10.965 ;
      RECT 0 10.795 29.44 10.965 ;
      RECT 91.08 8.075 92 8.245 ;
      RECT 25.76 8.075 29.44 8.245 ;
      RECT 88.32 5.355 92 5.525 ;
      RECT 25.76 5.355 27.6 5.525 ;
      RECT 88.32 2.635 92 2.805 ;
      RECT 25.76 2.635 29.44 2.805 ;
      RECT 25.76 -0.085 92 0.085 ;
    LAYER met3 ;
      POLYGON 81.125 98.085 81.125 98.08 81.34 98.08 81.34 97.76 81.125 97.76 81.125 97.755 80.795 97.755 80.795 97.76 80.58 97.76 80.58 98.08 80.795 98.08 80.795 98.085 ;
      POLYGON 51.685 98.085 51.685 98.08 51.9 98.08 51.9 97.76 51.685 97.76 51.685 97.755 51.355 97.755 51.355 97.76 51.14 97.76 51.14 98.08 51.355 98.08 51.355 98.085 ;
      POLYGON 11.205 98.085 11.205 98.08 11.42 98.08 11.42 97.76 11.205 97.76 11.205 97.755 10.875 97.755 10.875 97.76 10.66 97.76 10.66 98.08 10.875 98.08 10.875 98.085 ;
      POLYGON 28.67 68.83 28.67 68.53 1.23 68.53 1.23 68.81 1.78 68.81 1.78 68.83 ;
      POLYGON 2.03 18.52 2.03 18.51 6.13 18.51 6.13 18.21 2.03 18.21 2.03 18.2 1.65 18.2 1.65 18.52 ;
      POLYGON 24.53 17.15 24.53 16.85 1.23 16.85 1.23 17.13 1.78 17.13 1.78 17.15 ;
      POLYGON 11.205 11.045 11.205 11.04 11.42 11.04 11.42 10.72 11.205 10.72 11.205 10.715 10.875 10.715 10.875 10.72 10.66 10.72 10.66 11.04 10.875 11.04 10.875 11.045 ;
      POLYGON 81.125 0.165 81.125 0.16 81.34 0.16 81.34 -0.16 81.125 -0.16 81.125 -0.165 80.795 -0.165 80.795 -0.16 80.58 -0.16 80.58 0.16 80.795 0.16 80.795 0.165 ;
      POLYGON 51.685 0.165 51.685 0.16 51.9 0.16 51.9 -0.16 51.685 -0.16 51.685 -0.165 51.355 -0.165 51.355 -0.16 51.14 -0.16 51.14 0.16 51.355 0.16 51.355 0.165 ;
      POLYGON 91.6 97.52 91.6 0.4 26.16 0.4 26.16 11.28 0.4 11.28 0.4 14.41 1.78 14.41 1.78 15.51 0.4 15.51 0.4 15.77 1.78 15.77 1.78 16.87 0.4 16.87 0.4 17.13 1.78 17.13 1.78 18.23 0.4 18.23 0.4 18.49 1.78 18.49 1.78 19.59 0.4 19.59 0.4 19.85 1.78 19.85 1.78 20.95 0.4 20.95 0.4 21.21 1.78 21.21 1.78 22.31 0.4 22.31 0.4 22.57 1.78 22.57 1.78 23.67 0.4 23.67 0.4 23.93 1.78 23.93 1.78 25.03 0.4 25.03 0.4 25.97 1.78 25.97 1.78 27.07 0.4 27.07 0.4 27.33 1.78 27.33 1.78 28.43 0.4 28.43 0.4 28.69 1.78 28.69 1.78 29.79 0.4 29.79 0.4 30.05 1.78 30.05 1.78 31.15 0.4 31.15 0.4 31.41 1.78 31.41 1.78 32.51 0.4 32.51 0.4 32.77 1.78 32.77 1.78 33.87 0.4 33.87 0.4 34.81 1.78 34.81 1.78 35.91 0.4 35.91 0.4 36.85 1.78 36.85 1.78 37.95 0.4 37.95 0.4 38.21 1.78 38.21 1.78 39.31 0.4 39.31 0.4 39.57 1.78 39.57 1.78 40.67 0.4 40.67 0.4 40.93 1.78 40.93 1.78 42.03 0.4 42.03 0.4 42.29 1.78 42.29 1.78 43.39 0.4 43.39 0.4 43.65 1.78 43.65 1.78 44.75 0.4 44.75 0.4 45.01 1.78 45.01 1.78 46.11 0.4 46.11 0.4 46.37 1.78 46.37 1.78 47.47 0.4 47.47 0.4 47.73 1.78 47.73 1.78 48.83 0.4 48.83 0.4 49.09 1.78 49.09 1.78 50.19 0.4 50.19 0.4 50.45 1.78 50.45 1.78 51.55 0.4 51.55 0.4 51.81 1.78 51.81 1.78 52.91 0.4 52.91 0.4 53.17 1.78 53.17 1.78 54.27 0.4 54.27 0.4 54.53 1.78 54.53 1.78 55.63 0.4 55.63 0.4 55.89 1.78 55.89 1.78 56.99 0.4 56.99 0.4 57.25 1.78 57.25 1.78 58.35 0.4 58.35 0.4 58.61 1.78 58.61 1.78 59.71 0.4 59.71 0.4 60.65 1.78 60.65 1.78 61.75 0.4 61.75 0.4 62.69 1.78 62.69 1.78 63.79 0.4 63.79 0.4 64.05 1.78 64.05 1.78 65.15 0.4 65.15 0.4 65.41 1.78 65.41 1.78 66.51 0.4 66.51 0.4 67.45 1.78 67.45 1.78 68.55 0.4 68.55 0.4 68.81 1.78 68.81 1.78 69.91 0.4 69.91 0.4 70.17 1.78 70.17 1.78 71.27 0.4 71.27 0.4 71.53 1.78 71.53 1.78 72.63 0.4 72.63 0.4 72.89 1.78 72.89 1.78 73.99 0.4 73.99 0.4 74.25 1.78 74.25 1.78 75.35 0.4 75.35 0.4 75.61 1.78 75.61 1.78 76.71 0.4 76.71 0.4 76.97 1.78 76.97 1.78 78.07 0.4 78.07 0.4 78.33 1.78 78.33 1.78 79.43 0.4 79.43 0.4 89.21 1.78 89.21 1.78 90.31 0.4 90.31 0.4 97.52 ;
    LAYER met2 ;
      RECT 80.82 97.735 81.1 98.105 ;
      RECT 51.38 97.735 51.66 98.105 ;
      RECT 10.9 97.735 11.18 98.105 ;
      RECT 15.51 12.42 15.77 12.74 ;
      RECT 10.9 10.695 11.18 11.065 ;
      RECT 56.91 1.54 57.17 1.86 ;
      RECT 51.85 1.54 52.11 1.86 ;
      RECT 48.17 1.54 48.43 1.86 ;
      RECT 80.82 -0.185 81.1 0.185 ;
      RECT 51.38 -0.185 51.66 0.185 ;
      POLYGON 91.72 97.64 91.72 0.28 82.23 0.28 82.23 1.64 81.53 1.64 81.53 0.28 74.87 0.28 74.87 1.64 74.17 1.64 74.17 0.28 73.95 0.28 73.95 1.64 73.25 1.64 73.25 0.28 73.03 0.28 73.03 1.64 72.33 1.64 72.33 0.28 72.11 0.28 72.11 1.64 71.41 1.64 71.41 0.28 71.19 0.28 71.19 1.64 70.49 1.64 70.49 0.28 69.81 0.28 69.81 1.64 69.11 1.64 69.11 0.28 68.89 0.28 68.89 1.64 68.19 1.64 68.19 0.28 67.51 0.28 67.51 1.64 66.81 1.64 66.81 0.28 66.59 0.28 66.59 1.64 65.89 1.64 65.89 0.28 65.21 0.28 65.21 1.64 64.51 1.64 64.51 0.28 64.29 0.28 64.29 1.64 63.59 1.64 63.59 0.28 63.37 0.28 63.37 1.64 62.67 1.64 62.67 0.28 62.45 0.28 62.45 1.64 61.75 1.64 61.75 0.28 61.53 0.28 61.53 1.64 60.83 1.64 60.83 0.28 60.61 0.28 60.61 1.64 59.91 1.64 59.91 0.28 59.23 0.28 59.23 1.64 58.53 1.64 58.53 0.28 57.85 0.28 57.85 1.64 57.15 1.64 57.15 0.28 56.93 0.28 56.93 1.64 56.23 1.64 56.23 0.28 56.01 0.28 56.01 1.64 55.31 1.64 55.31 0.28 54.63 0.28 54.63 1.64 53.93 1.64 53.93 0.28 53.71 0.28 53.71 1.64 53.01 1.64 53.01 0.28 52.79 0.28 52.79 1.64 52.09 1.64 52.09 0.28 50.95 0.28 50.95 1.64 50.25 1.64 50.25 0.28 49.57 0.28 49.57 1.64 48.87 1.64 48.87 0.28 48.19 0.28 48.19 1.64 47.49 1.64 47.49 0.28 47.27 0.28 47.27 1.64 46.57 1.64 46.57 0.28 45.89 0.28 45.89 1.64 45.19 1.64 45.19 0.28 44.51 0.28 44.51 1.64 43.81 1.64 43.81 0.28 43.13 0.28 43.13 1.64 42.43 1.64 42.43 0.28 42.21 0.28 42.21 1.64 41.51 1.64 41.51 0.28 41.29 0.28 41.29 1.64 40.59 1.64 40.59 0.28 40.37 0.28 40.37 1.64 39.67 1.64 39.67 0.28 39.45 0.28 39.45 1.64 38.75 1.64 38.75 0.28 38.53 0.28 38.53 1.64 37.83 1.64 37.83 0.28 37.61 0.28 37.61 1.64 36.91 1.64 36.91 0.28 34.39 0.28 34.39 1.64 33.69 1.64 33.69 0.28 32.55 0.28 32.55 1.64 31.85 1.64 31.85 0.28 31.63 0.28 31.63 1.64 30.93 1.64 30.93 0.28 28.41 0.28 28.41 1.64 27.71 1.64 27.71 0.28 26.04 0.28 26.04 11.16 18.75 11.16 18.75 12.52 18.05 12.52 18.05 11.16 16.45 11.16 16.45 12.52 15.75 12.52 15.75 11.16 15.53 11.16 15.53 12.52 14.83 12.52 14.83 11.16 13.23 11.16 13.23 12.52 12.53 12.52 12.53 11.16 12.31 11.16 12.31 12.52 11.61 12.52 11.61 11.16 10.47 11.16 10.47 12.52 9.77 12.52 9.77 11.16 9.55 11.16 9.55 12.52 8.85 12.52 8.85 11.16 8.63 11.16 8.63 12.52 7.93 12.52 7.93 11.16 7.71 11.16 7.71 12.52 7.01 12.52 7.01 11.16 6.79 11.16 6.79 12.52 6.09 12.52 6.09 11.16 5.41 11.16 5.41 12.52 4.71 12.52 4.71 11.16 4.49 11.16 4.49 12.52 3.79 12.52 3.79 11.16 0.28 11.16 0.28 97.64 1.95 97.64 1.95 96.28 2.65 96.28 2.65 97.64 30.93 97.64 30.93 96.28 31.63 96.28 31.63 97.64 ;
    LAYER met4 ;
      POLYGON 91.6 97.52 91.6 0.4 81.66 0.4 81.66 1 80.26 1 80.26 0.4 66.94 0.4 66.94 1 65.54 1 65.54 0.4 59.43 0.4 59.43 1.76 58.33 1.76 58.33 0.4 57.59 0.4 57.59 1.76 56.49 1.76 56.49 0.4 52.22 0.4 52.22 1 50.82 1 50.82 0.4 37.5 0.4 37.5 1 36.1 1 36.1 0.4 26.16 0.4 26.16 11.28 13.43 11.28 13.43 12.64 12.33 12.64 12.33 11.28 11.74 11.28 11.74 11.88 10.34 11.88 10.34 11.28 9.75 11.28 9.75 12.64 8.65 12.64 8.65 11.28 5.15 11.28 5.15 12.64 4.05 12.64 4.05 11.28 0.4 11.28 0.4 97.52 10.34 97.52 10.34 96.92 11.74 96.92 11.74 97.52 36.1 97.52 36.1 96.92 37.5 96.92 37.5 97.52 50.82 97.52 50.82 96.92 52.22 96.92 52.22 97.52 65.54 97.52 65.54 96.92 66.94 96.92 66.94 97.52 80.26 97.52 80.26 96.92 81.66 96.92 81.66 97.52 ;
    LAYER met5 ;
      POLYGON 90.4 96.32 90.4 88.2 87.2 88.2 87.2 81.8 90.4 81.8 90.4 67.8 87.2 67.8 87.2 61.4 90.4 61.4 90.4 47.4 87.2 47.4 87.2 41 90.4 41 90.4 27 87.2 27 87.2 20.6 90.4 20.6 90.4 1.6 27.36 1.6 27.36 12.48 1.6 12.48 1.6 20.6 4.8 20.6 4.8 27 1.6 27 1.6 41 4.8 41 4.8 47.4 1.6 47.4 1.6 61.4 4.8 61.4 4.8 67.8 1.6 67.8 1.6 81.8 4.8 81.8 4.8 88.2 1.6 88.2 1.6 96.32 ;
    LAYER met1 ;
      POLYGON 91.72 97.4 91.72 95.72 91.24 95.72 91.24 94.68 91.72 94.68 91.72 93 91.24 93 91.24 91.96 91.72 91.96 91.72 90.28 91.24 90.28 91.24 89.24 91.72 89.24 91.72 87.56 91.24 87.56 91.24 86.52 91.72 86.52 91.72 84.84 91.24 84.84 91.24 83.8 91.72 83.8 91.72 82.12 91.24 82.12 91.24 81.08 91.72 81.08 91.72 79.4 91.24 79.4 91.24 78.36 91.72 78.36 91.72 76.68 91.24 76.68 91.24 75.64 91.72 75.64 91.72 73.96 91.24 73.96 91.24 72.92 91.72 72.92 91.72 71.24 91.24 71.24 91.24 70.2 91.72 70.2 91.72 68.52 91.24 68.52 91.24 67.48 91.72 67.48 91.72 65.8 91.24 65.8 91.24 64.76 91.72 64.76 91.72 63.08 91.24 63.08 91.24 62.04 91.72 62.04 91.72 60.36 91.24 60.36 91.24 59.32 91.72 59.32 91.72 57.64 91.24 57.64 91.24 56.6 91.72 56.6 91.72 54.92 91.24 54.92 91.24 53.88 91.72 53.88 91.72 52.2 91.24 52.2 91.24 51.16 91.72 51.16 91.72 49.48 91.24 49.48 91.24 48.44 91.72 48.44 91.72 46.76 91.24 46.76 91.24 45.72 91.72 45.72 91.72 44.04 91.24 44.04 91.24 43 91.72 43 91.72 41.32 91.24 41.32 91.24 40.28 91.72 40.28 91.72 38.6 91.24 38.6 91.24 37.56 91.72 37.56 91.72 35.88 91.24 35.88 91.24 34.84 91.72 34.84 91.72 33.16 91.24 33.16 91.24 32.12 91.72 32.12 91.72 30.44 91.24 30.44 91.24 29.4 91.72 29.4 91.72 27.72 91.24 27.72 91.24 26.68 91.72 26.68 91.72 25 91.24 25 91.24 23.96 91.72 23.96 91.72 22.28 91.24 22.28 91.24 21.24 91.72 21.24 91.72 19.56 91.24 19.56 91.24 18.52 91.72 18.52 91.72 16.84 91.24 16.84 91.24 15.8 91.72 15.8 91.72 14.12 91.24 14.12 91.24 13.08 91.72 13.08 91.72 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 ;
      POLYGON 91.72 10.36 91.72 8.68 91.24 8.68 91.24 7.64 91.72 7.64 91.72 5.96 91.24 5.96 91.24 4.92 91.72 4.92 91.72 3.24 91.24 3.24 91.24 2.2 91.72 2.2 91.72 0.52 26.04 0.52 26.04 2.2 26.52 2.2 26.52 3.24 26.04 3.24 26.04 4.92 26.52 4.92 26.52 5.96 26.04 5.96 26.04 7.64 26.52 7.64 26.52 8.68 26.04 8.68 26.04 10.36 ;
    LAYER li1 ;
      POLYGON 91.83 97.75 91.83 0.17 25.93 0.17 25.93 11.05 0.17 11.05 0.17 97.75 ;
    LAYER mcon ;
      RECT 91.685 97.835 91.855 98.005 ;
      RECT 91.225 97.835 91.395 98.005 ;
      RECT 90.765 97.835 90.935 98.005 ;
      RECT 90.305 97.835 90.475 98.005 ;
      RECT 89.845 97.835 90.015 98.005 ;
      RECT 89.385 97.835 89.555 98.005 ;
      RECT 88.925 97.835 89.095 98.005 ;
      RECT 88.465 97.835 88.635 98.005 ;
      RECT 88.005 97.835 88.175 98.005 ;
      RECT 87.545 97.835 87.715 98.005 ;
      RECT 87.085 97.835 87.255 98.005 ;
      RECT 86.625 97.835 86.795 98.005 ;
      RECT 86.165 97.835 86.335 98.005 ;
      RECT 85.705 97.835 85.875 98.005 ;
      RECT 85.245 97.835 85.415 98.005 ;
      RECT 84.785 97.835 84.955 98.005 ;
      RECT 84.325 97.835 84.495 98.005 ;
      RECT 83.865 97.835 84.035 98.005 ;
      RECT 83.405 97.835 83.575 98.005 ;
      RECT 82.945 97.835 83.115 98.005 ;
      RECT 82.485 97.835 82.655 98.005 ;
      RECT 82.025 97.835 82.195 98.005 ;
      RECT 81.565 97.835 81.735 98.005 ;
      RECT 81.105 97.835 81.275 98.005 ;
      RECT 80.645 97.835 80.815 98.005 ;
      RECT 80.185 97.835 80.355 98.005 ;
      RECT 79.725 97.835 79.895 98.005 ;
      RECT 79.265 97.835 79.435 98.005 ;
      RECT 78.805 97.835 78.975 98.005 ;
      RECT 78.345 97.835 78.515 98.005 ;
      RECT 77.885 97.835 78.055 98.005 ;
      RECT 77.425 97.835 77.595 98.005 ;
      RECT 76.965 97.835 77.135 98.005 ;
      RECT 76.505 97.835 76.675 98.005 ;
      RECT 76.045 97.835 76.215 98.005 ;
      RECT 75.585 97.835 75.755 98.005 ;
      RECT 75.125 97.835 75.295 98.005 ;
      RECT 74.665 97.835 74.835 98.005 ;
      RECT 74.205 97.835 74.375 98.005 ;
      RECT 73.745 97.835 73.915 98.005 ;
      RECT 73.285 97.835 73.455 98.005 ;
      RECT 72.825 97.835 72.995 98.005 ;
      RECT 72.365 97.835 72.535 98.005 ;
      RECT 71.905 97.835 72.075 98.005 ;
      RECT 71.445 97.835 71.615 98.005 ;
      RECT 70.985 97.835 71.155 98.005 ;
      RECT 70.525 97.835 70.695 98.005 ;
      RECT 70.065 97.835 70.235 98.005 ;
      RECT 69.605 97.835 69.775 98.005 ;
      RECT 69.145 97.835 69.315 98.005 ;
      RECT 68.685 97.835 68.855 98.005 ;
      RECT 68.225 97.835 68.395 98.005 ;
      RECT 67.765 97.835 67.935 98.005 ;
      RECT 67.305 97.835 67.475 98.005 ;
      RECT 66.845 97.835 67.015 98.005 ;
      RECT 66.385 97.835 66.555 98.005 ;
      RECT 65.925 97.835 66.095 98.005 ;
      RECT 65.465 97.835 65.635 98.005 ;
      RECT 65.005 97.835 65.175 98.005 ;
      RECT 64.545 97.835 64.715 98.005 ;
      RECT 64.085 97.835 64.255 98.005 ;
      RECT 63.625 97.835 63.795 98.005 ;
      RECT 63.165 97.835 63.335 98.005 ;
      RECT 62.705 97.835 62.875 98.005 ;
      RECT 62.245 97.835 62.415 98.005 ;
      RECT 61.785 97.835 61.955 98.005 ;
      RECT 61.325 97.835 61.495 98.005 ;
      RECT 60.865 97.835 61.035 98.005 ;
      RECT 60.405 97.835 60.575 98.005 ;
      RECT 59.945 97.835 60.115 98.005 ;
      RECT 59.485 97.835 59.655 98.005 ;
      RECT 59.025 97.835 59.195 98.005 ;
      RECT 58.565 97.835 58.735 98.005 ;
      RECT 58.105 97.835 58.275 98.005 ;
      RECT 57.645 97.835 57.815 98.005 ;
      RECT 57.185 97.835 57.355 98.005 ;
      RECT 56.725 97.835 56.895 98.005 ;
      RECT 56.265 97.835 56.435 98.005 ;
      RECT 55.805 97.835 55.975 98.005 ;
      RECT 55.345 97.835 55.515 98.005 ;
      RECT 54.885 97.835 55.055 98.005 ;
      RECT 54.425 97.835 54.595 98.005 ;
      RECT 53.965 97.835 54.135 98.005 ;
      RECT 53.505 97.835 53.675 98.005 ;
      RECT 53.045 97.835 53.215 98.005 ;
      RECT 52.585 97.835 52.755 98.005 ;
      RECT 52.125 97.835 52.295 98.005 ;
      RECT 51.665 97.835 51.835 98.005 ;
      RECT 51.205 97.835 51.375 98.005 ;
      RECT 50.745 97.835 50.915 98.005 ;
      RECT 50.285 97.835 50.455 98.005 ;
      RECT 49.825 97.835 49.995 98.005 ;
      RECT 49.365 97.835 49.535 98.005 ;
      RECT 48.905 97.835 49.075 98.005 ;
      RECT 48.445 97.835 48.615 98.005 ;
      RECT 47.985 97.835 48.155 98.005 ;
      RECT 47.525 97.835 47.695 98.005 ;
      RECT 47.065 97.835 47.235 98.005 ;
      RECT 46.605 97.835 46.775 98.005 ;
      RECT 46.145 97.835 46.315 98.005 ;
      RECT 45.685 97.835 45.855 98.005 ;
      RECT 45.225 97.835 45.395 98.005 ;
      RECT 44.765 97.835 44.935 98.005 ;
      RECT 44.305 97.835 44.475 98.005 ;
      RECT 43.845 97.835 44.015 98.005 ;
      RECT 43.385 97.835 43.555 98.005 ;
      RECT 42.925 97.835 43.095 98.005 ;
      RECT 42.465 97.835 42.635 98.005 ;
      RECT 42.005 97.835 42.175 98.005 ;
      RECT 41.545 97.835 41.715 98.005 ;
      RECT 41.085 97.835 41.255 98.005 ;
      RECT 40.625 97.835 40.795 98.005 ;
      RECT 40.165 97.835 40.335 98.005 ;
      RECT 39.705 97.835 39.875 98.005 ;
      RECT 39.245 97.835 39.415 98.005 ;
      RECT 38.785 97.835 38.955 98.005 ;
      RECT 38.325 97.835 38.495 98.005 ;
      RECT 37.865 97.835 38.035 98.005 ;
      RECT 37.405 97.835 37.575 98.005 ;
      RECT 36.945 97.835 37.115 98.005 ;
      RECT 36.485 97.835 36.655 98.005 ;
      RECT 36.025 97.835 36.195 98.005 ;
      RECT 35.565 97.835 35.735 98.005 ;
      RECT 35.105 97.835 35.275 98.005 ;
      RECT 34.645 97.835 34.815 98.005 ;
      RECT 34.185 97.835 34.355 98.005 ;
      RECT 33.725 97.835 33.895 98.005 ;
      RECT 33.265 97.835 33.435 98.005 ;
      RECT 32.805 97.835 32.975 98.005 ;
      RECT 32.345 97.835 32.515 98.005 ;
      RECT 31.885 97.835 32.055 98.005 ;
      RECT 31.425 97.835 31.595 98.005 ;
      RECT 30.965 97.835 31.135 98.005 ;
      RECT 30.505 97.835 30.675 98.005 ;
      RECT 30.045 97.835 30.215 98.005 ;
      RECT 29.585 97.835 29.755 98.005 ;
      RECT 29.125 97.835 29.295 98.005 ;
      RECT 28.665 97.835 28.835 98.005 ;
      RECT 28.205 97.835 28.375 98.005 ;
      RECT 27.745 97.835 27.915 98.005 ;
      RECT 27.285 97.835 27.455 98.005 ;
      RECT 26.825 97.835 26.995 98.005 ;
      RECT 26.365 97.835 26.535 98.005 ;
      RECT 25.905 97.835 26.075 98.005 ;
      RECT 25.445 97.835 25.615 98.005 ;
      RECT 24.985 97.835 25.155 98.005 ;
      RECT 24.525 97.835 24.695 98.005 ;
      RECT 24.065 97.835 24.235 98.005 ;
      RECT 23.605 97.835 23.775 98.005 ;
      RECT 23.145 97.835 23.315 98.005 ;
      RECT 22.685 97.835 22.855 98.005 ;
      RECT 22.225 97.835 22.395 98.005 ;
      RECT 21.765 97.835 21.935 98.005 ;
      RECT 21.305 97.835 21.475 98.005 ;
      RECT 20.845 97.835 21.015 98.005 ;
      RECT 20.385 97.835 20.555 98.005 ;
      RECT 19.925 97.835 20.095 98.005 ;
      RECT 19.465 97.835 19.635 98.005 ;
      RECT 19.005 97.835 19.175 98.005 ;
      RECT 18.545 97.835 18.715 98.005 ;
      RECT 18.085 97.835 18.255 98.005 ;
      RECT 17.625 97.835 17.795 98.005 ;
      RECT 17.165 97.835 17.335 98.005 ;
      RECT 16.705 97.835 16.875 98.005 ;
      RECT 16.245 97.835 16.415 98.005 ;
      RECT 15.785 97.835 15.955 98.005 ;
      RECT 15.325 97.835 15.495 98.005 ;
      RECT 14.865 97.835 15.035 98.005 ;
      RECT 14.405 97.835 14.575 98.005 ;
      RECT 13.945 97.835 14.115 98.005 ;
      RECT 13.485 97.835 13.655 98.005 ;
      RECT 13.025 97.835 13.195 98.005 ;
      RECT 12.565 97.835 12.735 98.005 ;
      RECT 12.105 97.835 12.275 98.005 ;
      RECT 11.645 97.835 11.815 98.005 ;
      RECT 11.185 97.835 11.355 98.005 ;
      RECT 10.725 97.835 10.895 98.005 ;
      RECT 10.265 97.835 10.435 98.005 ;
      RECT 9.805 97.835 9.975 98.005 ;
      RECT 9.345 97.835 9.515 98.005 ;
      RECT 8.885 97.835 9.055 98.005 ;
      RECT 8.425 97.835 8.595 98.005 ;
      RECT 7.965 97.835 8.135 98.005 ;
      RECT 7.505 97.835 7.675 98.005 ;
      RECT 7.045 97.835 7.215 98.005 ;
      RECT 6.585 97.835 6.755 98.005 ;
      RECT 6.125 97.835 6.295 98.005 ;
      RECT 5.665 97.835 5.835 98.005 ;
      RECT 5.205 97.835 5.375 98.005 ;
      RECT 4.745 97.835 4.915 98.005 ;
      RECT 4.285 97.835 4.455 98.005 ;
      RECT 3.825 97.835 3.995 98.005 ;
      RECT 3.365 97.835 3.535 98.005 ;
      RECT 2.905 97.835 3.075 98.005 ;
      RECT 2.445 97.835 2.615 98.005 ;
      RECT 1.985 97.835 2.155 98.005 ;
      RECT 1.525 97.835 1.695 98.005 ;
      RECT 1.065 97.835 1.235 98.005 ;
      RECT 0.605 97.835 0.775 98.005 ;
      RECT 0.145 97.835 0.315 98.005 ;
      RECT 91.685 95.115 91.855 95.285 ;
      RECT 91.225 95.115 91.395 95.285 ;
      RECT 0.605 95.115 0.775 95.285 ;
      RECT 0.145 95.115 0.315 95.285 ;
      RECT 91.685 92.395 91.855 92.565 ;
      RECT 91.225 92.395 91.395 92.565 ;
      RECT 0.605 92.395 0.775 92.565 ;
      RECT 0.145 92.395 0.315 92.565 ;
      RECT 91.685 89.675 91.855 89.845 ;
      RECT 91.225 89.675 91.395 89.845 ;
      RECT 0.605 89.675 0.775 89.845 ;
      RECT 0.145 89.675 0.315 89.845 ;
      RECT 91.685 86.955 91.855 87.125 ;
      RECT 91.225 86.955 91.395 87.125 ;
      RECT 0.605 86.955 0.775 87.125 ;
      RECT 0.145 86.955 0.315 87.125 ;
      RECT 91.685 84.235 91.855 84.405 ;
      RECT 91.225 84.235 91.395 84.405 ;
      RECT 0.605 84.235 0.775 84.405 ;
      RECT 0.145 84.235 0.315 84.405 ;
      RECT 91.685 81.515 91.855 81.685 ;
      RECT 91.225 81.515 91.395 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 91.685 78.795 91.855 78.965 ;
      RECT 91.225 78.795 91.395 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 91.685 76.075 91.855 76.245 ;
      RECT 91.225 76.075 91.395 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 91.685 73.355 91.855 73.525 ;
      RECT 91.225 73.355 91.395 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 91.685 70.635 91.855 70.805 ;
      RECT 91.225 70.635 91.395 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 91.685 67.915 91.855 68.085 ;
      RECT 91.225 67.915 91.395 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 91.685 65.195 91.855 65.365 ;
      RECT 91.225 65.195 91.395 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 91.685 62.475 91.855 62.645 ;
      RECT 91.225 62.475 91.395 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 91.685 59.755 91.855 59.925 ;
      RECT 91.225 59.755 91.395 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 91.685 57.035 91.855 57.205 ;
      RECT 91.225 57.035 91.395 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 91.685 54.315 91.855 54.485 ;
      RECT 91.225 54.315 91.395 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 91.685 51.595 91.855 51.765 ;
      RECT 91.225 51.595 91.395 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 91.685 48.875 91.855 49.045 ;
      RECT 91.225 48.875 91.395 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 91.685 46.155 91.855 46.325 ;
      RECT 91.225 46.155 91.395 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 91.685 43.435 91.855 43.605 ;
      RECT 91.225 43.435 91.395 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 91.685 40.715 91.855 40.885 ;
      RECT 91.225 40.715 91.395 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 91.685 37.995 91.855 38.165 ;
      RECT 91.225 37.995 91.395 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 91.685 35.275 91.855 35.445 ;
      RECT 91.225 35.275 91.395 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 91.685 32.555 91.855 32.725 ;
      RECT 91.225 32.555 91.395 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 91.685 29.835 91.855 30.005 ;
      RECT 91.225 29.835 91.395 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 91.685 27.115 91.855 27.285 ;
      RECT 91.225 27.115 91.395 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 91.685 24.395 91.855 24.565 ;
      RECT 91.225 24.395 91.395 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 91.685 21.675 91.855 21.845 ;
      RECT 91.225 21.675 91.395 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 91.685 18.955 91.855 19.125 ;
      RECT 91.225 18.955 91.395 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 91.685 16.235 91.855 16.405 ;
      RECT 91.225 16.235 91.395 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 91.685 13.515 91.855 13.685 ;
      RECT 91.225 13.515 91.395 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 91.685 10.795 91.855 10.965 ;
      RECT 91.225 10.795 91.395 10.965 ;
      RECT 90.765 10.795 90.935 10.965 ;
      RECT 90.305 10.795 90.475 10.965 ;
      RECT 89.845 10.795 90.015 10.965 ;
      RECT 89.385 10.795 89.555 10.965 ;
      RECT 88.925 10.795 89.095 10.965 ;
      RECT 88.465 10.795 88.635 10.965 ;
      RECT 88.005 10.795 88.175 10.965 ;
      RECT 87.545 10.795 87.715 10.965 ;
      RECT 87.085 10.795 87.255 10.965 ;
      RECT 86.625 10.795 86.795 10.965 ;
      RECT 86.165 10.795 86.335 10.965 ;
      RECT 85.705 10.795 85.875 10.965 ;
      RECT 85.245 10.795 85.415 10.965 ;
      RECT 84.785 10.795 84.955 10.965 ;
      RECT 84.325 10.795 84.495 10.965 ;
      RECT 83.865 10.795 84.035 10.965 ;
      RECT 83.405 10.795 83.575 10.965 ;
      RECT 82.945 10.795 83.115 10.965 ;
      RECT 82.485 10.795 82.655 10.965 ;
      RECT 82.025 10.795 82.195 10.965 ;
      RECT 81.565 10.795 81.735 10.965 ;
      RECT 81.105 10.795 81.275 10.965 ;
      RECT 80.645 10.795 80.815 10.965 ;
      RECT 80.185 10.795 80.355 10.965 ;
      RECT 79.725 10.795 79.895 10.965 ;
      RECT 79.265 10.795 79.435 10.965 ;
      RECT 78.805 10.795 78.975 10.965 ;
      RECT 78.345 10.795 78.515 10.965 ;
      RECT 77.885 10.795 78.055 10.965 ;
      RECT 77.425 10.795 77.595 10.965 ;
      RECT 76.965 10.795 77.135 10.965 ;
      RECT 76.505 10.795 76.675 10.965 ;
      RECT 76.045 10.795 76.215 10.965 ;
      RECT 75.585 10.795 75.755 10.965 ;
      RECT 75.125 10.795 75.295 10.965 ;
      RECT 74.665 10.795 74.835 10.965 ;
      RECT 74.205 10.795 74.375 10.965 ;
      RECT 73.745 10.795 73.915 10.965 ;
      RECT 73.285 10.795 73.455 10.965 ;
      RECT 72.825 10.795 72.995 10.965 ;
      RECT 72.365 10.795 72.535 10.965 ;
      RECT 71.905 10.795 72.075 10.965 ;
      RECT 71.445 10.795 71.615 10.965 ;
      RECT 70.985 10.795 71.155 10.965 ;
      RECT 70.525 10.795 70.695 10.965 ;
      RECT 70.065 10.795 70.235 10.965 ;
      RECT 69.605 10.795 69.775 10.965 ;
      RECT 69.145 10.795 69.315 10.965 ;
      RECT 68.685 10.795 68.855 10.965 ;
      RECT 68.225 10.795 68.395 10.965 ;
      RECT 67.765 10.795 67.935 10.965 ;
      RECT 67.305 10.795 67.475 10.965 ;
      RECT 66.845 10.795 67.015 10.965 ;
      RECT 66.385 10.795 66.555 10.965 ;
      RECT 65.925 10.795 66.095 10.965 ;
      RECT 65.465 10.795 65.635 10.965 ;
      RECT 65.005 10.795 65.175 10.965 ;
      RECT 64.545 10.795 64.715 10.965 ;
      RECT 64.085 10.795 64.255 10.965 ;
      RECT 63.625 10.795 63.795 10.965 ;
      RECT 63.165 10.795 63.335 10.965 ;
      RECT 62.705 10.795 62.875 10.965 ;
      RECT 62.245 10.795 62.415 10.965 ;
      RECT 61.785 10.795 61.955 10.965 ;
      RECT 61.325 10.795 61.495 10.965 ;
      RECT 60.865 10.795 61.035 10.965 ;
      RECT 60.405 10.795 60.575 10.965 ;
      RECT 59.945 10.795 60.115 10.965 ;
      RECT 59.485 10.795 59.655 10.965 ;
      RECT 59.025 10.795 59.195 10.965 ;
      RECT 58.565 10.795 58.735 10.965 ;
      RECT 58.105 10.795 58.275 10.965 ;
      RECT 57.645 10.795 57.815 10.965 ;
      RECT 57.185 10.795 57.355 10.965 ;
      RECT 56.725 10.795 56.895 10.965 ;
      RECT 56.265 10.795 56.435 10.965 ;
      RECT 55.805 10.795 55.975 10.965 ;
      RECT 55.345 10.795 55.515 10.965 ;
      RECT 54.885 10.795 55.055 10.965 ;
      RECT 54.425 10.795 54.595 10.965 ;
      RECT 53.965 10.795 54.135 10.965 ;
      RECT 53.505 10.795 53.675 10.965 ;
      RECT 53.045 10.795 53.215 10.965 ;
      RECT 52.585 10.795 52.755 10.965 ;
      RECT 52.125 10.795 52.295 10.965 ;
      RECT 51.665 10.795 51.835 10.965 ;
      RECT 51.205 10.795 51.375 10.965 ;
      RECT 50.745 10.795 50.915 10.965 ;
      RECT 50.285 10.795 50.455 10.965 ;
      RECT 49.825 10.795 49.995 10.965 ;
      RECT 49.365 10.795 49.535 10.965 ;
      RECT 48.905 10.795 49.075 10.965 ;
      RECT 48.445 10.795 48.615 10.965 ;
      RECT 47.985 10.795 48.155 10.965 ;
      RECT 47.525 10.795 47.695 10.965 ;
      RECT 47.065 10.795 47.235 10.965 ;
      RECT 46.605 10.795 46.775 10.965 ;
      RECT 46.145 10.795 46.315 10.965 ;
      RECT 45.685 10.795 45.855 10.965 ;
      RECT 45.225 10.795 45.395 10.965 ;
      RECT 44.765 10.795 44.935 10.965 ;
      RECT 44.305 10.795 44.475 10.965 ;
      RECT 43.845 10.795 44.015 10.965 ;
      RECT 43.385 10.795 43.555 10.965 ;
      RECT 42.925 10.795 43.095 10.965 ;
      RECT 42.465 10.795 42.635 10.965 ;
      RECT 42.005 10.795 42.175 10.965 ;
      RECT 41.545 10.795 41.715 10.965 ;
      RECT 41.085 10.795 41.255 10.965 ;
      RECT 40.625 10.795 40.795 10.965 ;
      RECT 40.165 10.795 40.335 10.965 ;
      RECT 39.705 10.795 39.875 10.965 ;
      RECT 39.245 10.795 39.415 10.965 ;
      RECT 38.785 10.795 38.955 10.965 ;
      RECT 38.325 10.795 38.495 10.965 ;
      RECT 37.865 10.795 38.035 10.965 ;
      RECT 37.405 10.795 37.575 10.965 ;
      RECT 36.945 10.795 37.115 10.965 ;
      RECT 36.485 10.795 36.655 10.965 ;
      RECT 36.025 10.795 36.195 10.965 ;
      RECT 35.565 10.795 35.735 10.965 ;
      RECT 35.105 10.795 35.275 10.965 ;
      RECT 34.645 10.795 34.815 10.965 ;
      RECT 34.185 10.795 34.355 10.965 ;
      RECT 33.725 10.795 33.895 10.965 ;
      RECT 33.265 10.795 33.435 10.965 ;
      RECT 32.805 10.795 32.975 10.965 ;
      RECT 32.345 10.795 32.515 10.965 ;
      RECT 31.885 10.795 32.055 10.965 ;
      RECT 31.425 10.795 31.595 10.965 ;
      RECT 30.965 10.795 31.135 10.965 ;
      RECT 30.505 10.795 30.675 10.965 ;
      RECT 30.045 10.795 30.215 10.965 ;
      RECT 29.585 10.795 29.755 10.965 ;
      RECT 29.125 10.795 29.295 10.965 ;
      RECT 28.665 10.795 28.835 10.965 ;
      RECT 28.205 10.795 28.375 10.965 ;
      RECT 27.745 10.795 27.915 10.965 ;
      RECT 27.285 10.795 27.455 10.965 ;
      RECT 26.825 10.795 26.995 10.965 ;
      RECT 26.365 10.795 26.535 10.965 ;
      RECT 25.905 10.795 26.075 10.965 ;
      RECT 25.445 10.795 25.615 10.965 ;
      RECT 24.985 10.795 25.155 10.965 ;
      RECT 24.525 10.795 24.695 10.965 ;
      RECT 24.065 10.795 24.235 10.965 ;
      RECT 23.605 10.795 23.775 10.965 ;
      RECT 23.145 10.795 23.315 10.965 ;
      RECT 22.685 10.795 22.855 10.965 ;
      RECT 22.225 10.795 22.395 10.965 ;
      RECT 21.765 10.795 21.935 10.965 ;
      RECT 21.305 10.795 21.475 10.965 ;
      RECT 20.845 10.795 21.015 10.965 ;
      RECT 20.385 10.795 20.555 10.965 ;
      RECT 19.925 10.795 20.095 10.965 ;
      RECT 19.465 10.795 19.635 10.965 ;
      RECT 19.005 10.795 19.175 10.965 ;
      RECT 18.545 10.795 18.715 10.965 ;
      RECT 18.085 10.795 18.255 10.965 ;
      RECT 17.625 10.795 17.795 10.965 ;
      RECT 17.165 10.795 17.335 10.965 ;
      RECT 16.705 10.795 16.875 10.965 ;
      RECT 16.245 10.795 16.415 10.965 ;
      RECT 15.785 10.795 15.955 10.965 ;
      RECT 15.325 10.795 15.495 10.965 ;
      RECT 14.865 10.795 15.035 10.965 ;
      RECT 14.405 10.795 14.575 10.965 ;
      RECT 13.945 10.795 14.115 10.965 ;
      RECT 13.485 10.795 13.655 10.965 ;
      RECT 13.025 10.795 13.195 10.965 ;
      RECT 12.565 10.795 12.735 10.965 ;
      RECT 12.105 10.795 12.275 10.965 ;
      RECT 11.645 10.795 11.815 10.965 ;
      RECT 11.185 10.795 11.355 10.965 ;
      RECT 10.725 10.795 10.895 10.965 ;
      RECT 10.265 10.795 10.435 10.965 ;
      RECT 9.805 10.795 9.975 10.965 ;
      RECT 9.345 10.795 9.515 10.965 ;
      RECT 8.885 10.795 9.055 10.965 ;
      RECT 8.425 10.795 8.595 10.965 ;
      RECT 7.965 10.795 8.135 10.965 ;
      RECT 7.505 10.795 7.675 10.965 ;
      RECT 7.045 10.795 7.215 10.965 ;
      RECT 6.585 10.795 6.755 10.965 ;
      RECT 6.125 10.795 6.295 10.965 ;
      RECT 5.665 10.795 5.835 10.965 ;
      RECT 5.205 10.795 5.375 10.965 ;
      RECT 4.745 10.795 4.915 10.965 ;
      RECT 4.285 10.795 4.455 10.965 ;
      RECT 3.825 10.795 3.995 10.965 ;
      RECT 3.365 10.795 3.535 10.965 ;
      RECT 2.905 10.795 3.075 10.965 ;
      RECT 2.445 10.795 2.615 10.965 ;
      RECT 1.985 10.795 2.155 10.965 ;
      RECT 1.525 10.795 1.695 10.965 ;
      RECT 1.065 10.795 1.235 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 91.685 8.075 91.855 8.245 ;
      RECT 91.225 8.075 91.395 8.245 ;
      RECT 26.365 8.075 26.535 8.245 ;
      RECT 25.905 8.075 26.075 8.245 ;
      RECT 91.685 5.355 91.855 5.525 ;
      RECT 91.225 5.355 91.395 5.525 ;
      RECT 26.365 5.355 26.535 5.525 ;
      RECT 25.905 5.355 26.075 5.525 ;
      RECT 91.685 2.635 91.855 2.805 ;
      RECT 91.225 2.635 91.395 2.805 ;
      RECT 26.365 2.635 26.535 2.805 ;
      RECT 25.905 2.635 26.075 2.805 ;
      RECT 91.685 -0.085 91.855 0.085 ;
      RECT 91.225 -0.085 91.395 0.085 ;
      RECT 90.765 -0.085 90.935 0.085 ;
      RECT 90.305 -0.085 90.475 0.085 ;
      RECT 89.845 -0.085 90.015 0.085 ;
      RECT 89.385 -0.085 89.555 0.085 ;
      RECT 88.925 -0.085 89.095 0.085 ;
      RECT 88.465 -0.085 88.635 0.085 ;
      RECT 88.005 -0.085 88.175 0.085 ;
      RECT 87.545 -0.085 87.715 0.085 ;
      RECT 87.085 -0.085 87.255 0.085 ;
      RECT 86.625 -0.085 86.795 0.085 ;
      RECT 86.165 -0.085 86.335 0.085 ;
      RECT 85.705 -0.085 85.875 0.085 ;
      RECT 85.245 -0.085 85.415 0.085 ;
      RECT 84.785 -0.085 84.955 0.085 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
    LAYER via ;
      RECT 80.885 97.845 81.035 97.995 ;
      RECT 51.445 97.845 51.595 97.995 ;
      RECT 10.965 97.845 11.115 97.995 ;
      RECT 31.205 96.145 31.355 96.295 ;
      RECT 9.125 12.505 9.275 12.655 ;
      RECT 80.885 10.805 81.035 10.955 ;
      RECT 51.445 10.805 51.595 10.955 ;
      RECT 10.965 10.805 11.115 10.955 ;
      RECT 52.365 1.625 52.515 1.775 ;
      RECT 49.145 1.625 49.295 1.775 ;
      RECT 45.465 1.625 45.615 1.775 ;
      RECT 39.945 1.625 40.095 1.775 ;
      RECT 80.885 -0.075 81.035 0.075 ;
      RECT 51.445 -0.075 51.595 0.075 ;
    LAYER via2 ;
      RECT 80.86 97.82 81.06 98.02 ;
      RECT 51.42 97.82 51.62 98.02 ;
      RECT 10.94 97.82 11.14 98.02 ;
      RECT 1.28 78.78 1.48 78.98 ;
      RECT 1.74 70.62 1.94 70.82 ;
      RECT 1.28 37.3 1.48 37.5 ;
      RECT 1.28 33.22 1.48 33.42 ;
      RECT 1.28 16.22 1.48 16.42 ;
      RECT 1.28 14.86 1.48 15.06 ;
      RECT 10.94 10.78 11.14 10.98 ;
      RECT 80.86 -0.1 81.06 0.1 ;
      RECT 51.42 -0.1 51.62 0.1 ;
    LAYER via3 ;
      RECT 80.86 97.82 81.06 98.02 ;
      RECT 51.42 97.82 51.62 98.02 ;
      RECT 10.94 97.82 11.14 98.02 ;
      RECT 1.74 59.06 1.94 59.26 ;
      RECT 10.94 10.78 11.14 10.98 ;
      RECT 80.86 -0.1 81.06 0.1 ;
      RECT 51.42 -0.1 51.62 0.1 ;
    LAYER OVERLAP ;
      POLYGON 25.76 0 25.76 10.88 0 10.88 0 97.92 92 97.92 92 0 ;
  END
END sb_2__2_

END LIBRARY
