//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module fpga_top
(
    ccff_head,
    clk,
    gfpga_pad_io_soc_in,
    isol_n,
    prog_clk,
    prog_reset,
    reset,
    scan_enable,
    ccff_tail,
    gfpga_pad_io_soc_dir,
    gfpga_pad_io_soc_out
);

    input ccff_head;
    input clk;
    input [0:127]gfpga_pad_io_soc_in;
    input isol_n;
    input prog_clk;
    input prog_reset;
    input reset;
    input scan_enable;
    output ccff_tail;
    output [0:127]gfpga_pad_io_soc_dir;
    output [0:127]gfpga_pad_io_soc_out;

    wire cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__0__0_ccff_tail;
    wire [0:29]cbx_1__0__0_chanx_left_out;
    wire [0:29]cbx_1__0__0_chanx_right_out;
    wire cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__0__1_ccff_tail;
    wire [0:29]cbx_1__0__1_chanx_left_out;
    wire [0:29]cbx_1__0__1_chanx_right_out;
    wire cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__0__2_ccff_tail;
    wire [0:29]cbx_1__0__2_chanx_left_out;
    wire [0:29]cbx_1__0__2_chanx_right_out;
    wire cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__0__3_ccff_tail;
    wire [0:29]cbx_1__0__3_chanx_left_out;
    wire [0:29]cbx_1__0__3_chanx_right_out;
    wire cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__0__4_ccff_tail;
    wire [0:29]cbx_1__0__4_chanx_left_out;
    wire [0:29]cbx_1__0__4_chanx_right_out;
    wire cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__0__5_ccff_tail;
    wire [0:29]cbx_1__0__5_chanx_left_out;
    wire [0:29]cbx_1__0__5_chanx_right_out;
    wire cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__0__6_ccff_tail;
    wire [0:29]cbx_1__0__6_chanx_left_out;
    wire [0:29]cbx_1__0__6_chanx_right_out;
    wire cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__0__7_ccff_tail;
    wire [0:29]cbx_1__0__7_chanx_left_out;
    wire [0:29]cbx_1__0__7_chanx_right_out;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__0_ccff_tail;
    wire [0:29]cbx_1__1__0_chanx_left_out;
    wire [0:29]cbx_1__1__0_chanx_right_out;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__10_ccff_tail;
    wire [0:29]cbx_1__1__10_chanx_left_out;
    wire [0:29]cbx_1__1__10_chanx_right_out;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__11_ccff_tail;
    wire [0:29]cbx_1__1__11_chanx_left_out;
    wire [0:29]cbx_1__1__11_chanx_right_out;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__12_ccff_tail;
    wire [0:29]cbx_1__1__12_chanx_left_out;
    wire [0:29]cbx_1__1__12_chanx_right_out;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__13_ccff_tail;
    wire [0:29]cbx_1__1__13_chanx_left_out;
    wire [0:29]cbx_1__1__13_chanx_right_out;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__14_ccff_tail;
    wire [0:29]cbx_1__1__14_chanx_left_out;
    wire [0:29]cbx_1__1__14_chanx_right_out;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__15_ccff_tail;
    wire [0:29]cbx_1__1__15_chanx_left_out;
    wire [0:29]cbx_1__1__15_chanx_right_out;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__16_ccff_tail;
    wire [0:29]cbx_1__1__16_chanx_left_out;
    wire [0:29]cbx_1__1__16_chanx_right_out;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__17_ccff_tail;
    wire [0:29]cbx_1__1__17_chanx_left_out;
    wire [0:29]cbx_1__1__17_chanx_right_out;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__18_ccff_tail;
    wire [0:29]cbx_1__1__18_chanx_left_out;
    wire [0:29]cbx_1__1__18_chanx_right_out;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__19_ccff_tail;
    wire [0:29]cbx_1__1__19_chanx_left_out;
    wire [0:29]cbx_1__1__19_chanx_right_out;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__1_ccff_tail;
    wire [0:29]cbx_1__1__1_chanx_left_out;
    wire [0:29]cbx_1__1__1_chanx_right_out;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__20_ccff_tail;
    wire [0:29]cbx_1__1__20_chanx_left_out;
    wire [0:29]cbx_1__1__20_chanx_right_out;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__21_ccff_tail;
    wire [0:29]cbx_1__1__21_chanx_left_out;
    wire [0:29]cbx_1__1__21_chanx_right_out;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__22_ccff_tail;
    wire [0:29]cbx_1__1__22_chanx_left_out;
    wire [0:29]cbx_1__1__22_chanx_right_out;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__23_ccff_tail;
    wire [0:29]cbx_1__1__23_chanx_left_out;
    wire [0:29]cbx_1__1__23_chanx_right_out;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__24_ccff_tail;
    wire [0:29]cbx_1__1__24_chanx_left_out;
    wire [0:29]cbx_1__1__24_chanx_right_out;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__25_ccff_tail;
    wire [0:29]cbx_1__1__25_chanx_left_out;
    wire [0:29]cbx_1__1__25_chanx_right_out;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__26_ccff_tail;
    wire [0:29]cbx_1__1__26_chanx_left_out;
    wire [0:29]cbx_1__1__26_chanx_right_out;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__27_ccff_tail;
    wire [0:29]cbx_1__1__27_chanx_left_out;
    wire [0:29]cbx_1__1__27_chanx_right_out;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__28_ccff_tail;
    wire [0:29]cbx_1__1__28_chanx_left_out;
    wire [0:29]cbx_1__1__28_chanx_right_out;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__29_ccff_tail;
    wire [0:29]cbx_1__1__29_chanx_left_out;
    wire [0:29]cbx_1__1__29_chanx_right_out;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__2_ccff_tail;
    wire [0:29]cbx_1__1__2_chanx_left_out;
    wire [0:29]cbx_1__1__2_chanx_right_out;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__30_ccff_tail;
    wire [0:29]cbx_1__1__30_chanx_left_out;
    wire [0:29]cbx_1__1__30_chanx_right_out;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__31_ccff_tail;
    wire [0:29]cbx_1__1__31_chanx_left_out;
    wire [0:29]cbx_1__1__31_chanx_right_out;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__32_ccff_tail;
    wire [0:29]cbx_1__1__32_chanx_left_out;
    wire [0:29]cbx_1__1__32_chanx_right_out;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__33_ccff_tail;
    wire [0:29]cbx_1__1__33_chanx_left_out;
    wire [0:29]cbx_1__1__33_chanx_right_out;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__34_ccff_tail;
    wire [0:29]cbx_1__1__34_chanx_left_out;
    wire [0:29]cbx_1__1__34_chanx_right_out;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__35_ccff_tail;
    wire [0:29]cbx_1__1__35_chanx_left_out;
    wire [0:29]cbx_1__1__35_chanx_right_out;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__36_ccff_tail;
    wire [0:29]cbx_1__1__36_chanx_left_out;
    wire [0:29]cbx_1__1__36_chanx_right_out;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__37_ccff_tail;
    wire [0:29]cbx_1__1__37_chanx_left_out;
    wire [0:29]cbx_1__1__37_chanx_right_out;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__38_ccff_tail;
    wire [0:29]cbx_1__1__38_chanx_left_out;
    wire [0:29]cbx_1__1__38_chanx_right_out;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__39_ccff_tail;
    wire [0:29]cbx_1__1__39_chanx_left_out;
    wire [0:29]cbx_1__1__39_chanx_right_out;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__3_ccff_tail;
    wire [0:29]cbx_1__1__3_chanx_left_out;
    wire [0:29]cbx_1__1__3_chanx_right_out;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__40_ccff_tail;
    wire [0:29]cbx_1__1__40_chanx_left_out;
    wire [0:29]cbx_1__1__40_chanx_right_out;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__41_ccff_tail;
    wire [0:29]cbx_1__1__41_chanx_left_out;
    wire [0:29]cbx_1__1__41_chanx_right_out;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__42_ccff_tail;
    wire [0:29]cbx_1__1__42_chanx_left_out;
    wire [0:29]cbx_1__1__42_chanx_right_out;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__43_ccff_tail;
    wire [0:29]cbx_1__1__43_chanx_left_out;
    wire [0:29]cbx_1__1__43_chanx_right_out;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__44_ccff_tail;
    wire [0:29]cbx_1__1__44_chanx_left_out;
    wire [0:29]cbx_1__1__44_chanx_right_out;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__45_ccff_tail;
    wire [0:29]cbx_1__1__45_chanx_left_out;
    wire [0:29]cbx_1__1__45_chanx_right_out;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__46_ccff_tail;
    wire [0:29]cbx_1__1__46_chanx_left_out;
    wire [0:29]cbx_1__1__46_chanx_right_out;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__47_ccff_tail;
    wire [0:29]cbx_1__1__47_chanx_left_out;
    wire [0:29]cbx_1__1__47_chanx_right_out;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__48_ccff_tail;
    wire [0:29]cbx_1__1__48_chanx_left_out;
    wire [0:29]cbx_1__1__48_chanx_right_out;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__49_ccff_tail;
    wire [0:29]cbx_1__1__49_chanx_left_out;
    wire [0:29]cbx_1__1__49_chanx_right_out;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__4_ccff_tail;
    wire [0:29]cbx_1__1__4_chanx_left_out;
    wire [0:29]cbx_1__1__4_chanx_right_out;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__50_ccff_tail;
    wire [0:29]cbx_1__1__50_chanx_left_out;
    wire [0:29]cbx_1__1__50_chanx_right_out;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__51_ccff_tail;
    wire [0:29]cbx_1__1__51_chanx_left_out;
    wire [0:29]cbx_1__1__51_chanx_right_out;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__52_ccff_tail;
    wire [0:29]cbx_1__1__52_chanx_left_out;
    wire [0:29]cbx_1__1__52_chanx_right_out;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__53_ccff_tail;
    wire [0:29]cbx_1__1__53_chanx_left_out;
    wire [0:29]cbx_1__1__53_chanx_right_out;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__54_ccff_tail;
    wire [0:29]cbx_1__1__54_chanx_left_out;
    wire [0:29]cbx_1__1__54_chanx_right_out;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__55_ccff_tail;
    wire [0:29]cbx_1__1__55_chanx_left_out;
    wire [0:29]cbx_1__1__55_chanx_right_out;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__5_ccff_tail;
    wire [0:29]cbx_1__1__5_chanx_left_out;
    wire [0:29]cbx_1__1__5_chanx_right_out;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__6_ccff_tail;
    wire [0:29]cbx_1__1__6_chanx_left_out;
    wire [0:29]cbx_1__1__6_chanx_right_out;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__7_ccff_tail;
    wire [0:29]cbx_1__1__7_chanx_left_out;
    wire [0:29]cbx_1__1__7_chanx_right_out;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__8_ccff_tail;
    wire [0:29]cbx_1__1__8_chanx_left_out;
    wire [0:29]cbx_1__1__8_chanx_right_out;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__1__9_ccff_tail;
    wire [0:29]cbx_1__1__9_chanx_left_out;
    wire [0:29]cbx_1__1__9_chanx_right_out;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__8__0_ccff_tail;
    wire [0:29]cbx_1__8__0_chanx_left_out;
    wire [0:29]cbx_1__8__0_chanx_right_out;
    wire cbx_1__8__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__8__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__8__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__8__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__8__1_ccff_tail;
    wire [0:29]cbx_1__8__1_chanx_left_out;
    wire [0:29]cbx_1__8__1_chanx_right_out;
    wire cbx_1__8__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__8__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__8__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__8__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__8__2_ccff_tail;
    wire [0:29]cbx_1__8__2_chanx_left_out;
    wire [0:29]cbx_1__8__2_chanx_right_out;
    wire cbx_1__8__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__8__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__8__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__8__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__8__3_ccff_tail;
    wire [0:29]cbx_1__8__3_chanx_left_out;
    wire [0:29]cbx_1__8__3_chanx_right_out;
    wire cbx_1__8__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__8__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__8__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__8__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__8__4_ccff_tail;
    wire [0:29]cbx_1__8__4_chanx_left_out;
    wire [0:29]cbx_1__8__4_chanx_right_out;
    wire cbx_1__8__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__8__4_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__8__4_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__8__4_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__8__5_ccff_tail;
    wire [0:29]cbx_1__8__5_chanx_left_out;
    wire [0:29]cbx_1__8__5_chanx_right_out;
    wire cbx_1__8__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__8__5_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__8__5_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__8__5_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__8__6_ccff_tail;
    wire [0:29]cbx_1__8__6_chanx_left_out;
    wire [0:29]cbx_1__8__6_chanx_right_out;
    wire cbx_1__8__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__8__6_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__8__6_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__8__6_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
    wire cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_;
    wire cbx_1__8__7_ccff_tail;
    wire [0:29]cbx_1__8__7_chanx_left_out;
    wire [0:29]cbx_1__8__7_chanx_right_out;
    wire cbx_1__8__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cbx_1__8__7_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cbx_1__8__7_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cbx_1__8__7_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_0__1__0_ccff_tail;
    wire [0:29]cby_0__1__0_chany_bottom_out;
    wire [0:29]cby_0__1__0_chany_top_out;
    wire cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_0__1__1_ccff_tail;
    wire [0:29]cby_0__1__1_chany_bottom_out;
    wire [0:29]cby_0__1__1_chany_top_out;
    wire cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_0__1__2_ccff_tail;
    wire [0:29]cby_0__1__2_chany_bottom_out;
    wire [0:29]cby_0__1__2_chany_top_out;
    wire cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_0__1__3_ccff_tail;
    wire [0:29]cby_0__1__3_chany_bottom_out;
    wire [0:29]cby_0__1__3_chany_top_out;
    wire cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_0__1__4_ccff_tail;
    wire [0:29]cby_0__1__4_chany_bottom_out;
    wire [0:29]cby_0__1__4_chany_top_out;
    wire cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_0__1__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_0__1__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_0__1__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_0__1__5_ccff_tail;
    wire [0:29]cby_0__1__5_chany_bottom_out;
    wire [0:29]cby_0__1__5_chany_top_out;
    wire cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_0__1__5_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_0__1__5_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_0__1__5_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_0__1__6_ccff_tail;
    wire [0:29]cby_0__1__6_chany_bottom_out;
    wire [0:29]cby_0__1__6_chany_top_out;
    wire cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_0__1__6_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_0__1__6_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_0__1__6_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_0__1__7_ccff_tail;
    wire [0:29]cby_0__1__7_chany_bottom_out;
    wire [0:29]cby_0__1__7_chany_top_out;
    wire cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_0__1__7_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_0__1__7_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_0__1__7_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_1__1__0_ccff_tail;
    wire [0:29]cby_1__1__0_chany_bottom_out;
    wire [0:29]cby_1__1__0_chany_top_out;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__10_ccff_tail;
    wire [0:29]cby_1__1__10_chany_bottom_out;
    wire [0:29]cby_1__1__10_chany_top_out;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__11_ccff_tail;
    wire [0:29]cby_1__1__11_chany_bottom_out;
    wire [0:29]cby_1__1__11_chany_top_out;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__12_ccff_tail;
    wire [0:29]cby_1__1__12_chany_bottom_out;
    wire [0:29]cby_1__1__12_chany_top_out;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__13_ccff_tail;
    wire [0:29]cby_1__1__13_chany_bottom_out;
    wire [0:29]cby_1__1__13_chany_top_out;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__14_ccff_tail;
    wire [0:29]cby_1__1__14_chany_bottom_out;
    wire [0:29]cby_1__1__14_chany_top_out;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__15_ccff_tail;
    wire [0:29]cby_1__1__15_chany_bottom_out;
    wire [0:29]cby_1__1__15_chany_top_out;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__16_ccff_tail;
    wire [0:29]cby_1__1__16_chany_bottom_out;
    wire [0:29]cby_1__1__16_chany_top_out;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__17_ccff_tail;
    wire [0:29]cby_1__1__17_chany_bottom_out;
    wire [0:29]cby_1__1__17_chany_top_out;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__18_ccff_tail;
    wire [0:29]cby_1__1__18_chany_bottom_out;
    wire [0:29]cby_1__1__18_chany_top_out;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__19_ccff_tail;
    wire [0:29]cby_1__1__19_chany_bottom_out;
    wire [0:29]cby_1__1__19_chany_top_out;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__1_ccff_tail;
    wire [0:29]cby_1__1__1_chany_bottom_out;
    wire [0:29]cby_1__1__1_chany_top_out;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__20_ccff_tail;
    wire [0:29]cby_1__1__20_chany_bottom_out;
    wire [0:29]cby_1__1__20_chany_top_out;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__21_ccff_tail;
    wire [0:29]cby_1__1__21_chany_bottom_out;
    wire [0:29]cby_1__1__21_chany_top_out;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__22_ccff_tail;
    wire [0:29]cby_1__1__22_chany_bottom_out;
    wire [0:29]cby_1__1__22_chany_top_out;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__23_ccff_tail;
    wire [0:29]cby_1__1__23_chany_bottom_out;
    wire [0:29]cby_1__1__23_chany_top_out;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__24_ccff_tail;
    wire [0:29]cby_1__1__24_chany_bottom_out;
    wire [0:29]cby_1__1__24_chany_top_out;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__25_ccff_tail;
    wire [0:29]cby_1__1__25_chany_bottom_out;
    wire [0:29]cby_1__1__25_chany_top_out;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__26_ccff_tail;
    wire [0:29]cby_1__1__26_chany_bottom_out;
    wire [0:29]cby_1__1__26_chany_top_out;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__27_ccff_tail;
    wire [0:29]cby_1__1__27_chany_bottom_out;
    wire [0:29]cby_1__1__27_chany_top_out;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__28_ccff_tail;
    wire [0:29]cby_1__1__28_chany_bottom_out;
    wire [0:29]cby_1__1__28_chany_top_out;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__29_ccff_tail;
    wire [0:29]cby_1__1__29_chany_bottom_out;
    wire [0:29]cby_1__1__29_chany_top_out;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__2_ccff_tail;
    wire [0:29]cby_1__1__2_chany_bottom_out;
    wire [0:29]cby_1__1__2_chany_top_out;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__30_ccff_tail;
    wire [0:29]cby_1__1__30_chany_bottom_out;
    wire [0:29]cby_1__1__30_chany_top_out;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__31_ccff_tail;
    wire [0:29]cby_1__1__31_chany_bottom_out;
    wire [0:29]cby_1__1__31_chany_top_out;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__32_ccff_tail;
    wire [0:29]cby_1__1__32_chany_bottom_out;
    wire [0:29]cby_1__1__32_chany_top_out;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__33_ccff_tail;
    wire [0:29]cby_1__1__33_chany_bottom_out;
    wire [0:29]cby_1__1__33_chany_top_out;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__34_ccff_tail;
    wire [0:29]cby_1__1__34_chany_bottom_out;
    wire [0:29]cby_1__1__34_chany_top_out;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__35_ccff_tail;
    wire [0:29]cby_1__1__35_chany_bottom_out;
    wire [0:29]cby_1__1__35_chany_top_out;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__36_ccff_tail;
    wire [0:29]cby_1__1__36_chany_bottom_out;
    wire [0:29]cby_1__1__36_chany_top_out;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__37_ccff_tail;
    wire [0:29]cby_1__1__37_chany_bottom_out;
    wire [0:29]cby_1__1__37_chany_top_out;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__38_ccff_tail;
    wire [0:29]cby_1__1__38_chany_bottom_out;
    wire [0:29]cby_1__1__38_chany_top_out;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__39_ccff_tail;
    wire [0:29]cby_1__1__39_chany_bottom_out;
    wire [0:29]cby_1__1__39_chany_top_out;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__3_ccff_tail;
    wire [0:29]cby_1__1__3_chany_bottom_out;
    wire [0:29]cby_1__1__3_chany_top_out;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__40_ccff_tail;
    wire [0:29]cby_1__1__40_chany_bottom_out;
    wire [0:29]cby_1__1__40_chany_top_out;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__41_ccff_tail;
    wire [0:29]cby_1__1__41_chany_bottom_out;
    wire [0:29]cby_1__1__41_chany_top_out;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__42_ccff_tail;
    wire [0:29]cby_1__1__42_chany_bottom_out;
    wire [0:29]cby_1__1__42_chany_top_out;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__43_ccff_tail;
    wire [0:29]cby_1__1__43_chany_bottom_out;
    wire [0:29]cby_1__1__43_chany_top_out;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__44_ccff_tail;
    wire [0:29]cby_1__1__44_chany_bottom_out;
    wire [0:29]cby_1__1__44_chany_top_out;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__45_ccff_tail;
    wire [0:29]cby_1__1__45_chany_bottom_out;
    wire [0:29]cby_1__1__45_chany_top_out;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__46_ccff_tail;
    wire [0:29]cby_1__1__46_chany_bottom_out;
    wire [0:29]cby_1__1__46_chany_top_out;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__47_ccff_tail;
    wire [0:29]cby_1__1__47_chany_bottom_out;
    wire [0:29]cby_1__1__47_chany_top_out;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__48_ccff_tail;
    wire [0:29]cby_1__1__48_chany_bottom_out;
    wire [0:29]cby_1__1__48_chany_top_out;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__49_ccff_tail;
    wire [0:29]cby_1__1__49_chany_bottom_out;
    wire [0:29]cby_1__1__49_chany_top_out;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__4_ccff_tail;
    wire [0:29]cby_1__1__4_chany_bottom_out;
    wire [0:29]cby_1__1__4_chany_top_out;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__50_ccff_tail;
    wire [0:29]cby_1__1__50_chany_bottom_out;
    wire [0:29]cby_1__1__50_chany_top_out;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__51_ccff_tail;
    wire [0:29]cby_1__1__51_chany_bottom_out;
    wire [0:29]cby_1__1__51_chany_top_out;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__52_ccff_tail;
    wire [0:29]cby_1__1__52_chany_bottom_out;
    wire [0:29]cby_1__1__52_chany_top_out;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__53_ccff_tail;
    wire [0:29]cby_1__1__53_chany_bottom_out;
    wire [0:29]cby_1__1__53_chany_top_out;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__54_ccff_tail;
    wire [0:29]cby_1__1__54_chany_bottom_out;
    wire [0:29]cby_1__1__54_chany_top_out;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__55_ccff_tail;
    wire [0:29]cby_1__1__55_chany_bottom_out;
    wire [0:29]cby_1__1__55_chany_top_out;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__5_ccff_tail;
    wire [0:29]cby_1__1__5_chany_bottom_out;
    wire [0:29]cby_1__1__5_chany_top_out;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__6_ccff_tail;
    wire [0:29]cby_1__1__6_chany_bottom_out;
    wire [0:29]cby_1__1__6_chany_top_out;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__7_ccff_tail;
    wire [0:29]cby_1__1__7_chany_bottom_out;
    wire [0:29]cby_1__1__7_chany_top_out;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__8_ccff_tail;
    wire [0:29]cby_1__1__8_chany_bottom_out;
    wire [0:29]cby_1__1__8_chany_top_out;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_1__1__9_ccff_tail;
    wire [0:29]cby_1__1__9_chany_bottom_out;
    wire [0:29]cby_1__1__9_chany_top_out;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_8__1__0_ccff_tail;
    wire [0:29]cby_8__1__0_chany_bottom_out;
    wire [0:29]cby_8__1__0_chany_top_out;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_8__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_8__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_8__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_8__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_8__1__1_ccff_tail;
    wire [0:29]cby_8__1__1_chany_bottom_out;
    wire [0:29]cby_8__1__1_chany_top_out;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_8__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_8__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_8__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_8__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_8__1__2_ccff_tail;
    wire [0:29]cby_8__1__2_chany_bottom_out;
    wire [0:29]cby_8__1__2_chany_top_out;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_8__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_8__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_8__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_8__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_8__1__3_ccff_tail;
    wire [0:29]cby_8__1__3_chany_bottom_out;
    wire [0:29]cby_8__1__3_chany_top_out;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_8__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_8__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_8__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_8__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_8__1__4_ccff_tail;
    wire [0:29]cby_8__1__4_chany_bottom_out;
    wire [0:29]cby_8__1__4_chany_top_out;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_8__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_8__1__4_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_8__1__4_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_8__1__4_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_8__1__5_ccff_tail;
    wire [0:29]cby_8__1__5_chany_bottom_out;
    wire [0:29]cby_8__1__5_chany_top_out;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_8__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_8__1__5_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_8__1__5_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_8__1__5_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_8__1__6_ccff_tail;
    wire [0:29]cby_8__1__6_chany_bottom_out;
    wire [0:29]cby_8__1__6_chany_top_out;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_8__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_8__1__6_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_8__1__6_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_8__1__6_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
    wire cby_8__1__7_ccff_tail;
    wire [0:29]cby_8__1__7_chany_bottom_out;
    wire [0:29]cby_8__1__7_chany_top_out;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
    wire cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_;
    wire cby_8__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
    wire cby_8__1__7_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
    wire cby_8__1__7_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
    wire cby_8__1__7_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
    wire ccff_head;
    wire ccff_tail;
    wire clk;
    wire direct_interc_0_out;
    wire direct_interc_100_out;
    wire direct_interc_101_out;
    wire direct_interc_102_out;
    wire direct_interc_103_out;
    wire direct_interc_104_out;
    wire direct_interc_105_out;
    wire direct_interc_106_out;
    wire direct_interc_107_out;
    wire direct_interc_108_out;
    wire direct_interc_109_out;
    wire direct_interc_10_out;
    wire direct_interc_110_out;
    wire direct_interc_111_out;
    wire direct_interc_112_out;
    wire direct_interc_113_out;
    wire direct_interc_114_out;
    wire direct_interc_115_out;
    wire direct_interc_116_out;
    wire direct_interc_117_out;
    wire direct_interc_118_out;
    wire direct_interc_119_out;
    wire direct_interc_11_out;
    wire direct_interc_120_out;
    wire direct_interc_121_out;
    wire direct_interc_122_out;
    wire direct_interc_123_out;
    wire direct_interc_124_out;
    wire direct_interc_125_out;
    wire direct_interc_126_out;
    wire direct_interc_127_out;
    wire direct_interc_128_out;
    wire direct_interc_129_out;
    wire direct_interc_12_out;
    wire direct_interc_130_out;
    wire direct_interc_131_out;
    wire direct_interc_132_out;
    wire direct_interc_133_out;
    wire direct_interc_134_out;
    wire direct_interc_135_out;
    wire direct_interc_136_out;
    wire direct_interc_137_out;
    wire direct_interc_138_out;
    wire direct_interc_139_out;
    wire direct_interc_13_out;
    wire direct_interc_140_out;
    wire direct_interc_141_out;
    wire direct_interc_142_out;
    wire direct_interc_143_out;
    wire direct_interc_144_out;
    wire direct_interc_145_out;
    wire direct_interc_146_out;
    wire direct_interc_147_out;
    wire direct_interc_148_out;
    wire direct_interc_149_out;
    wire direct_interc_14_out;
    wire direct_interc_150_out;
    wire direct_interc_151_out;
    wire direct_interc_152_out;
    wire direct_interc_153_out;
    wire direct_interc_154_out;
    wire direct_interc_155_out;
    wire direct_interc_156_out;
    wire direct_interc_157_out;
    wire direct_interc_158_out;
    wire direct_interc_159_out;
    wire direct_interc_15_out;
    wire direct_interc_160_out;
    wire direct_interc_161_out;
    wire direct_interc_162_out;
    wire direct_interc_163_out;
    wire direct_interc_164_out;
    wire direct_interc_165_out;
    wire direct_interc_166_out;
    wire direct_interc_167_out;
    wire direct_interc_168_out;
    wire direct_interc_169_out;
    wire direct_interc_16_out;
    wire direct_interc_170_out;
    wire direct_interc_171_out;
    wire direct_interc_172_out;
    wire direct_interc_173_out;
    wire direct_interc_174_out;
    wire direct_interc_17_out;
    wire direct_interc_18_out;
    wire direct_interc_19_out;
    wire direct_interc_1_out;
    wire direct_interc_20_out;
    wire direct_interc_21_out;
    wire direct_interc_22_out;
    wire direct_interc_23_out;
    wire direct_interc_24_out;
    wire direct_interc_25_out;
    wire direct_interc_26_out;
    wire direct_interc_27_out;
    wire direct_interc_28_out;
    wire direct_interc_29_out;
    wire direct_interc_2_out;
    wire direct_interc_30_out;
    wire direct_interc_31_out;
    wire direct_interc_32_out;
    wire direct_interc_33_out;
    wire direct_interc_34_out;
    wire direct_interc_35_out;
    wire direct_interc_36_out;
    wire direct_interc_37_out;
    wire direct_interc_38_out;
    wire direct_interc_39_out;
    wire direct_interc_3_out;
    wire direct_interc_40_out;
    wire direct_interc_41_out;
    wire direct_interc_42_out;
    wire direct_interc_43_out;
    wire direct_interc_44_out;
    wire direct_interc_45_out;
    wire direct_interc_46_out;
    wire direct_interc_47_out;
    wire direct_interc_48_out;
    wire direct_interc_49_out;
    wire direct_interc_4_out;
    wire direct_interc_50_out;
    wire direct_interc_51_out;
    wire direct_interc_52_out;
    wire direct_interc_53_out;
    wire direct_interc_54_out;
    wire direct_interc_55_out;
    wire direct_interc_56_out;
    wire direct_interc_57_out;
    wire direct_interc_58_out;
    wire direct_interc_59_out;
    wire direct_interc_5_out;
    wire direct_interc_60_out;
    wire direct_interc_61_out;
    wire direct_interc_62_out;
    wire direct_interc_63_out;
    wire direct_interc_64_out;
    wire direct_interc_65_out;
    wire direct_interc_66_out;
    wire direct_interc_67_out;
    wire direct_interc_68_out;
    wire direct_interc_69_out;
    wire direct_interc_6_out;
    wire direct_interc_70_out;
    wire direct_interc_71_out;
    wire direct_interc_72_out;
    wire direct_interc_73_out;
    wire direct_interc_74_out;
    wire direct_interc_75_out;
    wire direct_interc_76_out;
    wire direct_interc_77_out;
    wire direct_interc_78_out;
    wire direct_interc_79_out;
    wire direct_interc_7_out;
    wire direct_interc_80_out;
    wire direct_interc_81_out;
    wire direct_interc_82_out;
    wire direct_interc_83_out;
    wire direct_interc_84_out;
    wire direct_interc_85_out;
    wire direct_interc_86_out;
    wire direct_interc_87_out;
    wire direct_interc_88_out;
    wire direct_interc_89_out;
    wire direct_interc_8_out;
    wire direct_interc_90_out;
    wire direct_interc_91_out;
    wire direct_interc_92_out;
    wire direct_interc_93_out;
    wire direct_interc_94_out;
    wire direct_interc_95_out;
    wire direct_interc_96_out;
    wire direct_interc_97_out;
    wire direct_interc_98_out;
    wire direct_interc_99_out;
    wire direct_interc_9_out;
    wire [0:127]gfpga_pad_io_soc_dir;
    wire [0:127]gfpga_pad_io_soc_in;
    wire [0:127]gfpga_pad_io_soc_out;
    wire grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_0_ccff_tail;
    wire grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_10_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_10_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_10_ccff_tail;
    wire grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_10_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_10_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_10_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_10_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_10_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_11_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_11_ccff_tail;
    wire grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_11_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_11_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_11_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_11_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_11_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_12_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_12_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_12_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_12_ccff_tail;
    wire grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_12_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_12_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_12_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_12_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_12_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_13_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_13_ccff_tail;
    wire grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_13_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_13_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_13_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_13_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_13_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_14_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_14_ccff_tail;
    wire grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_14_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_14_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_14_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_14_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_14_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_15_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_15_ccff_tail;
    wire grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_15_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_15_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_15_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_15_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_15_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_16_ccff_tail;
    wire grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_16_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_16_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_16_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_16_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_16_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_17_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_17_ccff_tail;
    wire grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_17_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_17_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_17_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_17_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_17_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_18_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_18_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_18_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_18_ccff_tail;
    wire grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_18_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_18_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_18_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_18_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_18_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_19_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_19_ccff_tail;
    wire grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_19_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_19_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_19_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_19_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_19_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_1__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
    wire grid_clb_1__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
    wire grid_clb_1__8__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
    wire grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_1_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_1_ccff_tail;
    wire grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_20_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_20_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_20_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_20_ccff_tail;
    wire grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_20_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_20_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_20_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_20_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_20_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_21_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_21_ccff_tail;
    wire grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_21_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_21_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_21_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_21_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_21_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_22_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_22_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_22_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_22_ccff_tail;
    wire grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_22_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_22_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_22_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_22_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_22_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_22_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_23_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_23_ccff_tail;
    wire grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_23_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_23_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_23_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_23_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_23_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_23_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_24_ccff_tail;
    wire grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_24_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_24_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_24_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_24_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_24_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_24_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_25_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_25_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_25_ccff_tail;
    wire grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_25_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_25_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_25_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_25_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_25_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_25_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_26_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_26_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_26_ccff_tail;
    wire grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_26_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_26_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_26_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_26_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_26_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_26_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_27_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_27_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_27_ccff_tail;
    wire grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_27_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_27_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_27_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_27_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_27_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_27_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_28_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_28_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_28_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_28_ccff_tail;
    wire grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_28_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_28_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_28_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_28_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_28_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_28_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_29_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_29_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_29_ccff_tail;
    wire grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_29_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_29_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_29_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_29_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_29_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_29_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_2__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
    wire grid_clb_2__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
    wire grid_clb_2_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_2_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_2_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_2_ccff_tail;
    wire grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_30_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_30_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_30_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_30_ccff_tail;
    wire grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_30_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_30_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_30_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_30_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_30_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_30_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_31_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_31_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_31_ccff_tail;
    wire grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_31_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_31_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_31_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_31_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_31_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_31_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_32_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_32_ccff_tail;
    wire grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_32_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_32_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_32_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_32_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_32_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_32_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_33_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_33_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_33_ccff_tail;
    wire grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_33_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_33_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_33_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_33_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_33_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_33_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_34_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_34_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_34_ccff_tail;
    wire grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_34_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_34_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_34_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_34_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_34_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_34_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_35_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_35_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_35_ccff_tail;
    wire grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_35_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_35_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_35_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_35_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_35_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_35_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_36_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_36_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_36_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_36_ccff_tail;
    wire grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_36_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_36_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_36_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_36_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_36_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_36_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_37_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_37_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_37_ccff_tail;
    wire grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_37_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_37_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_37_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_37_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_37_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_37_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_38_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_38_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_38_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_38_ccff_tail;
    wire grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_38_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_38_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_38_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_38_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_38_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_38_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_39_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_39_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_39_ccff_tail;
    wire grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_39_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_39_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_39_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_39_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_39_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_39_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_3__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
    wire grid_clb_3__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
    wire grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_3_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_3_ccff_tail;
    wire grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_40_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_40_ccff_tail;
    wire grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_40_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_40_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_40_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_40_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_40_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_40_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_41_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_41_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_41_ccff_tail;
    wire grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_41_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_41_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_41_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_41_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_41_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_41_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_42_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_42_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_42_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_42_ccff_tail;
    wire grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_42_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_42_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_42_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_42_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_42_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_42_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_43_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_43_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_43_ccff_tail;
    wire grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_43_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_43_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_43_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_43_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_43_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_43_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_44_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_44_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_44_ccff_tail;
    wire grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_44_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_44_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_44_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_44_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_44_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_44_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_45_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_45_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_45_ccff_tail;
    wire grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_45_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_45_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_45_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_45_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_45_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_45_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_46_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_46_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_46_ccff_tail;
    wire grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_46_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_46_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_46_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_46_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_46_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_46_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_47_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_47_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_47_ccff_tail;
    wire grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_47_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_47_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_47_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_47_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_47_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_47_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_48_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_48_ccff_tail;
    wire grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_48_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_48_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_48_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_48_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_48_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_48_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_49_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_49_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_49_ccff_tail;
    wire grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_49_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_49_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_49_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_49_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_49_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_49_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_4__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
    wire grid_clb_4__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
    wire grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_4_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_4_ccff_tail;
    wire grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_4_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_4_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_4_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_4_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_4_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_50_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_50_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_50_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_50_ccff_tail;
    wire grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_50_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_50_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_50_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_50_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_50_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_50_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_51_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_51_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_51_ccff_tail;
    wire grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_51_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_51_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_51_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_51_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_51_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_51_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_52_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_52_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_52_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_52_ccff_tail;
    wire grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_52_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_52_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_52_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_52_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_52_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_52_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_53_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_53_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_53_ccff_tail;
    wire grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_53_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_53_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_53_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_53_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_53_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_53_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_54_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_54_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_54_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_54_ccff_tail;
    wire grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_54_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_54_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_54_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_54_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_54_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_54_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_55_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_55_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_55_ccff_tail;
    wire grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_55_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_55_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_55_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_55_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_55_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_55_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_56_ccff_tail;
    wire grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_56_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_56_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_56_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_56_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_56_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_56_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_57_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_57_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_57_ccff_tail;
    wire grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_57_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_57_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_57_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_57_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_57_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_57_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_58_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_58_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_58_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_58_ccff_tail;
    wire grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_58_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_58_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_58_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_58_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_58_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_58_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_59_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_59_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_59_ccff_tail;
    wire grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_59_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_59_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_59_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_59_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_59_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_59_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_5__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
    wire grid_clb_5__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
    wire grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_5_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_5_ccff_tail;
    wire grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_5_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_5_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_5_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_5_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_5_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_60_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_60_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_60_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_60_ccff_tail;
    wire grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_60_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_60_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_60_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_60_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_60_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_60_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_61_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_61_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_61_ccff_tail;
    wire grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_61_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_61_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_61_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_61_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_61_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_61_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_62_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_62_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_62_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_62_ccff_tail;
    wire grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_62_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_62_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_62_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_62_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_62_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_62_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_63_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_63_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_63_ccff_tail;
    wire grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_63_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_63_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_63_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_63_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_63_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_63_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_6__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_6__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_6__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
    wire grid_clb_6__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
    wire grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_6_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_6_ccff_tail;
    wire grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_6_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_6_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_6_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_6_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_6_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_7__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
    wire grid_clb_7__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
    wire grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_7_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_7_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_7_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_7_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_7_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_7_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_8__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
    wire grid_clb_8__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
    wire grid_clb_8_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_8_ccff_tail;
    wire grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_8_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_8_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_8_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_8_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_8_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_;
    wire grid_clb_9_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
    wire grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
    wire grid_clb_9_ccff_tail;
    wire grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_;
    wire grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_;
    wire grid_clb_9_right_width_0_height_0_subtile_0__pin_O_12_;
    wire grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_;
    wire grid_clb_9_right_width_0_height_0_subtile_0__pin_O_14_;
    wire grid_clb_9_right_width_0_height_0_subtile_0__pin_O_15_;
    wire grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_;
    wire grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_;
    wire grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_;
    wire grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_;
    wire grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_;
    wire grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_;
    wire grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_;
    wire grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_;
    wire grid_clb_9_top_width_0_height_0_subtile_0__pin_O_6_;
    wire grid_clb_9_top_width_0_height_0_subtile_0__pin_O_7_;
    wire grid_io_bottom_bottom_0_ccff_tail;
    wire grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_bottom_bottom_1_ccff_tail;
    wire grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_bottom_bottom_2_ccff_tail;
    wire grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_bottom_bottom_3_ccff_tail;
    wire grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_bottom_bottom_4_ccff_tail;
    wire grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_bottom_bottom_5_ccff_tail;
    wire grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_bottom_bottom_6_ccff_tail;
    wire grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_bottom_bottom_7_ccff_tail;
    wire grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_left_left_0_ccff_tail;
    wire grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_left_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_left_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_left_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_left_left_1_ccff_tail;
    wire grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_left_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_left_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_left_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_left_left_2_ccff_tail;
    wire grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_left_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_left_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_left_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_left_left_3_ccff_tail;
    wire grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_left_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_left_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_left_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_left_left_4_ccff_tail;
    wire grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_left_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_left_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_left_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_left_left_5_ccff_tail;
    wire grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_left_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_left_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_left_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_left_left_6_ccff_tail;
    wire grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_left_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_left_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_left_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_left_left_7_ccff_tail;
    wire grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_left_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_left_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_left_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_right_right_0_ccff_tail;
    wire grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_right_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_right_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_right_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_right_right_1_ccff_tail;
    wire grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_right_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_right_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_right_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_right_right_2_ccff_tail;
    wire grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_right_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_right_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_right_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_right_right_3_ccff_tail;
    wire grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_right_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_right_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_right_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_right_right_4_ccff_tail;
    wire grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_right_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_right_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_right_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_right_right_5_ccff_tail;
    wire grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_right_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_right_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_right_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_right_right_6_ccff_tail;
    wire grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_right_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_right_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_right_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_right_right_7_ccff_tail;
    wire grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_right_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_right_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_right_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_top_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_top_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_top_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_top_top_0_ccff_tail;
    wire grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_top_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_top_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_top_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_top_top_1_ccff_tail;
    wire grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_top_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_top_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_top_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_top_top_2_ccff_tail;
    wire grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_top_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_top_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_top_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_top_top_3_ccff_tail;
    wire grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_top_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_top_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_top_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_top_top_4_ccff_tail;
    wire grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_top_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_top_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_top_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_top_top_5_ccff_tail;
    wire grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_top_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_top_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_top_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_top_top_6_ccff_tail;
    wire grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
    wire grid_io_top_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
    wire grid_io_top_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
    wire grid_io_top_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
    wire grid_io_top_top_7_ccff_tail;
    wire isol_n;
    wire prog_clk;
    wire prog_reset;
    wire [63:0]prog_reset_ft;
    wire reset;
    wire [63:0]reset_ft;
    wire sb_0__0__0_ccff_tail;
    wire [0:29]sb_0__0__0_chanx_right_out;
    wire [0:29]sb_0__0__0_chany_top_out;
    wire sb_0__1__0_ccff_tail;
    wire [0:29]sb_0__1__0_chanx_right_out;
    wire [0:29]sb_0__1__0_chany_bottom_out;
    wire [0:29]sb_0__1__0_chany_top_out;
    wire sb_0__1__1_ccff_tail;
    wire [0:29]sb_0__1__1_chanx_right_out;
    wire [0:29]sb_0__1__1_chany_bottom_out;
    wire [0:29]sb_0__1__1_chany_top_out;
    wire sb_0__1__2_ccff_tail;
    wire [0:29]sb_0__1__2_chanx_right_out;
    wire [0:29]sb_0__1__2_chany_bottom_out;
    wire [0:29]sb_0__1__2_chany_top_out;
    wire sb_0__1__3_ccff_tail;
    wire [0:29]sb_0__1__3_chanx_right_out;
    wire [0:29]sb_0__1__3_chany_bottom_out;
    wire [0:29]sb_0__1__3_chany_top_out;
    wire sb_0__1__4_ccff_tail;
    wire [0:29]sb_0__1__4_chanx_right_out;
    wire [0:29]sb_0__1__4_chany_bottom_out;
    wire [0:29]sb_0__1__4_chany_top_out;
    wire sb_0__1__5_ccff_tail;
    wire [0:29]sb_0__1__5_chanx_right_out;
    wire [0:29]sb_0__1__5_chany_bottom_out;
    wire [0:29]sb_0__1__5_chany_top_out;
    wire sb_0__1__6_ccff_tail;
    wire [0:29]sb_0__1__6_chanx_right_out;
    wire [0:29]sb_0__1__6_chany_bottom_out;
    wire [0:29]sb_0__1__6_chany_top_out;
    wire sb_0__8__0_ccff_tail;
    wire [0:29]sb_0__8__0_chanx_right_out;
    wire [0:29]sb_0__8__0_chany_bottom_out;
    wire sb_1__0__0_ccff_tail;
    wire [0:29]sb_1__0__0_chanx_left_out;
    wire [0:29]sb_1__0__0_chanx_right_out;
    wire [0:29]sb_1__0__0_chany_top_out;
    wire sb_1__0__1_ccff_tail;
    wire [0:29]sb_1__0__1_chanx_left_out;
    wire [0:29]sb_1__0__1_chanx_right_out;
    wire [0:29]sb_1__0__1_chany_top_out;
    wire sb_1__0__2_ccff_tail;
    wire [0:29]sb_1__0__2_chanx_left_out;
    wire [0:29]sb_1__0__2_chanx_right_out;
    wire [0:29]sb_1__0__2_chany_top_out;
    wire sb_1__0__3_ccff_tail;
    wire [0:29]sb_1__0__3_chanx_left_out;
    wire [0:29]sb_1__0__3_chanx_right_out;
    wire [0:29]sb_1__0__3_chany_top_out;
    wire sb_1__0__4_ccff_tail;
    wire [0:29]sb_1__0__4_chanx_left_out;
    wire [0:29]sb_1__0__4_chanx_right_out;
    wire [0:29]sb_1__0__4_chany_top_out;
    wire sb_1__0__5_ccff_tail;
    wire [0:29]sb_1__0__5_chanx_left_out;
    wire [0:29]sb_1__0__5_chanx_right_out;
    wire [0:29]sb_1__0__5_chany_top_out;
    wire sb_1__0__6_ccff_tail;
    wire [0:29]sb_1__0__6_chanx_left_out;
    wire [0:29]sb_1__0__6_chanx_right_out;
    wire [0:29]sb_1__0__6_chany_top_out;
    wire sb_1__1__0_ccff_tail;
    wire [0:29]sb_1__1__0_chanx_left_out;
    wire [0:29]sb_1__1__0_chanx_right_out;
    wire [0:29]sb_1__1__0_chany_bottom_out;
    wire [0:29]sb_1__1__0_chany_top_out;
    wire sb_1__1__10_ccff_tail;
    wire [0:29]sb_1__1__10_chanx_left_out;
    wire [0:29]sb_1__1__10_chanx_right_out;
    wire [0:29]sb_1__1__10_chany_bottom_out;
    wire [0:29]sb_1__1__10_chany_top_out;
    wire sb_1__1__11_ccff_tail;
    wire [0:29]sb_1__1__11_chanx_left_out;
    wire [0:29]sb_1__1__11_chanx_right_out;
    wire [0:29]sb_1__1__11_chany_bottom_out;
    wire [0:29]sb_1__1__11_chany_top_out;
    wire sb_1__1__12_ccff_tail;
    wire [0:29]sb_1__1__12_chanx_left_out;
    wire [0:29]sb_1__1__12_chanx_right_out;
    wire [0:29]sb_1__1__12_chany_bottom_out;
    wire [0:29]sb_1__1__12_chany_top_out;
    wire sb_1__1__13_ccff_tail;
    wire [0:29]sb_1__1__13_chanx_left_out;
    wire [0:29]sb_1__1__13_chanx_right_out;
    wire [0:29]sb_1__1__13_chany_bottom_out;
    wire [0:29]sb_1__1__13_chany_top_out;
    wire sb_1__1__14_ccff_tail;
    wire [0:29]sb_1__1__14_chanx_left_out;
    wire [0:29]sb_1__1__14_chanx_right_out;
    wire [0:29]sb_1__1__14_chany_bottom_out;
    wire [0:29]sb_1__1__14_chany_top_out;
    wire sb_1__1__15_ccff_tail;
    wire [0:29]sb_1__1__15_chanx_left_out;
    wire [0:29]sb_1__1__15_chanx_right_out;
    wire [0:29]sb_1__1__15_chany_bottom_out;
    wire [0:29]sb_1__1__15_chany_top_out;
    wire sb_1__1__16_ccff_tail;
    wire [0:29]sb_1__1__16_chanx_left_out;
    wire [0:29]sb_1__1__16_chanx_right_out;
    wire [0:29]sb_1__1__16_chany_bottom_out;
    wire [0:29]sb_1__1__16_chany_top_out;
    wire sb_1__1__17_ccff_tail;
    wire [0:29]sb_1__1__17_chanx_left_out;
    wire [0:29]sb_1__1__17_chanx_right_out;
    wire [0:29]sb_1__1__17_chany_bottom_out;
    wire [0:29]sb_1__1__17_chany_top_out;
    wire sb_1__1__18_ccff_tail;
    wire [0:29]sb_1__1__18_chanx_left_out;
    wire [0:29]sb_1__1__18_chanx_right_out;
    wire [0:29]sb_1__1__18_chany_bottom_out;
    wire [0:29]sb_1__1__18_chany_top_out;
    wire sb_1__1__19_ccff_tail;
    wire [0:29]sb_1__1__19_chanx_left_out;
    wire [0:29]sb_1__1__19_chanx_right_out;
    wire [0:29]sb_1__1__19_chany_bottom_out;
    wire [0:29]sb_1__1__19_chany_top_out;
    wire sb_1__1__1_ccff_tail;
    wire [0:29]sb_1__1__1_chanx_left_out;
    wire [0:29]sb_1__1__1_chanx_right_out;
    wire [0:29]sb_1__1__1_chany_bottom_out;
    wire [0:29]sb_1__1__1_chany_top_out;
    wire sb_1__1__20_ccff_tail;
    wire [0:29]sb_1__1__20_chanx_left_out;
    wire [0:29]sb_1__1__20_chanx_right_out;
    wire [0:29]sb_1__1__20_chany_bottom_out;
    wire [0:29]sb_1__1__20_chany_top_out;
    wire sb_1__1__21_ccff_tail;
    wire [0:29]sb_1__1__21_chanx_left_out;
    wire [0:29]sb_1__1__21_chanx_right_out;
    wire [0:29]sb_1__1__21_chany_bottom_out;
    wire [0:29]sb_1__1__21_chany_top_out;
    wire sb_1__1__22_ccff_tail;
    wire [0:29]sb_1__1__22_chanx_left_out;
    wire [0:29]sb_1__1__22_chanx_right_out;
    wire [0:29]sb_1__1__22_chany_bottom_out;
    wire [0:29]sb_1__1__22_chany_top_out;
    wire sb_1__1__23_ccff_tail;
    wire [0:29]sb_1__1__23_chanx_left_out;
    wire [0:29]sb_1__1__23_chanx_right_out;
    wire [0:29]sb_1__1__23_chany_bottom_out;
    wire [0:29]sb_1__1__23_chany_top_out;
    wire sb_1__1__24_ccff_tail;
    wire [0:29]sb_1__1__24_chanx_left_out;
    wire [0:29]sb_1__1__24_chanx_right_out;
    wire [0:29]sb_1__1__24_chany_bottom_out;
    wire [0:29]sb_1__1__24_chany_top_out;
    wire sb_1__1__25_ccff_tail;
    wire [0:29]sb_1__1__25_chanx_left_out;
    wire [0:29]sb_1__1__25_chanx_right_out;
    wire [0:29]sb_1__1__25_chany_bottom_out;
    wire [0:29]sb_1__1__25_chany_top_out;
    wire sb_1__1__26_ccff_tail;
    wire [0:29]sb_1__1__26_chanx_left_out;
    wire [0:29]sb_1__1__26_chanx_right_out;
    wire [0:29]sb_1__1__26_chany_bottom_out;
    wire [0:29]sb_1__1__26_chany_top_out;
    wire sb_1__1__27_ccff_tail;
    wire [0:29]sb_1__1__27_chanx_left_out;
    wire [0:29]sb_1__1__27_chanx_right_out;
    wire [0:29]sb_1__1__27_chany_bottom_out;
    wire [0:29]sb_1__1__27_chany_top_out;
    wire sb_1__1__28_ccff_tail;
    wire [0:29]sb_1__1__28_chanx_left_out;
    wire [0:29]sb_1__1__28_chanx_right_out;
    wire [0:29]sb_1__1__28_chany_bottom_out;
    wire [0:29]sb_1__1__28_chany_top_out;
    wire sb_1__1__29_ccff_tail;
    wire [0:29]sb_1__1__29_chanx_left_out;
    wire [0:29]sb_1__1__29_chanx_right_out;
    wire [0:29]sb_1__1__29_chany_bottom_out;
    wire [0:29]sb_1__1__29_chany_top_out;
    wire sb_1__1__2_ccff_tail;
    wire [0:29]sb_1__1__2_chanx_left_out;
    wire [0:29]sb_1__1__2_chanx_right_out;
    wire [0:29]sb_1__1__2_chany_bottom_out;
    wire [0:29]sb_1__1__2_chany_top_out;
    wire sb_1__1__30_ccff_tail;
    wire [0:29]sb_1__1__30_chanx_left_out;
    wire [0:29]sb_1__1__30_chanx_right_out;
    wire [0:29]sb_1__1__30_chany_bottom_out;
    wire [0:29]sb_1__1__30_chany_top_out;
    wire sb_1__1__31_ccff_tail;
    wire [0:29]sb_1__1__31_chanx_left_out;
    wire [0:29]sb_1__1__31_chanx_right_out;
    wire [0:29]sb_1__1__31_chany_bottom_out;
    wire [0:29]sb_1__1__31_chany_top_out;
    wire sb_1__1__32_ccff_tail;
    wire [0:29]sb_1__1__32_chanx_left_out;
    wire [0:29]sb_1__1__32_chanx_right_out;
    wire [0:29]sb_1__1__32_chany_bottom_out;
    wire [0:29]sb_1__1__32_chany_top_out;
    wire sb_1__1__33_ccff_tail;
    wire [0:29]sb_1__1__33_chanx_left_out;
    wire [0:29]sb_1__1__33_chanx_right_out;
    wire [0:29]sb_1__1__33_chany_bottom_out;
    wire [0:29]sb_1__1__33_chany_top_out;
    wire sb_1__1__34_ccff_tail;
    wire [0:29]sb_1__1__34_chanx_left_out;
    wire [0:29]sb_1__1__34_chanx_right_out;
    wire [0:29]sb_1__1__34_chany_bottom_out;
    wire [0:29]sb_1__1__34_chany_top_out;
    wire sb_1__1__35_ccff_tail;
    wire [0:29]sb_1__1__35_chanx_left_out;
    wire [0:29]sb_1__1__35_chanx_right_out;
    wire [0:29]sb_1__1__35_chany_bottom_out;
    wire [0:29]sb_1__1__35_chany_top_out;
    wire sb_1__1__36_ccff_tail;
    wire [0:29]sb_1__1__36_chanx_left_out;
    wire [0:29]sb_1__1__36_chanx_right_out;
    wire [0:29]sb_1__1__36_chany_bottom_out;
    wire [0:29]sb_1__1__36_chany_top_out;
    wire sb_1__1__37_ccff_tail;
    wire [0:29]sb_1__1__37_chanx_left_out;
    wire [0:29]sb_1__1__37_chanx_right_out;
    wire [0:29]sb_1__1__37_chany_bottom_out;
    wire [0:29]sb_1__1__37_chany_top_out;
    wire sb_1__1__38_ccff_tail;
    wire [0:29]sb_1__1__38_chanx_left_out;
    wire [0:29]sb_1__1__38_chanx_right_out;
    wire [0:29]sb_1__1__38_chany_bottom_out;
    wire [0:29]sb_1__1__38_chany_top_out;
    wire sb_1__1__39_ccff_tail;
    wire [0:29]sb_1__1__39_chanx_left_out;
    wire [0:29]sb_1__1__39_chanx_right_out;
    wire [0:29]sb_1__1__39_chany_bottom_out;
    wire [0:29]sb_1__1__39_chany_top_out;
    wire sb_1__1__3_ccff_tail;
    wire [0:29]sb_1__1__3_chanx_left_out;
    wire [0:29]sb_1__1__3_chanx_right_out;
    wire [0:29]sb_1__1__3_chany_bottom_out;
    wire [0:29]sb_1__1__3_chany_top_out;
    wire sb_1__1__40_ccff_tail;
    wire [0:29]sb_1__1__40_chanx_left_out;
    wire [0:29]sb_1__1__40_chanx_right_out;
    wire [0:29]sb_1__1__40_chany_bottom_out;
    wire [0:29]sb_1__1__40_chany_top_out;
    wire sb_1__1__41_ccff_tail;
    wire [0:29]sb_1__1__41_chanx_left_out;
    wire [0:29]sb_1__1__41_chanx_right_out;
    wire [0:29]sb_1__1__41_chany_bottom_out;
    wire [0:29]sb_1__1__41_chany_top_out;
    wire sb_1__1__42_ccff_tail;
    wire [0:29]sb_1__1__42_chanx_left_out;
    wire [0:29]sb_1__1__42_chanx_right_out;
    wire [0:29]sb_1__1__42_chany_bottom_out;
    wire [0:29]sb_1__1__42_chany_top_out;
    wire sb_1__1__43_ccff_tail;
    wire [0:29]sb_1__1__43_chanx_left_out;
    wire [0:29]sb_1__1__43_chanx_right_out;
    wire [0:29]sb_1__1__43_chany_bottom_out;
    wire [0:29]sb_1__1__43_chany_top_out;
    wire sb_1__1__44_ccff_tail;
    wire [0:29]sb_1__1__44_chanx_left_out;
    wire [0:29]sb_1__1__44_chanx_right_out;
    wire [0:29]sb_1__1__44_chany_bottom_out;
    wire [0:29]sb_1__1__44_chany_top_out;
    wire sb_1__1__45_ccff_tail;
    wire [0:29]sb_1__1__45_chanx_left_out;
    wire [0:29]sb_1__1__45_chanx_right_out;
    wire [0:29]sb_1__1__45_chany_bottom_out;
    wire [0:29]sb_1__1__45_chany_top_out;
    wire sb_1__1__46_ccff_tail;
    wire [0:29]sb_1__1__46_chanx_left_out;
    wire [0:29]sb_1__1__46_chanx_right_out;
    wire [0:29]sb_1__1__46_chany_bottom_out;
    wire [0:29]sb_1__1__46_chany_top_out;
    wire sb_1__1__47_ccff_tail;
    wire [0:29]sb_1__1__47_chanx_left_out;
    wire [0:29]sb_1__1__47_chanx_right_out;
    wire [0:29]sb_1__1__47_chany_bottom_out;
    wire [0:29]sb_1__1__47_chany_top_out;
    wire sb_1__1__48_ccff_tail;
    wire [0:29]sb_1__1__48_chanx_left_out;
    wire [0:29]sb_1__1__48_chanx_right_out;
    wire [0:29]sb_1__1__48_chany_bottom_out;
    wire [0:29]sb_1__1__48_chany_top_out;
    wire sb_1__1__4_ccff_tail;
    wire [0:29]sb_1__1__4_chanx_left_out;
    wire [0:29]sb_1__1__4_chanx_right_out;
    wire [0:29]sb_1__1__4_chany_bottom_out;
    wire [0:29]sb_1__1__4_chany_top_out;
    wire sb_1__1__5_ccff_tail;
    wire [0:29]sb_1__1__5_chanx_left_out;
    wire [0:29]sb_1__1__5_chanx_right_out;
    wire [0:29]sb_1__1__5_chany_bottom_out;
    wire [0:29]sb_1__1__5_chany_top_out;
    wire sb_1__1__6_ccff_tail;
    wire [0:29]sb_1__1__6_chanx_left_out;
    wire [0:29]sb_1__1__6_chanx_right_out;
    wire [0:29]sb_1__1__6_chany_bottom_out;
    wire [0:29]sb_1__1__6_chany_top_out;
    wire sb_1__1__7_ccff_tail;
    wire [0:29]sb_1__1__7_chanx_left_out;
    wire [0:29]sb_1__1__7_chanx_right_out;
    wire [0:29]sb_1__1__7_chany_bottom_out;
    wire [0:29]sb_1__1__7_chany_top_out;
    wire sb_1__1__8_ccff_tail;
    wire [0:29]sb_1__1__8_chanx_left_out;
    wire [0:29]sb_1__1__8_chanx_right_out;
    wire [0:29]sb_1__1__8_chany_bottom_out;
    wire [0:29]sb_1__1__8_chany_top_out;
    wire sb_1__1__9_ccff_tail;
    wire [0:29]sb_1__1__9_chanx_left_out;
    wire [0:29]sb_1__1__9_chanx_right_out;
    wire [0:29]sb_1__1__9_chany_bottom_out;
    wire [0:29]sb_1__1__9_chany_top_out;
    wire sb_1__8__0_ccff_tail;
    wire [0:29]sb_1__8__0_chanx_left_out;
    wire [0:29]sb_1__8__0_chanx_right_out;
    wire [0:29]sb_1__8__0_chany_bottom_out;
    wire sb_1__8__1_ccff_tail;
    wire [0:29]sb_1__8__1_chanx_left_out;
    wire [0:29]sb_1__8__1_chanx_right_out;
    wire [0:29]sb_1__8__1_chany_bottom_out;
    wire sb_1__8__2_ccff_tail;
    wire [0:29]sb_1__8__2_chanx_left_out;
    wire [0:29]sb_1__8__2_chanx_right_out;
    wire [0:29]sb_1__8__2_chany_bottom_out;
    wire sb_1__8__3_ccff_tail;
    wire [0:29]sb_1__8__3_chanx_left_out;
    wire [0:29]sb_1__8__3_chanx_right_out;
    wire [0:29]sb_1__8__3_chany_bottom_out;
    wire sb_1__8__4_ccff_tail;
    wire [0:29]sb_1__8__4_chanx_left_out;
    wire [0:29]sb_1__8__4_chanx_right_out;
    wire [0:29]sb_1__8__4_chany_bottom_out;
    wire sb_1__8__5_ccff_tail;
    wire [0:29]sb_1__8__5_chanx_left_out;
    wire [0:29]sb_1__8__5_chanx_right_out;
    wire [0:29]sb_1__8__5_chany_bottom_out;
    wire sb_1__8__6_ccff_tail;
    wire [0:29]sb_1__8__6_chanx_left_out;
    wire [0:29]sb_1__8__6_chanx_right_out;
    wire [0:29]sb_1__8__6_chany_bottom_out;
    wire sb_8__0__0_ccff_tail;
    wire [0:29]sb_8__0__0_chanx_left_out;
    wire [0:29]sb_8__0__0_chany_top_out;
    wire sb_8__1__0_ccff_tail;
    wire [0:29]sb_8__1__0_chanx_left_out;
    wire [0:29]sb_8__1__0_chany_bottom_out;
    wire [0:29]sb_8__1__0_chany_top_out;
    wire sb_8__1__1_ccff_tail;
    wire [0:29]sb_8__1__1_chanx_left_out;
    wire [0:29]sb_8__1__1_chany_bottom_out;
    wire [0:29]sb_8__1__1_chany_top_out;
    wire sb_8__1__2_ccff_tail;
    wire [0:29]sb_8__1__2_chanx_left_out;
    wire [0:29]sb_8__1__2_chany_bottom_out;
    wire [0:29]sb_8__1__2_chany_top_out;
    wire sb_8__1__3_ccff_tail;
    wire [0:29]sb_8__1__3_chanx_left_out;
    wire [0:29]sb_8__1__3_chany_bottom_out;
    wire [0:29]sb_8__1__3_chany_top_out;
    wire sb_8__1__4_ccff_tail;
    wire [0:29]sb_8__1__4_chanx_left_out;
    wire [0:29]sb_8__1__4_chany_bottom_out;
    wire [0:29]sb_8__1__4_chany_top_out;
    wire sb_8__1__5_ccff_tail;
    wire [0:29]sb_8__1__5_chanx_left_out;
    wire [0:29]sb_8__1__5_chany_bottom_out;
    wire [0:29]sb_8__1__5_chany_top_out;
    wire sb_8__1__6_ccff_tail;
    wire [0:29]sb_8__1__6_chanx_left_out;
    wire [0:29]sb_8__1__6_chany_bottom_out;
    wire [0:29]sb_8__1__6_chany_top_out;
    wire sb_8__8__0_ccff_tail;
    wire [0:29]sb_8__8__0_chanx_left_out;
    wire [0:29]sb_8__8__0_chany_bottom_out;
    wire scan_enable;

assign prog_reset_ft[0] = prog_reset;
assign reset_ft[0] = reset;
    bottom_left_tile tile_1__1_
    (
        .ccff_head(grid_io_left_left_1_ccff_tail),
        .chanx_right_in(cbx_1__0__0_chanx_left_out),
        .chany_top_in(cby_0__1__0_chany_bottom_out),
        .prog_clk(prog_clk),
        .prog_reset_top_in(prog_reset_ft[4]),
        .reset_top_in(reset_ft[63]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(sb_0__0__0_ccff_tail),
        .chanx_right_out(sb_0__0__0_chanx_right_out),
        .chany_top_out(sb_0__0__0_chany_top_out)
    );
    left_tile tile_1__2_
    (
        .ccff_head(grid_io_left_left_2_ccff_tail),
        .ccff_head_0(sb_0__0__0_ccff_tail),
        .chanx_right_in(cbx_1__1__0_chanx_left_out),
        .chany_bottom_in(sb_0__0__0_chany_top_out),
        .chany_top_in_0(cby_0__1__1_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[96:99]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[3]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[62]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_io_left_left_0_ccff_tail),
        .ccff_tail_0(sb_0__1__0_ccff_tail),
        .chanx_right_out(sb_0__1__0_chanx_right_out),
        .chany_bottom_out(cby_0__1__0_chany_bottom_out),
        .chany_top_out_0(sb_0__1__0_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[96:99]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[96:99]),
        .prog_reset_bottom_out(prog_reset_ft[4]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[63]),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    left_tile tile_1__3_
    (
        .ccff_head(grid_io_left_left_3_ccff_tail),
        .ccff_head_0(sb_0__1__0_ccff_tail),
        .chanx_right_in(cbx_1__1__1_chanx_left_out),
        .chany_bottom_in(sb_0__1__0_chany_top_out),
        .chany_top_in_0(cby_0__1__2_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[100:103]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[2]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[61]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_io_left_left_1_ccff_tail),
        .ccff_tail_0(sb_0__1__1_ccff_tail),
        .chanx_right_out(sb_0__1__1_chanx_right_out),
        .chany_bottom_out(cby_0__1__1_chany_bottom_out),
        .chany_top_out_0(sb_0__1__1_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[100:103]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[100:103]),
        .prog_reset_bottom_out(prog_reset_ft[3]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[62]),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    left_tile tile_1__4_
    (
        .ccff_head(grid_io_left_left_4_ccff_tail),
        .ccff_head_0(sb_0__1__1_ccff_tail),
        .chanx_right_in(cbx_1__1__2_chanx_left_out),
        .chany_bottom_in(sb_0__1__1_chany_top_out),
        .chany_top_in_0(cby_0__1__3_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[104:107]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[1]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[60]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_io_left_left_2_ccff_tail),
        .ccff_tail_0(sb_0__1__2_ccff_tail),
        .chanx_right_out(sb_0__1__2_chanx_right_out),
        .chany_bottom_out(cby_0__1__2_chany_bottom_out),
        .chany_top_out_0(sb_0__1__2_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[104:107]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[104:107]),
        .prog_reset_bottom_out(prog_reset_ft[2]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[61]),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    left_tile tile_1__5_
    (
        .ccff_head(grid_io_left_left_5_ccff_tail),
        .ccff_head_0(sb_0__1__2_ccff_tail),
        .chanx_right_in(cbx_1__1__3_chanx_left_out),
        .chany_bottom_in(sb_0__1__2_chany_top_out),
        .chany_top_in_0(cby_0__1__4_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[108:111]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(prog_reset_ft[0]),
        .prog_reset_top_in(),
        .reset_bottom_in(),
        .reset_right_in(reset_ft[56]),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_io_left_left_3_ccff_tail),
        .ccff_tail_0(sb_0__1__3_ccff_tail),
        .chanx_right_out(sb_0__1__3_chanx_right_out),
        .chany_bottom_out(cby_0__1__3_chany_bottom_out),
        .chany_top_out_0(sb_0__1__3_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[108:111]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[108:111]),
        .prog_reset_bottom_out(prog_reset_ft[1]),
        .prog_reset_right_out(prog_reset_ft[8]),
        .prog_reset_top_out(prog_reset_ft[5]),
        .reset_bottom_out(reset_ft[60]),
        .reset_top_out(reset_ft[57]),
        .right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    left_tile tile_1__6_
    (
        .ccff_head(grid_io_left_left_6_ccff_tail),
        .ccff_head_0(sb_0__1__3_ccff_tail),
        .chanx_right_in(cbx_1__1__4_chanx_left_out),
        .chany_bottom_in(sb_0__1__3_chany_top_out),
        .chany_top_in_0(cby_0__1__5_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[112:115]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[5]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[57]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_7_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_io_left_left_4_ccff_tail),
        .ccff_tail_0(sb_0__1__4_ccff_tail),
        .chanx_right_out(sb_0__1__4_chanx_right_out),
        .chany_bottom_out(cby_0__1__4_chany_bottom_out),
        .chany_top_out_0(sb_0__1__4_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[112:115]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[112:115]),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[6]),
        .reset_bottom_out(),
        .reset_top_out(reset_ft[58]),
        .right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    left_tile tile_1__7_
    (
        .ccff_head(grid_io_left_left_7_ccff_tail),
        .ccff_head_0(sb_0__1__4_ccff_tail),
        .chanx_right_in(cbx_1__1__5_chanx_left_out),
        .chany_bottom_in(sb_0__1__4_chany_top_out),
        .chany_top_in_0(cby_0__1__6_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[116:119]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[6]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[58]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_7_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_io_left_left_5_ccff_tail),
        .ccff_tail_0(sb_0__1__5_ccff_tail),
        .chanx_right_out(sb_0__1__5_chanx_right_out),
        .chany_bottom_out(cby_0__1__5_chany_bottom_out),
        .chany_top_out_0(sb_0__1__5_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[116:119]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[116:119]),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[7]),
        .reset_bottom_out(),
        .reset_top_out(reset_ft[59]),
        .right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    left_tile tile_1__8_
    (
        .ccff_head(sb_0__8__0_ccff_tail),
        .ccff_head_0(sb_0__1__5_ccff_tail),
        .chanx_right_in(cbx_1__1__6_chanx_left_out),
        .chany_bottom_in(sb_0__1__5_chany_top_out),
        .chany_top_in_0(cby_0__1__7_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[120:123]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[7]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[59]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_7_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_io_left_left_6_ccff_tail),
        .ccff_tail_0(sb_0__1__6_ccff_tail),
        .chanx_right_out(sb_0__1__6_chanx_right_out),
        .chany_bottom_out(cby_0__1__6_chany_bottom_out),
        .chany_top_out_0(sb_0__1__6_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[120:123]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[120:123]),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    top_left_tile tile_1__9_
    (
        .ccff_head(grid_io_top_top_0_ccff_tail),
        .ccff_head_0(sb_0__1__6_ccff_tail),
        .chanx_right_in(cbx_1__8__0_chanx_left_out),
        .chany_bottom_in_0(sb_0__1__6_chany_top_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[124:127]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_7_),
        .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(sb_0__8__0_ccff_tail),
        .ccff_tail_0(grid_io_left_left_7_ccff_tail),
        .chanx_right_out(sb_0__8__0_chanx_right_out),
        .chany_bottom_out_0(cby_0__1__7_chany_bottom_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[124:127]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[124:127]),
        .right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    bottom_tile tile_2__1_
    (
        .ccff_head(ccff_head),
        .ccff_head_1(grid_io_left_left_0_ccff_tail),
        .chanx_left_in(sb_0__0__0_chanx_right_out),
        .chanx_right_in_0(cbx_1__0__1_chanx_left_out),
        .chany_top_in(cby_1__1__0_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[92:95]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_top_in(prog_reset_ft[12]),
        .reset_top_in(reset_ft[55]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
        .ccff_tail(grid_io_bottom_bottom_7_ccff_tail),
        .ccff_tail_0(cbx_1__0__0_ccff_tail),
        .chanx_left_out(cbx_1__0__0_chanx_left_out),
        .chanx_right_out_0(sb_1__0__0_chanx_right_out),
        .chany_top_out(sb_1__0__0_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[92:95]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[92:95]),
        .top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    tile tile_2__2_
    (
        .ccff_head_1(cbx_1__0__0_ccff_tail),
        .ccff_head_2(grid_clb_9_ccff_tail),
        .chanx_left_in(sb_0__1__0_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__7_chanx_left_out),
        .chany_bottom_in(sb_1__0__0_chany_top_out),
        .chany_top_in_0(cby_1__1__1_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[11]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[54]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_0_ccff_tail),
        .ccff_tail_0(cbx_1__1__0_ccff_tail),
        .chanx_left_out(cbx_1__1__0_chanx_left_out),
        .chanx_right_out_0(sb_1__1__0_chanx_right_out),
        .chany_bottom_out(cby_1__1__0_chany_bottom_out),
        .chany_top_out_0(sb_1__1__0_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[12]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[55]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_2__3_
    (
        .ccff_head_1(cbx_1__1__0_ccff_tail),
        .ccff_head_2(grid_clb_1_ccff_tail),
        .chanx_left_in(sb_0__1__1_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__8_chanx_left_out),
        .chany_bottom_in(sb_1__1__0_chany_top_out),
        .chany_top_in_0(cby_1__1__2_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[10]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[53]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_1_ccff_tail),
        .ccff_tail_0(cbx_1__1__1_ccff_tail),
        .chanx_left_out(cbx_1__1__1_chanx_left_out),
        .chanx_right_out_0(sb_1__1__1_chanx_right_out),
        .chany_bottom_out(cby_1__1__1_chany_bottom_out),
        .chany_top_out_0(sb_1__1__1_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[11]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[54]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_2__4_
    (
        .ccff_head_1(cbx_1__1__1_ccff_tail),
        .ccff_head_2(grid_clb_11_ccff_tail),
        .chanx_left_in(sb_0__1__2_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__9_chanx_left_out),
        .chany_bottom_in(sb_1__1__1_chany_top_out),
        .chany_top_in_0(cby_1__1__3_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[9]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[52]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_2_ccff_tail),
        .ccff_tail_0(cbx_1__1__2_ccff_tail),
        .chanx_left_out(cbx_1__1__2_chanx_left_out),
        .chanx_right_out_0(sb_1__1__2_chanx_right_out),
        .chany_bottom_out(cby_1__1__2_chany_bottom_out),
        .chany_top_out_0(sb_1__1__2_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[10]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[53]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_2__5_
    (
        .ccff_head_1(cbx_1__1__2_ccff_tail),
        .ccff_head_2(grid_clb_3_ccff_tail),
        .chanx_left_in(sb_0__1__3_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__10_chanx_left_out),
        .chany_bottom_in(sb_1__1__2_chany_top_out),
        .chany_top_in_0(cby_1__1__4_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(prog_reset_ft[8]),
        .prog_reset_top_in(),
        .reset_bottom_in(),
        .reset_right_in(reset_ft[48]),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_3_ccff_tail),
        .ccff_tail_0(cbx_1__1__3_ccff_tail),
        .chanx_left_out(cbx_1__1__3_chanx_left_out),
        .chanx_right_out_0(sb_1__1__3_chanx_right_out),
        .chany_bottom_out(cby_1__1__3_chany_bottom_out),
        .chany_top_out_0(sb_1__1__3_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[9]),
        .prog_reset_right_out(prog_reset_ft[16]),
        .prog_reset_top_out(prog_reset_ft[13]),
        .reset_bottom_out(reset_ft[52]),
        .reset_left_out(reset_ft[56]),
        .reset_top_out(reset_ft[49]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_2__6_
    (
        .ccff_head_1(cbx_1__1__3_ccff_tail),
        .ccff_head_2(grid_clb_13_ccff_tail),
        .chanx_left_in(sb_0__1__4_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__11_chanx_left_out),
        .chany_bottom_in(sb_1__1__3_chany_top_out),
        .chany_top_in_0(cby_1__1__5_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[13]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[49]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_4_ccff_tail),
        .ccff_tail_0(cbx_1__1__4_ccff_tail),
        .chanx_left_out(cbx_1__1__4_chanx_left_out),
        .chanx_right_out_0(sb_1__1__4_chanx_right_out),
        .chany_bottom_out(cby_1__1__4_chany_bottom_out),
        .chany_top_out_0(sb_1__1__4_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[14]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[50]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_2__7_
    (
        .ccff_head_1(cbx_1__1__4_ccff_tail),
        .ccff_head_2(grid_clb_5_ccff_tail),
        .chanx_left_in(sb_0__1__5_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__12_chanx_left_out),
        .chany_bottom_in(sb_1__1__4_chany_top_out),
        .chany_top_in_0(cby_1__1__6_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[14]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[50]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_5_ccff_tail),
        .ccff_tail_0(cbx_1__1__5_ccff_tail),
        .chanx_left_out(cbx_1__1__5_chanx_left_out),
        .chanx_right_out_0(sb_1__1__5_chanx_right_out),
        .chany_bottom_out(cby_1__1__5_chany_bottom_out),
        .chany_top_out_0(sb_1__1__5_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[15]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[51]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_2__8_
    (
        .ccff_head_1(cbx_1__1__5_ccff_tail),
        .ccff_head_2(grid_clb_15_ccff_tail),
        .chanx_left_in(sb_0__1__6_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__13_chanx_left_out),
        .chany_bottom_in(sb_1__1__5_chany_top_out),
        .chany_top_in_0(cby_1__1__7_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[15]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[51]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_6_ccff_tail),
        .ccff_tail_0(cbx_1__1__6_ccff_tail),
        .chanx_left_out(cbx_1__1__6_chanx_left_out),
        .chanx_right_out_0(sb_1__1__6_chanx_right_out),
        .chany_bottom_out(cby_1__1__6_chany_bottom_out),
        .chany_top_out_0(sb_1__1__6_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    top_tile tile_2__9_
    (
        .ccff_head_1(cbx_1__1__6_ccff_tail),
        .ccff_head_2(grid_io_top_top_1_ccff_tail),
        .chanx_left_in(sb_0__8__0_chanx_right_out),
        .chanx_right_in_0(cbx_1__8__1_chanx_left_out),
        .chany_bottom_in(sb_1__1__6_chany_top_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[0:3]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_7_),
        .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .scan_enable(scan_enable),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_1__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_1__8__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(ccff_tail),
        .ccff_tail_0(grid_io_top_top_0_ccff_tail),
        .chanx_left_out(cbx_1__8__0_chanx_left_out),
        .chanx_right_out_0(sb_1__8__0_chanx_right_out),
        .chany_bottom_out(cby_1__1__7_chany_bottom_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[0:3]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[0:3]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    bottom_tile tile_3__1_
    (
        .ccff_head(grid_io_bottom_bottom_7_ccff_tail),
        .ccff_head_1(grid_clb_0_ccff_tail),
        .chanx_left_in(sb_1__0__0_chanx_right_out),
        .chanx_right_in_0(cbx_1__0__2_chanx_left_out),
        .chany_top_in(cby_1__1__8_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[88:91]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_top_in(prog_reset_ft[20]),
        .reset_top_in(reset_ft[47]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
        .ccff_tail(grid_io_bottom_bottom_6_ccff_tail),
        .ccff_tail_0(cbx_1__0__1_ccff_tail),
        .chanx_left_out(cbx_1__0__1_chanx_left_out),
        .chanx_right_out_0(sb_1__0__1_chanx_right_out),
        .chany_top_out(sb_1__0__1_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[88:91]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[88:91]),
        .top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    tile tile_3__2_
    (
        .ccff_head_1(cbx_1__0__1_ccff_tail),
        .ccff_head_2(grid_clb_17_ccff_tail),
        .chanx_left_in(sb_1__1__0_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__14_chanx_left_out),
        .chany_bottom_in(sb_1__0__1_chany_top_out),
        .chany_top_in_0(cby_1__1__9_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[19]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[46]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_8_ccff_tail),
        .ccff_tail_0(cbx_1__1__7_ccff_tail),
        .chanx_left_out(cbx_1__1__7_chanx_left_out),
        .chanx_right_out_0(sb_1__1__7_chanx_right_out),
        .chany_bottom_out(cby_1__1__8_chany_bottom_out),
        .chany_top_out_0(sb_1__1__7_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[20]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[47]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_3__3_
    (
        .ccff_head_1(cbx_1__1__7_ccff_tail),
        .ccff_head_2(grid_clb_2_ccff_tail),
        .chanx_left_in(sb_1__1__1_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__15_chanx_left_out),
        .chany_bottom_in(sb_1__1__7_chany_top_out),
        .chany_top_in_0(cby_1__1__10_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[18]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[45]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_9_ccff_tail),
        .ccff_tail_0(cbx_1__1__8_ccff_tail),
        .chanx_left_out(cbx_1__1__8_chanx_left_out),
        .chanx_right_out_0(sb_1__1__8_chanx_right_out),
        .chany_bottom_out(cby_1__1__9_chany_bottom_out),
        .chany_top_out_0(sb_1__1__8_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[19]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[46]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_3__4_
    (
        .ccff_head_1(cbx_1__1__8_ccff_tail),
        .ccff_head_2(grid_clb_19_ccff_tail),
        .chanx_left_in(sb_1__1__2_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__16_chanx_left_out),
        .chany_bottom_in(sb_1__1__8_chany_top_out),
        .chany_top_in_0(cby_1__1__11_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[17]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[44]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_10_ccff_tail),
        .ccff_tail_0(cbx_1__1__9_ccff_tail),
        .chanx_left_out(cbx_1__1__9_chanx_left_out),
        .chanx_right_out_0(sb_1__1__9_chanx_right_out),
        .chany_bottom_out(cby_1__1__10_chany_bottom_out),
        .chany_top_out_0(sb_1__1__9_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[18]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[45]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_3__5_
    (
        .ccff_head_1(cbx_1__1__9_ccff_tail),
        .ccff_head_2(grid_clb_4_ccff_tail),
        .chanx_left_in(sb_1__1__3_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__17_chanx_left_out),
        .chany_bottom_in(sb_1__1__9_chany_top_out),
        .chany_top_in_0(cby_1__1__12_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(prog_reset_ft[16]),
        .prog_reset_top_in(),
        .reset_bottom_in(),
        .reset_right_in(reset_ft[40]),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_11_ccff_tail),
        .ccff_tail_0(cbx_1__1__10_ccff_tail),
        .chanx_left_out(cbx_1__1__10_chanx_left_out),
        .chanx_right_out_0(sb_1__1__10_chanx_right_out),
        .chany_bottom_out(cby_1__1__11_chany_bottom_out),
        .chany_top_out_0(sb_1__1__10_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[17]),
        .prog_reset_right_out(prog_reset_ft[24]),
        .prog_reset_top_out(prog_reset_ft[21]),
        .reset_bottom_out(reset_ft[44]),
        .reset_left_out(reset_ft[48]),
        .reset_top_out(reset_ft[41]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_3__6_
    (
        .ccff_head_1(cbx_1__1__10_ccff_tail),
        .ccff_head_2(grid_clb_21_ccff_tail),
        .chanx_left_in(sb_1__1__4_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__18_chanx_left_out),
        .chany_bottom_in(sb_1__1__10_chany_top_out),
        .chany_top_in_0(cby_1__1__13_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[21]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[41]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_12_ccff_tail),
        .ccff_tail_0(cbx_1__1__11_ccff_tail),
        .chanx_left_out(cbx_1__1__11_chanx_left_out),
        .chanx_right_out_0(sb_1__1__11_chanx_right_out),
        .chany_bottom_out(cby_1__1__12_chany_bottom_out),
        .chany_top_out_0(sb_1__1__11_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[22]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[42]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_3__7_
    (
        .ccff_head_1(cbx_1__1__11_ccff_tail),
        .ccff_head_2(grid_clb_6_ccff_tail),
        .chanx_left_in(sb_1__1__5_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__19_chanx_left_out),
        .chany_bottom_in(sb_1__1__11_chany_top_out),
        .chany_top_in_0(cby_1__1__14_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[22]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[42]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_13_ccff_tail),
        .ccff_tail_0(cbx_1__1__12_ccff_tail),
        .chanx_left_out(cbx_1__1__12_chanx_left_out),
        .chanx_right_out_0(sb_1__1__12_chanx_right_out),
        .chany_bottom_out(cby_1__1__13_chany_bottom_out),
        .chany_top_out_0(sb_1__1__12_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[23]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[43]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_3__8_
    (
        .ccff_head_1(cbx_1__1__12_ccff_tail),
        .ccff_head_2(grid_clb_23_ccff_tail),
        .chanx_left_in(sb_1__1__6_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__20_chanx_left_out),
        .chany_bottom_in(sb_1__1__12_chany_top_out),
        .chany_top_in_0(cby_1__1__15_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[23]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[43]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_14_ccff_tail),
        .ccff_tail_0(cbx_1__1__13_ccff_tail),
        .chanx_left_out(cbx_1__1__13_chanx_left_out),
        .chanx_right_out_0(sb_1__1__13_chanx_right_out),
        .chany_bottom_out(cby_1__1__14_chany_bottom_out),
        .chany_top_out_0(sb_1__1__13_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    top_tile tile_3__9_
    (
        .ccff_head_1(cbx_1__1__13_ccff_tail),
        .ccff_head_2(grid_io_top_top_2_ccff_tail),
        .chanx_left_in(sb_1__8__0_chanx_right_out),
        .chanx_right_in_0(cbx_1__8__2_chanx_left_out),
        .chany_bottom_in(sb_1__1__13_chany_top_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[4:7]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_7_),
        .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .scan_enable(scan_enable),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_2__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_2__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_clb_15_ccff_tail),
        .ccff_tail_0(grid_io_top_top_1_ccff_tail),
        .chanx_left_out(cbx_1__8__1_chanx_left_out),
        .chanx_right_out_0(sb_1__8__1_chanx_right_out),
        .chany_bottom_out(cby_1__1__15_chany_bottom_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[4:7]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[4:7]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    bottom_tile tile_4__1_
    (
        .ccff_head(grid_io_bottom_bottom_6_ccff_tail),
        .ccff_head_1(grid_clb_8_ccff_tail),
        .chanx_left_in(sb_1__0__1_chanx_right_out),
        .chanx_right_in_0(cbx_1__0__3_chanx_left_out),
        .chany_top_in(cby_1__1__16_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[84:87]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_top_in(prog_reset_ft[28]),
        .reset_top_in(reset_ft[39]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_),
        .ccff_tail(grid_io_bottom_bottom_5_ccff_tail),
        .ccff_tail_0(cbx_1__0__2_ccff_tail),
        .chanx_left_out(cbx_1__0__2_chanx_left_out),
        .chanx_right_out_0(sb_1__0__2_chanx_right_out),
        .chany_top_out(sb_1__0__2_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[84:87]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[84:87]),
        .top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    tile tile_4__2_
    (
        .ccff_head_1(cbx_1__0__2_ccff_tail),
        .ccff_head_2(grid_clb_25_ccff_tail),
        .chanx_left_in(sb_1__1__7_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__21_chanx_left_out),
        .chany_bottom_in(sb_1__0__2_chany_top_out),
        .chany_top_in_0(cby_1__1__17_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[27]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[38]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_16_ccff_tail),
        .ccff_tail_0(cbx_1__1__14_ccff_tail),
        .chanx_left_out(cbx_1__1__14_chanx_left_out),
        .chanx_right_out_0(sb_1__1__14_chanx_right_out),
        .chany_bottom_out(cby_1__1__16_chany_bottom_out),
        .chany_top_out_0(sb_1__1__14_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[28]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[39]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_4__3_
    (
        .ccff_head_1(cbx_1__1__14_ccff_tail),
        .ccff_head_2(grid_clb_10_ccff_tail),
        .chanx_left_in(sb_1__1__8_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__22_chanx_left_out),
        .chany_bottom_in(sb_1__1__14_chany_top_out),
        .chany_top_in_0(cby_1__1__18_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[26]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[37]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_17_ccff_tail),
        .ccff_tail_0(cbx_1__1__15_ccff_tail),
        .chanx_left_out(cbx_1__1__15_chanx_left_out),
        .chanx_right_out_0(sb_1__1__15_chanx_right_out),
        .chany_bottom_out(cby_1__1__17_chany_bottom_out),
        .chany_top_out_0(sb_1__1__15_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[27]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[38]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_4__4_
    (
        .ccff_head_1(cbx_1__1__15_ccff_tail),
        .ccff_head_2(grid_clb_27_ccff_tail),
        .chanx_left_in(sb_1__1__9_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__23_chanx_left_out),
        .chany_bottom_in(sb_1__1__15_chany_top_out),
        .chany_top_in_0(cby_1__1__19_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[25]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[36]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_18_ccff_tail),
        .ccff_tail_0(cbx_1__1__16_ccff_tail),
        .chanx_left_out(cbx_1__1__16_chanx_left_out),
        .chanx_right_out_0(sb_1__1__16_chanx_right_out),
        .chany_bottom_out(cby_1__1__18_chany_bottom_out),
        .chany_top_out_0(sb_1__1__16_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[26]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[37]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_4__5_
    (
        .ccff_head_1(cbx_1__1__16_ccff_tail),
        .ccff_head_2(grid_clb_12_ccff_tail),
        .chanx_left_in(sb_1__1__10_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__24_chanx_left_out),
        .chany_bottom_in(sb_1__1__16_chany_top_out),
        .chany_top_in_0(cby_1__1__20_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(prog_reset_ft[24]),
        .prog_reset_top_in(),
        .reset_bottom_in(),
        .reset_right_in(reset_ft[32]),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_19_ccff_tail),
        .ccff_tail_0(cbx_1__1__17_ccff_tail),
        .chanx_left_out(cbx_1__1__17_chanx_left_out),
        .chanx_right_out_0(sb_1__1__17_chanx_right_out),
        .chany_bottom_out(cby_1__1__19_chany_bottom_out),
        .chany_top_out_0(sb_1__1__17_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[25]),
        .prog_reset_right_out(prog_reset_ft[32]),
        .prog_reset_top_out(prog_reset_ft[29]),
        .reset_bottom_out(reset_ft[36]),
        .reset_left_out(reset_ft[40]),
        .reset_top_out(reset_ft[33]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_4__6_
    (
        .ccff_head_1(cbx_1__1__17_ccff_tail),
        .ccff_head_2(grid_clb_29_ccff_tail),
        .chanx_left_in(sb_1__1__11_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__25_chanx_left_out),
        .chany_bottom_in(sb_1__1__17_chany_top_out),
        .chany_top_in_0(cby_1__1__21_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[29]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[33]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_20_ccff_tail),
        .ccff_tail_0(cbx_1__1__18_ccff_tail),
        .chanx_left_out(cbx_1__1__18_chanx_left_out),
        .chanx_right_out_0(sb_1__1__18_chanx_right_out),
        .chany_bottom_out(cby_1__1__20_chany_bottom_out),
        .chany_top_out_0(sb_1__1__18_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[30]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[34]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_4__7_
    (
        .ccff_head_1(cbx_1__1__18_ccff_tail),
        .ccff_head_2(grid_clb_14_ccff_tail),
        .chanx_left_in(sb_1__1__12_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__26_chanx_left_out),
        .chany_bottom_in(sb_1__1__18_chany_top_out),
        .chany_top_in_0(cby_1__1__22_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[30]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[34]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_21_ccff_tail),
        .ccff_tail_0(cbx_1__1__19_ccff_tail),
        .chanx_left_out(cbx_1__1__19_chanx_left_out),
        .chanx_right_out_0(sb_1__1__19_chanx_right_out),
        .chany_bottom_out(cby_1__1__21_chany_bottom_out),
        .chany_top_out_0(sb_1__1__19_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[31]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[35]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_4__8_
    (
        .ccff_head_1(cbx_1__1__19_ccff_tail),
        .ccff_head_2(grid_clb_31_ccff_tail),
        .chanx_left_in(sb_1__1__13_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__27_chanx_left_out),
        .chany_bottom_in(sb_1__1__19_chany_top_out),
        .chany_top_in_0(cby_1__1__23_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[31]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[35]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_22_ccff_tail),
        .ccff_tail_0(cbx_1__1__20_ccff_tail),
        .chanx_left_out(cbx_1__1__20_chanx_left_out),
        .chanx_right_out_0(sb_1__1__20_chanx_right_out),
        .chany_bottom_out(cby_1__1__22_chany_bottom_out),
        .chany_top_out_0(sb_1__1__20_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    top_tile tile_4__9_
    (
        .ccff_head_1(cbx_1__1__20_ccff_tail),
        .ccff_head_2(grid_io_top_top_3_ccff_tail),
        .chanx_left_in(sb_1__8__1_chanx_right_out),
        .chanx_right_in_0(cbx_1__8__3_chanx_left_out),
        .chany_bottom_in(sb_1__1__20_chany_top_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[8:11]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_7_),
        .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .scan_enable(scan_enable),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_3__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_clb_23_ccff_tail),
        .ccff_tail_0(grid_io_top_top_2_ccff_tail),
        .chanx_left_out(cbx_1__8__2_chanx_left_out),
        .chanx_right_out_0(sb_1__8__2_chanx_right_out),
        .chany_bottom_out(cby_1__1__23_chany_bottom_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[8:11]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[8:11]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    bottom_tile tile_5__1_
    (
        .ccff_head(grid_io_bottom_bottom_5_ccff_tail),
        .ccff_head_1(grid_clb_16_ccff_tail),
        .chanx_left_in(sb_1__0__2_chanx_right_out),
        .chanx_right_in_0(cbx_1__0__4_chanx_left_out),
        .chany_top_in(cby_1__1__24_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[80:83]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_top_in(prog_reset_ft[36]),
        .reset_top_in(reset_ft[31]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_),
        .ccff_tail(grid_io_bottom_bottom_4_ccff_tail),
        .ccff_tail_0(cbx_1__0__3_ccff_tail),
        .chanx_left_out(cbx_1__0__3_chanx_left_out),
        .chanx_right_out_0(sb_1__0__3_chanx_right_out),
        .chany_top_out(sb_1__0__3_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[80:83]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[80:83]),
        .top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    tile tile_5__2_
    (
        .ccff_head_1(cbx_1__0__3_ccff_tail),
        .ccff_head_2(grid_clb_33_ccff_tail),
        .chanx_left_in(sb_1__1__14_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__28_chanx_left_out),
        .chany_bottom_in(sb_1__0__3_chany_top_out),
        .chany_top_in_0(cby_1__1__25_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[35]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[30]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_24_ccff_tail),
        .ccff_tail_0(cbx_1__1__21_ccff_tail),
        .chanx_left_out(cbx_1__1__21_chanx_left_out),
        .chanx_right_out_0(sb_1__1__21_chanx_right_out),
        .chany_bottom_out(cby_1__1__24_chany_bottom_out),
        .chany_top_out_0(sb_1__1__21_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[36]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[31]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_5__3_
    (
        .ccff_head_1(cbx_1__1__21_ccff_tail),
        .ccff_head_2(grid_clb_18_ccff_tail),
        .chanx_left_in(sb_1__1__15_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__29_chanx_left_out),
        .chany_bottom_in(sb_1__1__21_chany_top_out),
        .chany_top_in_0(cby_1__1__26_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[34]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[29]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_25_ccff_tail),
        .ccff_tail_0(cbx_1__1__22_ccff_tail),
        .chanx_left_out(cbx_1__1__22_chanx_left_out),
        .chanx_right_out_0(sb_1__1__22_chanx_right_out),
        .chany_bottom_out(cby_1__1__25_chany_bottom_out),
        .chany_top_out_0(sb_1__1__22_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[35]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[30]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_5__4_
    (
        .ccff_head_1(cbx_1__1__22_ccff_tail),
        .ccff_head_2(grid_clb_35_ccff_tail),
        .chanx_left_in(sb_1__1__16_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__30_chanx_left_out),
        .chany_bottom_in(sb_1__1__22_chany_top_out),
        .chany_top_in_0(cby_1__1__27_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[33]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[28]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_26_ccff_tail),
        .ccff_tail_0(cbx_1__1__23_ccff_tail),
        .chanx_left_out(cbx_1__1__23_chanx_left_out),
        .chanx_right_out_0(sb_1__1__23_chanx_right_out),
        .chany_bottom_out(cby_1__1__26_chany_bottom_out),
        .chany_top_out_0(sb_1__1__23_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[34]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[29]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_5__5_
    (
        .ccff_head_1(cbx_1__1__23_ccff_tail),
        .ccff_head_2(grid_clb_20_ccff_tail),
        .chanx_left_in(sb_1__1__17_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__31_chanx_left_out),
        .chany_bottom_in(sb_1__1__23_chany_top_out),
        .chany_top_in_0(cby_1__1__28_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(prog_reset_ft[32]),
        .prog_reset_top_in(),
        .reset_bottom_in(),
        .reset_right_in(reset_ft[24]),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_27_ccff_tail),
        .ccff_tail_0(cbx_1__1__24_ccff_tail),
        .chanx_left_out(cbx_1__1__24_chanx_left_out),
        .chanx_right_out_0(sb_1__1__24_chanx_right_out),
        .chany_bottom_out(cby_1__1__27_chany_bottom_out),
        .chany_top_out_0(sb_1__1__24_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[33]),
        .prog_reset_right_out(prog_reset_ft[40]),
        .prog_reset_top_out(prog_reset_ft[37]),
        .reset_bottom_out(reset_ft[28]),
        .reset_left_out(reset_ft[32]),
        .reset_top_out(reset_ft[25]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_5__6_
    (
        .ccff_head_1(cbx_1__1__24_ccff_tail),
        .ccff_head_2(grid_clb_37_ccff_tail),
        .chanx_left_in(sb_1__1__18_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__32_chanx_left_out),
        .chany_bottom_in(sb_1__1__24_chany_top_out),
        .chany_top_in_0(cby_1__1__29_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[37]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[25]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_28_ccff_tail),
        .ccff_tail_0(cbx_1__1__25_ccff_tail),
        .chanx_left_out(cbx_1__1__25_chanx_left_out),
        .chanx_right_out_0(sb_1__1__25_chanx_right_out),
        .chany_bottom_out(cby_1__1__28_chany_bottom_out),
        .chany_top_out_0(sb_1__1__25_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[38]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[26]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_5__7_
    (
        .ccff_head_1(cbx_1__1__25_ccff_tail),
        .ccff_head_2(grid_clb_22_ccff_tail),
        .chanx_left_in(sb_1__1__19_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__33_chanx_left_out),
        .chany_bottom_in(sb_1__1__25_chany_top_out),
        .chany_top_in_0(cby_1__1__30_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[38]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[26]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_29_ccff_tail),
        .ccff_tail_0(cbx_1__1__26_ccff_tail),
        .chanx_left_out(cbx_1__1__26_chanx_left_out),
        .chanx_right_out_0(sb_1__1__26_chanx_right_out),
        .chany_bottom_out(cby_1__1__29_chany_bottom_out),
        .chany_top_out_0(sb_1__1__26_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[39]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[27]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_5__8_
    (
        .ccff_head_1(cbx_1__1__26_ccff_tail),
        .ccff_head_2(grid_clb_39_ccff_tail),
        .chanx_left_in(sb_1__1__20_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__34_chanx_left_out),
        .chany_bottom_in(sb_1__1__26_chany_top_out),
        .chany_top_in_0(cby_1__1__31_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[39]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[27]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_30_ccff_tail),
        .ccff_tail_0(cbx_1__1__27_ccff_tail),
        .chanx_left_out(cbx_1__1__27_chanx_left_out),
        .chanx_right_out_0(sb_1__1__27_chanx_right_out),
        .chany_bottom_out(cby_1__1__30_chany_bottom_out),
        .chany_top_out_0(sb_1__1__27_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    top_tile tile_5__9_
    (
        .ccff_head_1(cbx_1__1__27_ccff_tail),
        .ccff_head_2(grid_io_top_top_4_ccff_tail),
        .chanx_left_in(sb_1__8__2_chanx_right_out),
        .chanx_right_in_0(cbx_1__8__4_chanx_left_out),
        .chany_bottom_in(sb_1__1__27_chany_top_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[12:15]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_7_),
        .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .scan_enable(scan_enable),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_4__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_4__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_clb_31_ccff_tail),
        .ccff_tail_0(grid_io_top_top_3_ccff_tail),
        .chanx_left_out(cbx_1__8__3_chanx_left_out),
        .chanx_right_out_0(sb_1__8__3_chanx_right_out),
        .chany_bottom_out(cby_1__1__31_chany_bottom_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[12:15]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[12:15]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    bottom_tile tile_6__1_
    (
        .ccff_head(grid_io_bottom_bottom_4_ccff_tail),
        .ccff_head_1(grid_clb_24_ccff_tail),
        .chanx_left_in(sb_1__0__3_chanx_right_out),
        .chanx_right_in_0(cbx_1__0__5_chanx_left_out),
        .chany_top_in(cby_1__1__32_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[76:79]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_top_in(prog_reset_ft[44]),
        .reset_top_in(reset_ft[23]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_),
        .ccff_tail(grid_io_bottom_bottom_3_ccff_tail),
        .ccff_tail_0(cbx_1__0__4_ccff_tail),
        .chanx_left_out(cbx_1__0__4_chanx_left_out),
        .chanx_right_out_0(sb_1__0__4_chanx_right_out),
        .chany_top_out(sb_1__0__4_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[76:79]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[76:79]),
        .top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    tile tile_6__2_
    (
        .ccff_head_1(cbx_1__0__4_ccff_tail),
        .ccff_head_2(grid_clb_41_ccff_tail),
        .chanx_left_in(sb_1__1__21_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__35_chanx_left_out),
        .chany_bottom_in(sb_1__0__4_chany_top_out),
        .chany_top_in_0(cby_1__1__33_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[43]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[22]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_32_ccff_tail),
        .ccff_tail_0(cbx_1__1__28_ccff_tail),
        .chanx_left_out(cbx_1__1__28_chanx_left_out),
        .chanx_right_out_0(sb_1__1__28_chanx_right_out),
        .chany_bottom_out(cby_1__1__32_chany_bottom_out),
        .chany_top_out_0(sb_1__1__28_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[44]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[23]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_6__3_
    (
        .ccff_head_1(cbx_1__1__28_ccff_tail),
        .ccff_head_2(grid_clb_26_ccff_tail),
        .chanx_left_in(sb_1__1__22_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__36_chanx_left_out),
        .chany_bottom_in(sb_1__1__28_chany_top_out),
        .chany_top_in_0(cby_1__1__34_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[42]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[21]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_33_ccff_tail),
        .ccff_tail_0(cbx_1__1__29_ccff_tail),
        .chanx_left_out(cbx_1__1__29_chanx_left_out),
        .chanx_right_out_0(sb_1__1__29_chanx_right_out),
        .chany_bottom_out(cby_1__1__33_chany_bottom_out),
        .chany_top_out_0(sb_1__1__29_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[43]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[22]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_6__4_
    (
        .ccff_head_1(cbx_1__1__29_ccff_tail),
        .ccff_head_2(grid_clb_43_ccff_tail),
        .chanx_left_in(sb_1__1__23_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__37_chanx_left_out),
        .chany_bottom_in(sb_1__1__29_chany_top_out),
        .chany_top_in_0(cby_1__1__35_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[41]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[20]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_34_ccff_tail),
        .ccff_tail_0(cbx_1__1__30_ccff_tail),
        .chanx_left_out(cbx_1__1__30_chanx_left_out),
        .chanx_right_out_0(sb_1__1__30_chanx_right_out),
        .chany_bottom_out(cby_1__1__34_chany_bottom_out),
        .chany_top_out_0(sb_1__1__30_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[42]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[21]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_6__5_
    (
        .ccff_head_1(cbx_1__1__30_ccff_tail),
        .ccff_head_2(grid_clb_28_ccff_tail),
        .chanx_left_in(sb_1__1__24_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__38_chanx_left_out),
        .chany_bottom_in(sb_1__1__30_chany_top_out),
        .chany_top_in_0(cby_1__1__36_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(prog_reset_ft[40]),
        .prog_reset_top_in(),
        .reset_bottom_in(),
        .reset_right_in(reset_ft[16]),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_35_ccff_tail),
        .ccff_tail_0(cbx_1__1__31_ccff_tail),
        .chanx_left_out(cbx_1__1__31_chanx_left_out),
        .chanx_right_out_0(sb_1__1__31_chanx_right_out),
        .chany_bottom_out(cby_1__1__35_chany_bottom_out),
        .chany_top_out_0(sb_1__1__31_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[41]),
        .prog_reset_right_out(prog_reset_ft[48]),
        .prog_reset_top_out(prog_reset_ft[45]),
        .reset_bottom_out(reset_ft[20]),
        .reset_left_out(reset_ft[24]),
        .reset_top_out(reset_ft[17]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_6__6_
    (
        .ccff_head_1(cbx_1__1__31_ccff_tail),
        .ccff_head_2(grid_clb_45_ccff_tail),
        .chanx_left_in(sb_1__1__25_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__39_chanx_left_out),
        .chany_bottom_in(sb_1__1__31_chany_top_out),
        .chany_top_in_0(cby_1__1__37_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[45]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[17]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_36_ccff_tail),
        .ccff_tail_0(cbx_1__1__32_ccff_tail),
        .chanx_left_out(cbx_1__1__32_chanx_left_out),
        .chanx_right_out_0(sb_1__1__32_chanx_right_out),
        .chany_bottom_out(cby_1__1__36_chany_bottom_out),
        .chany_top_out_0(sb_1__1__32_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[46]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[18]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_6__7_
    (
        .ccff_head_1(cbx_1__1__32_ccff_tail),
        .ccff_head_2(grid_clb_30_ccff_tail),
        .chanx_left_in(sb_1__1__26_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__40_chanx_left_out),
        .chany_bottom_in(sb_1__1__32_chany_top_out),
        .chany_top_in_0(cby_1__1__38_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[46]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[18]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_37_ccff_tail),
        .ccff_tail_0(cbx_1__1__33_ccff_tail),
        .chanx_left_out(cbx_1__1__33_chanx_left_out),
        .chanx_right_out_0(sb_1__1__33_chanx_right_out),
        .chany_bottom_out(cby_1__1__37_chany_bottom_out),
        .chany_top_out_0(sb_1__1__33_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[47]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[19]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_6__8_
    (
        .ccff_head_1(cbx_1__1__33_ccff_tail),
        .ccff_head_2(grid_clb_47_ccff_tail),
        .chanx_left_in(sb_1__1__27_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__41_chanx_left_out),
        .chany_bottom_in(sb_1__1__33_chany_top_out),
        .chany_top_in_0(cby_1__1__39_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[47]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[19]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_38_ccff_tail),
        .ccff_tail_0(cbx_1__1__34_ccff_tail),
        .chanx_left_out(cbx_1__1__34_chanx_left_out),
        .chanx_right_out_0(sb_1__1__34_chanx_right_out),
        .chany_bottom_out(cby_1__1__38_chany_bottom_out),
        .chany_top_out_0(sb_1__1__34_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    top_tile tile_6__9_
    (
        .ccff_head_1(cbx_1__1__34_ccff_tail),
        .ccff_head_2(grid_io_top_top_5_ccff_tail),
        .chanx_left_in(sb_1__8__3_chanx_right_out),
        .chanx_right_in_0(cbx_1__8__5_chanx_left_out),
        .chany_bottom_in(sb_1__1__34_chany_top_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[16:19]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_7_),
        .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .scan_enable(scan_enable),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_5__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_clb_39_ccff_tail),
        .ccff_tail_0(grid_io_top_top_4_ccff_tail),
        .chanx_left_out(cbx_1__8__4_chanx_left_out),
        .chanx_right_out_0(sb_1__8__4_chanx_right_out),
        .chany_bottom_out(cby_1__1__39_chany_bottom_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[16:19]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[16:19]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    bottom_tile tile_7__1_
    (
        .ccff_head(grid_io_bottom_bottom_3_ccff_tail),
        .ccff_head_1(grid_clb_32_ccff_tail),
        .chanx_left_in(sb_1__0__4_chanx_right_out),
        .chanx_right_in_0(cbx_1__0__6_chanx_left_out),
        .chany_top_in(cby_1__1__40_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[72:75]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_top_in(prog_reset_ft[52]),
        .reset_top_in(reset_ft[15]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_),
        .ccff_tail(grid_io_bottom_bottom_2_ccff_tail),
        .ccff_tail_0(cbx_1__0__5_ccff_tail),
        .chanx_left_out(cbx_1__0__5_chanx_left_out),
        .chanx_right_out_0(sb_1__0__5_chanx_right_out),
        .chany_top_out(sb_1__0__5_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[72:75]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[72:75]),
        .top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    tile tile_7__2_
    (
        .ccff_head_1(cbx_1__0__5_ccff_tail),
        .ccff_head_2(grid_clb_49_ccff_tail),
        .chanx_left_in(sb_1__1__28_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__42_chanx_left_out),
        .chany_bottom_in(sb_1__0__5_chany_top_out),
        .chany_top_in_0(cby_1__1__41_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[51]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[14]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_6__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_6__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_40_ccff_tail),
        .ccff_tail_0(cbx_1__1__35_ccff_tail),
        .chanx_left_out(cbx_1__1__35_chanx_left_out),
        .chanx_right_out_0(sb_1__1__35_chanx_right_out),
        .chany_bottom_out(cby_1__1__40_chany_bottom_out),
        .chany_top_out_0(sb_1__1__35_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[52]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[15]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_7__3_
    (
        .ccff_head_1(cbx_1__1__35_ccff_tail),
        .ccff_head_2(grid_clb_34_ccff_tail),
        .chanx_left_in(sb_1__1__29_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__43_chanx_left_out),
        .chany_bottom_in(sb_1__1__35_chany_top_out),
        .chany_top_in_0(cby_1__1__42_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[50]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[13]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_41_ccff_tail),
        .ccff_tail_0(cbx_1__1__36_ccff_tail),
        .chanx_left_out(cbx_1__1__36_chanx_left_out),
        .chanx_right_out_0(sb_1__1__36_chanx_right_out),
        .chany_bottom_out(cby_1__1__41_chany_bottom_out),
        .chany_top_out_0(sb_1__1__36_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[51]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[14]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_7__4_
    (
        .ccff_head_1(cbx_1__1__36_ccff_tail),
        .ccff_head_2(grid_clb_51_ccff_tail),
        .chanx_left_in(sb_1__1__30_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__44_chanx_left_out),
        .chany_bottom_in(sb_1__1__36_chany_top_out),
        .chany_top_in_0(cby_1__1__43_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[49]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[12]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_42_ccff_tail),
        .ccff_tail_0(cbx_1__1__37_ccff_tail),
        .chanx_left_out(cbx_1__1__37_chanx_left_out),
        .chanx_right_out_0(sb_1__1__37_chanx_right_out),
        .chany_bottom_out(cby_1__1__42_chany_bottom_out),
        .chany_top_out_0(sb_1__1__37_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[50]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[13]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_7__5_
    (
        .ccff_head_1(cbx_1__1__37_ccff_tail),
        .ccff_head_2(grid_clb_36_ccff_tail),
        .chanx_left_in(sb_1__1__31_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__45_chanx_left_out),
        .chany_bottom_in(sb_1__1__37_chany_top_out),
        .chany_top_in_0(cby_1__1__44_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(prog_reset_ft[48]),
        .prog_reset_top_in(),
        .reset_bottom_in(),
        .reset_right_in(reset_ft[8]),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_43_ccff_tail),
        .ccff_tail_0(cbx_1__1__38_ccff_tail),
        .chanx_left_out(cbx_1__1__38_chanx_left_out),
        .chanx_right_out_0(sb_1__1__38_chanx_right_out),
        .chany_bottom_out(cby_1__1__43_chany_bottom_out),
        .chany_top_out_0(sb_1__1__38_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[49]),
        .prog_reset_right_out(prog_reset_ft[56]),
        .prog_reset_top_out(prog_reset_ft[53]),
        .reset_bottom_out(reset_ft[12]),
        .reset_left_out(reset_ft[16]),
        .reset_top_out(reset_ft[9]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_7__6_
    (
        .ccff_head_1(cbx_1__1__38_ccff_tail),
        .ccff_head_2(grid_clb_53_ccff_tail),
        .chanx_left_in(sb_1__1__32_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__46_chanx_left_out),
        .chany_bottom_in(sb_1__1__38_chany_top_out),
        .chany_top_in_0(cby_1__1__45_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[53]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[9]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_44_ccff_tail),
        .ccff_tail_0(cbx_1__1__39_ccff_tail),
        .chanx_left_out(cbx_1__1__39_chanx_left_out),
        .chanx_right_out_0(sb_1__1__39_chanx_right_out),
        .chany_bottom_out(cby_1__1__44_chany_bottom_out),
        .chany_top_out_0(sb_1__1__39_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[54]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[10]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_7__7_
    (
        .ccff_head_1(cbx_1__1__39_ccff_tail),
        .ccff_head_2(grid_clb_38_ccff_tail),
        .chanx_left_in(sb_1__1__33_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__47_chanx_left_out),
        .chany_bottom_in(sb_1__1__39_chany_top_out),
        .chany_top_in_0(cby_1__1__46_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[54]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[10]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_45_ccff_tail),
        .ccff_tail_0(cbx_1__1__40_ccff_tail),
        .chanx_left_out(cbx_1__1__40_chanx_left_out),
        .chanx_right_out_0(sb_1__1__40_chanx_right_out),
        .chany_bottom_out(cby_1__1__45_chany_bottom_out),
        .chany_top_out_0(sb_1__1__40_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[55]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[11]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_7__8_
    (
        .ccff_head_1(cbx_1__1__40_ccff_tail),
        .ccff_head_2(grid_clb_55_ccff_tail),
        .chanx_left_in(sb_1__1__34_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__48_chanx_left_out),
        .chany_bottom_in(sb_1__1__40_chany_top_out),
        .chany_top_in_0(cby_1__1__47_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[55]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[11]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_46_ccff_tail),
        .ccff_tail_0(cbx_1__1__41_ccff_tail),
        .chanx_left_out(cbx_1__1__41_chanx_left_out),
        .chanx_right_out_0(sb_1__1__41_chanx_right_out),
        .chany_bottom_out(cby_1__1__46_chany_bottom_out),
        .chany_top_out_0(sb_1__1__41_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    top_tile tile_7__9_
    (
        .ccff_head_1(cbx_1__1__41_ccff_tail),
        .ccff_head_2(grid_io_top_top_6_ccff_tail),
        .chanx_left_in(sb_1__8__4_chanx_right_out),
        .chanx_right_in_0(cbx_1__8__6_chanx_left_out),
        .chany_bottom_in(sb_1__1__41_chany_top_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[20:23]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_7_),
        .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .scan_enable(scan_enable),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_6__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_6__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_clb_47_ccff_tail),
        .ccff_tail_0(grid_io_top_top_5_ccff_tail),
        .chanx_left_out(cbx_1__8__5_chanx_left_out),
        .chanx_right_out_0(sb_1__8__5_chanx_right_out),
        .chany_bottom_out(cby_1__1__47_chany_bottom_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[20:23]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[20:23]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    bottom_tile tile_8__1_
    (
        .ccff_head(grid_io_bottom_bottom_2_ccff_tail),
        .ccff_head_1(grid_clb_40_ccff_tail),
        .chanx_left_in(sb_1__0__5_chanx_right_out),
        .chanx_right_in_0(cbx_1__0__7_chanx_left_out),
        .chany_top_in(cby_1__1__48_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[68:71]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset_top_in(prog_reset_ft[60]),
        .reset_top_in(reset_ft[7]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_),
        .ccff_tail(grid_io_bottom_bottom_1_ccff_tail),
        .ccff_tail_0(cbx_1__0__6_ccff_tail),
        .chanx_left_out(cbx_1__0__6_chanx_left_out),
        .chanx_right_out_0(sb_1__0__6_chanx_right_out),
        .chany_top_out(sb_1__0__6_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[68:71]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[68:71]),
        .top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    tile tile_8__2_
    (
        .ccff_head_1(cbx_1__0__6_ccff_tail),
        .ccff_head_2(grid_clb_57_ccff_tail),
        .chanx_left_in(sb_1__1__35_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__49_chanx_left_out),
        .chany_bottom_in(sb_1__0__6_chany_top_out),
        .chany_top_in_0(cby_1__1__49_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[59]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[6]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_48_ccff_tail),
        .ccff_tail_0(cbx_1__1__42_ccff_tail),
        .chanx_left_out(cbx_1__1__42_chanx_left_out),
        .chanx_right_out_0(sb_1__1__42_chanx_right_out),
        .chany_bottom_out(cby_1__1__48_chany_bottom_out),
        .chany_top_out_0(sb_1__1__42_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[60]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[7]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_8__3_
    (
        .ccff_head_1(cbx_1__1__42_ccff_tail),
        .ccff_head_2(grid_clb_42_ccff_tail),
        .chanx_left_in(sb_1__1__36_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__50_chanx_left_out),
        .chany_bottom_in(sb_1__1__42_chany_top_out),
        .chany_top_in_0(cby_1__1__50_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[58]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[5]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_49_ccff_tail),
        .ccff_tail_0(cbx_1__1__43_ccff_tail),
        .chanx_left_out(cbx_1__1__43_chanx_left_out),
        .chanx_right_out_0(sb_1__1__43_chanx_right_out),
        .chany_bottom_out(cby_1__1__49_chany_bottom_out),
        .chany_top_out_0(sb_1__1__43_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[59]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[6]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_8__4_
    (
        .ccff_head_1(cbx_1__1__43_ccff_tail),
        .ccff_head_2(grid_clb_59_ccff_tail),
        .chanx_left_in(sb_1__1__37_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__51_chanx_left_out),
        .chany_bottom_in(sb_1__1__43_chany_top_out),
        .chany_top_in_0(cby_1__1__51_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(),
        .prog_reset_top_in(prog_reset_ft[57]),
        .reset_bottom_in(),
        .reset_right_in(),
        .reset_top_in(reset_ft[4]),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_50_ccff_tail),
        .ccff_tail_0(cbx_1__1__44_ccff_tail),
        .chanx_left_out(cbx_1__1__44_chanx_left_out),
        .chanx_right_out_0(sb_1__1__44_chanx_right_out),
        .chany_bottom_out(cby_1__1__50_chany_bottom_out),
        .chany_top_out_0(sb_1__1__44_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[58]),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(reset_ft[5]),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_8__5_
    (
        .ccff_head_1(cbx_1__1__44_ccff_tail),
        .ccff_head_2(grid_clb_44_ccff_tail),
        .chanx_left_in(sb_1__1__38_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__52_chanx_left_out),
        .chany_bottom_in(sb_1__1__44_chany_top_out),
        .chany_top_in_0(cby_1__1__52_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(),
        .prog_reset_left_in(prog_reset_ft[56]),
        .prog_reset_top_in(),
        .reset_bottom_in(),
        .reset_right_in(reset_ft[0]),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_51_ccff_tail),
        .ccff_tail_0(cbx_1__1__45_ccff_tail),
        .chanx_left_out(cbx_1__1__45_chanx_left_out),
        .chanx_right_out_0(sb_1__1__45_chanx_right_out),
        .chany_bottom_out(cby_1__1__51_chany_bottom_out),
        .chany_top_out_0(sb_1__1__45_chany_top_out),
        .prog_reset_bottom_out(prog_reset_ft[57]),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[61]),
        .reset_bottom_out(reset_ft[4]),
        .reset_left_out(reset_ft[8]),
        .reset_top_out(reset_ft[1]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_8__6_
    (
        .ccff_head_1(cbx_1__1__45_ccff_tail),
        .ccff_head_2(grid_clb_61_ccff_tail),
        .chanx_left_in(sb_1__1__39_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__53_chanx_left_out),
        .chany_bottom_in(sb_1__1__45_chany_top_out),
        .chany_top_in_0(cby_1__1__53_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[61]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[1]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_52_ccff_tail),
        .ccff_tail_0(cbx_1__1__46_ccff_tail),
        .chanx_left_out(cbx_1__1__46_chanx_left_out),
        .chanx_right_out_0(sb_1__1__46_chanx_right_out),
        .chany_bottom_out(cby_1__1__52_chany_bottom_out),
        .chany_top_out_0(sb_1__1__46_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[62]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[2]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_8__7_
    (
        .ccff_head_1(cbx_1__1__46_ccff_tail),
        .ccff_head_2(grid_clb_46_ccff_tail),
        .chanx_left_in(sb_1__1__40_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__54_chanx_left_out),
        .chany_bottom_in(sb_1__1__46_chany_top_out),
        .chany_top_in_0(cby_1__1__54_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[62]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[2]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_53_ccff_tail),
        .ccff_tail_0(cbx_1__1__47_ccff_tail),
        .chanx_left_out(cbx_1__1__47_chanx_left_out),
        .chanx_right_out_0(sb_1__1__47_chanx_right_out),
        .chany_bottom_out(cby_1__1__53_chany_bottom_out),
        .chany_top_out_0(sb_1__1__47_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(prog_reset_ft[63]),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(reset_ft[3]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    tile tile_8__8_
    (
        .ccff_head_1(cbx_1__1__47_ccff_tail),
        .ccff_head_2(grid_clb_63_ccff_tail),
        .chanx_left_in(sb_1__1__41_chanx_right_out),
        .chanx_right_in_0(cbx_1__1__55_chanx_left_out),
        .chany_bottom_in(sb_1__1__47_chany_top_out),
        .chany_top_in_0(cby_1__1__55_chany_bottom_out),
        .clk0(clk),
        .prog_clk(prog_clk),
        .prog_reset_bottom_in(prog_reset_ft[63]),
        .prog_reset_left_in(),
        .prog_reset_top_in(),
        .reset_bottom_in(reset_ft[3]),
        .reset_right_in(),
        .reset_top_in(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_7_),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_54_ccff_tail),
        .ccff_tail_0(cbx_1__1__48_ccff_tail),
        .chanx_left_out(cbx_1__1__48_chanx_left_out),
        .chanx_right_out_0(sb_1__1__48_chanx_right_out),
        .chany_bottom_out(cby_1__1__54_chany_bottom_out),
        .chany_top_out_0(sb_1__1__48_chany_top_out),
        .prog_reset_bottom_out(),
        .prog_reset_right_out(),
        .prog_reset_top_out(),
        .reset_bottom_out(),
        .reset_left_out(),
        .reset_top_out(),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    top_tile tile_8__9_
    (
        .ccff_head_1(cbx_1__1__48_ccff_tail),
        .ccff_head_2(grid_io_top_top_7_ccff_tail),
        .chanx_left_in(sb_1__8__5_chanx_right_out),
        .chanx_right_in_0(cbx_1__8__7_chanx_left_out),
        .chany_bottom_in(sb_1__1__48_chany_top_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[24:27]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_6_),
        .right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_7_),
        .right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .scan_enable(scan_enable),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_7__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_clb_55_ccff_tail),
        .ccff_tail_0(grid_io_top_top_6_ccff_tail),
        .chanx_left_out(cbx_1__8__6_chanx_left_out),
        .chanx_right_out_0(sb_1__8__6_chanx_right_out),
        .chany_bottom_out(cby_1__1__55_chany_bottom_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[24:27]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[24:27]),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    bottom_right_tile tile_9__1_
    (
        .ccff_head(grid_io_bottom_bottom_1_ccff_tail),
        .ccff_head_1(grid_clb_48_ccff_tail),
        .chanx_left_in(sb_1__0__6_chanx_right_out),
        .chany_top_in(cby_8__1__0_chany_bottom_out),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[64:67]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_io_bottom_bottom_0_ccff_tail),
        .ccff_tail_0(cbx_1__0__7_ccff_tail),
        .chanx_left_out(cbx_1__0__7_chanx_left_out),
        .chany_top_out(sb_8__0__0_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[64:67]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[64:67]),
        .top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_)
    );
    right_tile tile_9__2_
    (
        .ccff_head_0_0(cbx_1__0__7_ccff_tail),
        .ccff_head_1(grid_io_bottom_bottom_0_ccff_tail),
        .ccff_head_2(grid_clb_56_ccff_tail),
        .chanx_left_in(sb_1__1__42_chanx_right_out),
        .chany_bottom_in(sb_8__0__0_chany_top_out),
        .chany_top_in_0(cby_8__1__1_chany_bottom_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[60:63]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_56_ccff_tail),
        .ccff_tail_0(cbx_1__1__49_ccff_tail),
        .ccff_tail_1(grid_io_right_right_7_ccff_tail),
        .chanx_left_out(cbx_1__1__49_chanx_left_out),
        .chany_bottom_out(cby_8__1__0_chany_bottom_out),
        .chany_top_out_0(sb_8__1__0_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[60:63]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[60:63]),
        .left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    right_tile tile_9__3_
    (
        .ccff_head_0_0(cbx_1__1__49_ccff_tail),
        .ccff_head_1(grid_io_right_right_7_ccff_tail),
        .ccff_head_2(grid_clb_50_ccff_tail),
        .chanx_left_in(sb_1__1__43_chanx_right_out),
        .chany_bottom_in(sb_8__1__0_chany_top_out),
        .chany_top_in_0(cby_8__1__2_chany_bottom_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[56:59]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_57_ccff_tail),
        .ccff_tail_0(cbx_1__1__50_ccff_tail),
        .ccff_tail_1(grid_io_right_right_6_ccff_tail),
        .chanx_left_out(cbx_1__1__50_chanx_left_out),
        .chany_bottom_out(cby_8__1__1_chany_bottom_out),
        .chany_top_out_0(sb_8__1__1_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[56:59]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[56:59]),
        .left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    right_tile tile_9__4_
    (
        .ccff_head_0_0(cbx_1__1__50_ccff_tail),
        .ccff_head_1(grid_io_right_right_6_ccff_tail),
        .ccff_head_2(grid_clb_58_ccff_tail),
        .chanx_left_in(sb_1__1__44_chanx_right_out),
        .chany_bottom_in(sb_8__1__1_chany_top_out),
        .chany_top_in_0(cby_8__1__3_chany_bottom_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[52:55]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_58_ccff_tail),
        .ccff_tail_0(cbx_1__1__51_ccff_tail),
        .ccff_tail_1(grid_io_right_right_5_ccff_tail),
        .chanx_left_out(cbx_1__1__51_chanx_left_out),
        .chany_bottom_out(cby_8__1__2_chany_bottom_out),
        .chany_top_out_0(sb_8__1__2_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[52:55]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[52:55]),
        .left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    right_tile tile_9__5_
    (
        .ccff_head_0_0(cbx_1__1__51_ccff_tail),
        .ccff_head_1(grid_io_right_right_5_ccff_tail),
        .ccff_head_2(grid_clb_52_ccff_tail),
        .chanx_left_in(sb_1__1__45_chanx_right_out),
        .chany_bottom_in(sb_8__1__2_chany_top_out),
        .chany_top_in_0(cby_8__1__4_chany_bottom_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[48:51]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_59_ccff_tail),
        .ccff_tail_0(cbx_1__1__52_ccff_tail),
        .ccff_tail_1(grid_io_right_right_4_ccff_tail),
        .chanx_left_out(cbx_1__1__52_chanx_left_out),
        .chany_bottom_out(cby_8__1__3_chany_bottom_out),
        .chany_top_out_0(sb_8__1__3_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[48:51]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[48:51]),
        .left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    right_tile tile_9__6_
    (
        .ccff_head_0_0(cbx_1__1__52_ccff_tail),
        .ccff_head_1(grid_io_right_right_4_ccff_tail),
        .ccff_head_2(grid_clb_60_ccff_tail),
        .chanx_left_in(sb_1__1__46_chanx_right_out),
        .chany_bottom_in(sb_8__1__3_chany_top_out),
        .chany_top_in_0(cby_8__1__5_chany_bottom_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[44:47]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_60_ccff_tail),
        .ccff_tail_0(cbx_1__1__53_ccff_tail),
        .ccff_tail_1(grid_io_right_right_3_ccff_tail),
        .chanx_left_out(cbx_1__1__53_chanx_left_out),
        .chany_bottom_out(cby_8__1__4_chany_bottom_out),
        .chany_top_out_0(sb_8__1__4_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[44:47]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[44:47]),
        .left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    right_tile tile_9__7_
    (
        .ccff_head_0_0(cbx_1__1__53_ccff_tail),
        .ccff_head_1(grid_io_right_right_3_ccff_tail),
        .ccff_head_2(grid_clb_54_ccff_tail),
        .chanx_left_in(sb_1__1__47_chanx_right_out),
        .chany_bottom_in(sb_8__1__4_chany_top_out),
        .chany_top_in_0(cby_8__1__6_chany_bottom_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[40:43]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_61_ccff_tail),
        .ccff_tail_0(cbx_1__1__54_ccff_tail),
        .ccff_tail_1(grid_io_right_right_2_ccff_tail),
        .chanx_left_out(cbx_1__1__54_chanx_left_out),
        .chany_bottom_out(cby_8__1__5_chany_bottom_out),
        .chany_top_out_0(sb_8__1__5_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[40:43]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[40:43]),
        .left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    right_tile tile_9__8_
    (
        .ccff_head_0_0(cbx_1__1__54_ccff_tail),
        .ccff_head_1(grid_io_right_right_2_ccff_tail),
        .ccff_head_2(grid_clb_62_ccff_tail),
        .chanx_left_in(sb_1__1__48_chanx_right_out),
        .chany_bottom_in(sb_8__1__5_chany_top_out),
        .chany_top_in_0(cby_8__1__7_chany_bottom_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[36:39]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .scan_enable(scan_enable),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_12_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_13_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_14_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_15_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_),
        .top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .ccff_tail(grid_clb_62_ccff_tail),
        .ccff_tail_0(cbx_1__1__55_ccff_tail),
        .ccff_tail_1(grid_io_right_right_1_ccff_tail),
        .chanx_left_out(cbx_1__1__55_chanx_left_out),
        .chany_bottom_out(cby_8__1__6_chany_bottom_out),
        .chany_top_out_0(sb_8__1__6_chany_top_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[36:39]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[36:39]),
        .left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_7_)
    );
    top_right_tile tile_9__9_
    (
        .ccff_head_0_0(cbx_1__1__55_ccff_tail),
        .ccff_head_1(grid_io_right_right_1_ccff_tail),
        .chanx_left_in(sb_1__8__6_chanx_right_out),
        .chany_bottom_in(sb_8__1__6_chany_top_out),
        .clk0(clk),
        .gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[28:31]),
        .gfpga_pad_io_soc_in_0(gfpga_pad_io_soc_in[32:35]),
        .isol_n(isol_n),
        .prog_clk(prog_clk),
        .prog_reset(),
        .reset(),
        .scan_enable(scan_enable),
        .top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_8__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
        .top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_8__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
        .top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_),
        .bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
        .bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
        .bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
        .bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
        .ccff_tail(grid_clb_63_ccff_tail),
        .ccff_tail_0(grid_io_top_top_7_ccff_tail),
        .chanx_left_out(cbx_1__8__7_chanx_left_out),
        .chany_bottom_out(cby_8__1__7_chany_bottom_out),
        .gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[28:31]),
        .gfpga_pad_io_soc_dir_0(gfpga_pad_io_soc_dir[32:35]),
        .gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[28:31]),
        .gfpga_pad_io_soc_out_0(gfpga_pad_io_soc_out[32:35]),
        .left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
        .left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
        .left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
        .left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
        .right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_),
        .right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_),
        .right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_12_),
        .right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_13_),
        .right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_14_),
        .right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_15_),
        .right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_),
        .right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_),
        .top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_),
        .top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_),
        .top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_),
        .top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_),
        .top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_),
        .top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_),
        .top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_6_),
        .top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_7_)
    );
endmodule

